// This is the unpowered netlist.
module fp_sqr (act,
    clk,
    done,
    inexact,
    inv,
    ov,
    rst,
    un,
    in1,
    out,
    round_m);
 input act;
 input clk;
 output done;
 output inexact;
 output inv;
 output ov;
 input rst;
 output un;
 input [31:0] in1;
 output [31:0] out;
 input [2:0] round_m;

 wire net82;
 wire \M00r[10] ;
 wire \M00r[11] ;
 wire \M00r[12] ;
 wire \M00r[13] ;
 wire \M00r[14] ;
 wire \M00r[15] ;
 wire \M00r[16] ;
 wire \M00r[17] ;
 wire \M00r[18] ;
 wire \M00r[19] ;
 wire \M00r[1] ;
 wire \M00r[20] ;
 wire \M00r[21] ;
 wire \M00r[22] ;
 wire \M00r[23] ;
 wire \M00r[24] ;
 wire \M00r[2] ;
 wire \M00r[3] ;
 wire \M00r[4] ;
 wire \M00r[5] ;
 wire \M00r[6] ;
 wire \M00r[7] ;
 wire \M00r[8] ;
 wire \M00r[9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire done0_r;
 wire forward;
 wire forward_c;
 wire inv_f;
 wire inv_f_c;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net242;
 wire net245;
 wire net248;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \out_f[22] ;
 wire \out_f_c[22] ;
 wire ov_f;
 wire ov_f_c;
 wire \sq.out[10] ;
 wire \sq.out[11] ;
 wire \sq.out[12] ;
 wire \sq.out[13] ;
 wire \sq.out[14] ;
 wire \sq.out[15] ;
 wire \sq.out[16] ;
 wire \sq.out[17] ;
 wire \sq.out[18] ;
 wire \sq.out[19] ;
 wire \sq.out[1] ;
 wire \sq.out[20] ;
 wire \sq.out[21] ;
 wire \sq.out[22] ;
 wire \sq.out[23] ;
 wire \sq.out[24] ;
 wire \sq.out[2] ;
 wire \sq.out[3] ;
 wire \sq.out[4] ;
 wire \sq.out[5] ;
 wire \sq.out[6] ;
 wire \sq.out[7] ;
 wire \sq.out[8] ;
 wire \sq.out[9] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__B (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06142__B (.DIODE(_00578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06148__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__A (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06158__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06159__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06161__A1 (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06166__A (.DIODE(_00837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06167__A (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06168__B (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06170__A (.DIODE(_00837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06170__B (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06171__A1 (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06175__B (.DIODE(_00933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06176__A (.DIODE(_00933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__A (.DIODE(_00933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__B (.DIODE(_00740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__C (.DIODE(_00837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06183__A (.DIODE(_01008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06184__B (.DIODE(_01008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06190__A (.DIODE(_01095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06197__B (.DIODE(_01095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06198__A (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06199__B (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06202__B_N (.DIODE(_01171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06203__A (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06204__B (.DIODE(_01223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06207__A1 (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06361__C (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06367__B (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06381__B (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06388__B (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__C (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06438__A (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06444__B (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06453__B (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06459__B (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06460__B (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__B (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06478__B (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__S (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__A2 (.DIODE(_04484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__C (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__A (.DIODE(_04484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06514__A (.DIODE(_04484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__A (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__A (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__B (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__C (.DIODE(_04484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__B (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06592__B (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__C (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__B (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__C (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__C (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__C (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__B (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__C (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06633__S (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__A (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__B (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__B (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__C (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__C (.DIODE(_04484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__B (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__C (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__B (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__C (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__A (.DIODE(_04484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__B (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__C (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__C (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__C (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__C (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__S (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__B (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__C (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__B (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__B (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__C (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__A1 (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__A2 (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__B (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__B (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__B (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__C (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__A (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__C (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A (.DIODE(_04484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__C (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__C (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__C (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__C (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__B (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__C (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__C (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__C (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__B (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A (.DIODE(_02961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__C (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__B (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__A (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__C (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__B (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__C (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__S (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__C (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__B (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__C (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__C (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__C (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__C (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__B (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__C (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__C (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__C (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__A (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__C (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__B (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__B (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__B (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__C (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__C (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A1 (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A2 (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__B1 (.DIODE(_05761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07165__C (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__C (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__B (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__C (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__B (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A0 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__S (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__S (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__B (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__C (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__C (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__C (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__B (.DIODE(_00238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__B (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__B (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B (.DIODE(_00086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__C (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__C (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__A (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__C (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__C (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__C (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__C (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__C (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__C (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__B (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__C (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__C (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__C (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__C (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__C (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__C (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__A (.DIODE(_04220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__B (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__A (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A (.DIODE(_03782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07451__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__A (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__B (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__C (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B (.DIODE(_00578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A1 (.DIODE(_00578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__S (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__C (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__B (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A (.DIODE(_00237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__C (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__B (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__A (.DIODE(_06036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__C (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__C (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__C (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__C (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__C (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__C (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__C (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__C (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__C (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__C (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__B (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__B (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__B (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__B (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__B (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__B (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__A (.DIODE(_00749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__C (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__B (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__B (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A (.DIODE(_00749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A (.DIODE(_00749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__A1 (.DIODE(_00749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__B (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__C (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__A (.DIODE(_00718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__C (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__C (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__C (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__C (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__C (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__A (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__C (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__C (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__B (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__B (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__C (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__B (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__C (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__A (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__C (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__A (.DIODE(_06020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__C (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__C (.DIODE(_05119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__C (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__C (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__A (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__C (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__B (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__B (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__C (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__C (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__B (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A1 (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__B (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__A2 (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__B (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__C (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__B (.DIODE(_00845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__B (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__C (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__C (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__B (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__C (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__C (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__C (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__B (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__C (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__C (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__C (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__C (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__B (.DIODE(_00749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__B (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__C (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__A (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__C (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__C (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__C (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__C (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__C (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__C (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__C (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__B (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__C (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__A (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__B (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__A (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__B (.DIODE(_00749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A (.DIODE(_00425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08169__B (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__B (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A (.DIODE(_00283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08223__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__B1 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__B1 (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__C (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__B (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A1 (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__B (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__B (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__B (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__B (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__B (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__B (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__B (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__B (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__B (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__B (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__B (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__B (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__B (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__C (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__B (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__C (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__C (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A1 (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__B (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__B (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A2 (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__B (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A (.DIODE(_00749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__B (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__B (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__C (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__B (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__B (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08469__B (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08471__B (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__B (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08484__B (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08496__A (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08498__B (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__C (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08512__B (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__B (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__B (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__B (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__B1 (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__B (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08549__B (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__B (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A (.DIODE(_00214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__B (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__B (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__B (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B_N (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__A (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__A (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__B (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A1 (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__B (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08651__A (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__B (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A2 (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__C (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08678__C1 (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__B (.DIODE(_01843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A (.DIODE(_01843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__A (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__C (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08690__A (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__A (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__A (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__B (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08694__B (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08696__B (.DIODE(_01843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__B (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__B (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__C (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__A1 (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__A2 (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__B (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__C (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__A (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__B (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__C (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__B (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08712__B (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__A (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__B (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__B (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__A (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__B (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__B (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__A (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A2 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__B (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__B (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__B (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__B (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__B (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__A1 (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__A (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__B (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__A1 (.DIODE(_01758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__A2 (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__A (.DIODE(_00743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A (.DIODE(_01855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08828__B (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08830__A (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08838__A (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08844__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A (.DIODE(_00460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__B (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__B (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__A (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__B (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A1 (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__A (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A1 (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A (.DIODE(_02050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__B (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A2 (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__B (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__A (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A2 (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A (.DIODE(_01344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__B (.DIODE(_01843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A (.DIODE(_02050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__B (.DIODE(_01843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08912__B1 (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08914__C (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__D (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__B (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__B_N (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__A (.DIODE(_01524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__B (.DIODE(_01843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A1 (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__B1 (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__C1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__B (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08944__B (.DIODE(_00091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__B (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__B (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__B (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__B (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__A (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08964__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__B (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__B (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__A (.DIODE(_06002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09008__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__C (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__C (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__B (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__B (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__B (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__C (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__A (.DIODE(_02050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09067__A (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A2 (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__B (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09085__B (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09089__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__C (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__B (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__B (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__B (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__B (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__A (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__B (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__C (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__A (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__B (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__A (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__B (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__B (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__A (.DIODE(_02108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__B (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__C (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__B (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__B (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__B (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09193__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(_01846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A2 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__B2 (.DIODE(_02109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__C1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__B (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__B (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__B (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__C (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A1 (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09278__A2 (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__A (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09280__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__A (.DIODE(_01644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__B (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__B (.DIODE(_02016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__B (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__C (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__C (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__B (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__B (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__B (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__A (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__A (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__B (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__B (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__B (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__B1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__B (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__A (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__B (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__B (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__A (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B (.DIODE(_02085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__C (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__B (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__A (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__B (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__B (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__A (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__A (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__B (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__B1 (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A1 (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__C (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__A (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A (.DIODE(_00843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__A (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__A2 (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09577__A (.DIODE(_01363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09578__B (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__A (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__A (.DIODE(_01286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__B (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__B (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A1 (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__A (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A (.DIODE(_01587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__B (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__S (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__B (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A2 (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A (.DIODE(_01240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__B (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__B (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09642__A (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__B1 (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09644__A (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__B (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A (.DIODE(_05130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__B (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A (.DIODE(_00455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__B (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A1 (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__B (.DIODE(_02767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__B (.DIODE(_02744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__A (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__B (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__B (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09714__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09728__S (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A1 (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__A2 (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__A (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__B (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A2 (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__C1 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__C (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__A (.DIODE(_03090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__A (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__B (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__A (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A (.DIODE(_03113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__B (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__B (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__A (.DIODE(_03090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__B (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A1 (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__A2 (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__B (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__C (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__A (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__B (.DIODE(_03090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__B (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__B (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09855__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09857__B (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__B (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B (.DIODE(_03090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__B (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__B1 (.DIODE(_03090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__B (.DIODE(_03113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__C (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__B (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__A (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__A (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A (.DIODE(_03113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__B (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__B (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__B (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__B (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__A (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A2 (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__A (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__B (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__A (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A2 (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__A (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09990__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__B (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__A (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10012__B (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__B (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A2 (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B1 (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A2 (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__B (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A1 (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__C (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10067__A (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__A2 (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__A (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__A (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A2 (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__A (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A1 (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A (.DIODE(_03117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A1 (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__B (.DIODE(_03204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__A (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A2 (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__B (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__A (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__C (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__A (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__B (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__A (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__B (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__B (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__C (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__A (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__B (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__A (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__B (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__B (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__C (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10191__B (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__B (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__B (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10285__B (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__B (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__A (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A2 (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__B (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__B1 (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A2 (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__B (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__B (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__B (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__B (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10368__A2 (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__B (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__B (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__A2 (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10389__A (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__A1 (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A (.DIODE(_03438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__B (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__A1 (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__B (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__A1 (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__S (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__B (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__A1 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__A (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__A (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__B (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__B (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__A (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__B (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__A1 (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__A2 (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__B (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__C (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10532__B (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10532__C (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10535__B (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__B (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__B (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__B (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__B (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__A (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A2 (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__B (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A1 (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A2 (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__A (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__B (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__B (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__S (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__B (.DIODE(_01712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__B (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__B (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A1 (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__B1 (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A2 (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__A1 (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__B (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__A1 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__B (.DIODE(_03662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10695__B (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__A2 (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__B (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10699__A2 (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__D1 (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__B (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__B (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__A2 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10756__A2 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10758__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__B (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__B (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__A (.DIODE(_03821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__A (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__A (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10838__B (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A2 (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__B (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__B (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__B1 (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__B (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__B (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__B (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__B (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__C (.DIODE(_03843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__B (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__C (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__B (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__A (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__A (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__B (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__B (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__B (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__B (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__B (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__B (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__B (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__B (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__B (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__B (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__A (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__B (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__B (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__B (.DIODE(_01081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__B (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__C (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A2 (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A2 (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__B1 (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11028__B (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__A (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__B (.DIODE(_04421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A (.DIODE(_04421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__B (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__B (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__B (.DIODE(_03439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__B (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__B (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__B (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__B (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__A (.DIODE(_03373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__A (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__B (.DIODE(_02898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__B (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__B (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__B (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__A2 (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__A (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__B (.DIODE(_02504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__A (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__A (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__B (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11220__B (.DIODE(_02345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__A1 (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__A (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__B (.DIODE(_02856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__A (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__B (.DIODE(_00844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__A2 (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__B (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__A (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B (.DIODE(_02843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__B (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__B (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__B (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11302__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__B (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__B (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__B (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11316__B (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__B (.DIODE(_02009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11320__B (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__A (.DIODE(_04421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11322__B (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__A (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__A (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11328__B (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__B (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__B (.DIODE(_01730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__B (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__B (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11346__A (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__B (.DIODE(_05140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__C1 (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__B (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A (.DIODE(_04601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A1 (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__B (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__A1 (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__A (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__B1 (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__B (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__B (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A1 (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__B (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11614__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11614__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11618__A2 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11618__B1 (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__A (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__11646__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__B1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__A (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11661__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A2 (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__B1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A2 (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__B1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__A1 (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A2 (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__B1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__B (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A2 (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11700__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11701__A2 (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11701__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__B (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11723__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__A (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__A1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__B (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__S (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__A1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__B (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__A (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__A1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__B1 (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11816__B (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__A (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__A1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__B1 (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__B (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__A (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__B (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__B1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A1 (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__B (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11893__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__B1 (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__A2 (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__B1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11918__B1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__B1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__A1 (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__B1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__A1 (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__B1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11962__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__A2 (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__B1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11982__A1 (.DIODE(_05057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__12003__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__B1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__B1 (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__B (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__A (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__B1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__B1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__B1 (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A2 (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__B1 (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__B1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__B (.DIODE(_05182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__B (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__B1 (.DIODE(_05177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__A2 (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__B (.DIODE(_05159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__A (.DIODE(_05162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A1 (.DIODE(_05164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__B1 (.DIODE(_05110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__A (.DIODE(_05094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__B (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__A (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__B (.DIODE(_05175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12124__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__B1 (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__B (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__B (.DIODE(_05106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A (.DIODE(_05085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__B (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A (.DIODE(_05124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__B (.DIODE(_05095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__B (.DIODE(_05063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__B1 (.DIODE(_05058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__A1 (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__A (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12180__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12188__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__C (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__B1 (.DIODE(_05170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__C (.DIODE(_05087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__C (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12214__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__C (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__C1 (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A (.DIODE(_01277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__A (.DIODE(\out_f_c[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__D (.DIODE(\out_f_c[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__D (.DIODE(\sq.out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__D (.DIODE(\sq.out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__D (.DIODE(\sq.out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__D (.DIODE(\sq.out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__D (.DIODE(\sq.out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__D (.DIODE(\sq.out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__D (.DIODE(\sq.out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__D (.DIODE(\sq.out[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__D (.DIODE(\sq.out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__D (.DIODE(\sq.out[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__D (.DIODE(\sq.out[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__D (.DIODE(\sq.out[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__D (.DIODE(\sq.out[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__D (.DIODE(\sq.out[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__D (.DIODE(\sq.out[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__D (.DIODE(\sq.out[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__D (.DIODE(\sq.out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__D (.DIODE(\sq.out[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__D (.DIODE(\sq.out[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__D (.DIODE(\sq.out[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__D (.DIODE(\sq.out[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__D (.DIODE(\sq.out[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__D (.DIODE(\sq.out[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__D (.DIODE(\sq.out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__RESET_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__RESET_B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__RESET_B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_split17_A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split18_A (.DIODE(_05173_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split1_A (.DIODE(_03090_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_992 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06118_ (.A(net11),
    .Y(_00325_));
 sky130_fd_sc_hd__inv_2 _06119_ (.A(net10),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _06120_ (.A(_00325_),
    .B(_00336_),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_2 _06121_ (.A(net14),
    .Y(_00358_));
 sky130_fd_sc_hd__inv_2 _06122_ (.A(net13),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _06123_ (.A(_00358_),
    .B(_00369_),
    .Y(_00380_));
 sky130_fd_sc_hd__or2_1 _06124_ (.A(net7),
    .B(net6),
    .X(_00391_));
 sky130_fd_sc_hd__or2_1 _06125_ (.A(net9),
    .B(net8),
    .X(_00402_));
 sky130_fd_sc_hd__or4_1 _06126_ (.A(_00347_),
    .B(_00380_),
    .C(_00391_),
    .D(_00402_),
    .X(_00413_));
 sky130_fd_sc_hd__nand2_1 _06127_ (.A(net18),
    .B(net19),
    .Y(_00424_));
 sky130_fd_sc_hd__inv_2 _06128_ (.A(net15),
    .Y(_00435_));
 sky130_fd_sc_hd__buf_8 _06129_ (.A(net16),
    .X(_00446_));
 sky130_fd_sc_hd__nand2_1 _06130_ (.A(_00435_),
    .B(_00446_),
    .Y(_00457_));
 sky130_fd_sc_hd__or2_1 _06131_ (.A(net28),
    .B(net27),
    .X(_00468_));
 sky130_fd_sc_hd__or2_1 _06132_ (.A(net26),
    .B(net23),
    .X(_00479_));
 sky130_fd_sc_hd__or4_1 _06133_ (.A(_00424_),
    .B(_00457_),
    .C(_00468_),
    .D(_00479_),
    .X(_00490_));
 sky130_fd_sc_hd__or2_1 _06134_ (.A(net3),
    .B(net2),
    .X(_00501_));
 sky130_fd_sc_hd__or2_1 _06135_ (.A(net5),
    .B(net4),
    .X(_00512_));
 sky130_fd_sc_hd__or2_1 _06136_ (.A(net30),
    .B(net29),
    .X(_00523_));
 sky130_fd_sc_hd__or2_1 _06137_ (.A(net32),
    .B(net31),
    .X(_00534_));
 sky130_fd_sc_hd__or4_1 _06138_ (.A(_00501_),
    .B(_00512_),
    .C(_00523_),
    .D(_00534_),
    .X(_00545_));
 sky130_fd_sc_hd__inv_2 _06139_ (.A(net24),
    .Y(_00556_));
 sky130_fd_sc_hd__inv_2 _06140_ (.A(net1),
    .Y(_00567_));
 sky130_fd_sc_hd__inv_2 _06141_ (.A(net12),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _06142_ (.A(_00567_),
    .B(_00578_),
    .Y(_00589_));
 sky130_fd_sc_hd__inv_2 _06143_ (.A(net17),
    .Y(_00599_));
 sky130_fd_sc_hd__inv_2 _06144_ (.A(net20),
    .Y(_00610_));
 sky130_fd_sc_hd__inv_2 _06145_ (.A(net22),
    .Y(_00620_));
 sky130_fd_sc_hd__inv_2 _06146_ (.A(net21),
    .Y(_00631_));
 sky130_fd_sc_hd__or4_1 _06147_ (.A(_00599_),
    .B(_00610_),
    .C(_00620_),
    .D(_00631_),
    .X(_00642_));
 sky130_fd_sc_hd__or4_1 _06148_ (.A(net25),
    .B(_00556_),
    .C(_00589_),
    .D(_00642_),
    .X(_00653_));
 sky130_fd_sc_hd__or4_1 _06149_ (.A(_00413_),
    .B(_00490_),
    .C(_00545_),
    .D(_00653_),
    .X(_00664_));
 sky130_fd_sc_hd__clkbuf_4 _06150_ (.A(_00664_),
    .X(\out_f_c[22] ));
 sky130_fd_sc_hd__clkinv_4 _06151_ (.A(net16),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_2 _06152_ (.A(_00685_),
    .B(_00599_),
    .Y(_00696_));
 sky130_fd_sc_hd__buf_6 _06153_ (.A(net113),
    .X(_00707_));
 sky130_fd_sc_hd__buf_6 _06154_ (.A(_00707_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_2 _06155_ (.A(_00718_),
    .B(net17),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_8 _06156_ (.A(_00696_),
    .B(_00729_),
    .Y(_00740_));
 sky130_fd_sc_hd__clkbuf_1 _06157_ (.A(net132),
    .X(_00751_));
 sky130_fd_sc_hd__inv_2 _06158_ (.A(net133),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _06159_ (.A(net123),
    .B(net133),
    .Y(_00773_));
 sky130_fd_sc_hd__inv_2 _06160_ (.A(net134),
    .Y(_00783_));
 sky130_fd_sc_hd__a21o_1 _06161_ (.A1(_00740_),
    .A2(_00762_),
    .B1(_00783_),
    .X(_00017_));
 sky130_fd_sc_hd__inv_2 _06162_ (.A(net18),
    .Y(_00804_));
 sky130_fd_sc_hd__or2_1 _06163_ (.A(_00804_),
    .B(_00729_),
    .X(_00815_));
 sky130_fd_sc_hd__nand2_1 _06164_ (.A(_00729_),
    .B(_00804_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_4 _06165_ (.A(_00815_),
    .B(_00826_),
    .Y(_00837_));
 sky130_fd_sc_hd__inv_2 _06166_ (.A(_00837_),
    .Y(_00847_));
 sky130_fd_sc_hd__or2_1 _06167_ (.A(_00740_),
    .B(_00847_),
    .X(_00858_));
 sky130_fd_sc_hd__nand2_1 _06168_ (.A(_00847_),
    .B(_00740_),
    .Y(_00869_));
 sky130_fd_sc_hd__a31o_1 _06169_ (.A1(_00858_),
    .A2(_00762_),
    .A3(_00869_),
    .B1(_00783_),
    .X(_00018_));
 sky130_fd_sc_hd__nand2_1 _06170_ (.A(_00837_),
    .B(_00740_),
    .Y(_00890_));
 sky130_fd_sc_hd__a31o_1 _06171_ (.A1(_00718_),
    .A2(net18),
    .A3(net17),
    .B1(net19),
    .X(_00900_));
 sky130_fd_sc_hd__nor2_1 _06172_ (.A(_00424_),
    .B(_00729_),
    .Y(_00911_));
 sky130_fd_sc_hd__inv_2 _06173_ (.A(_00911_),
    .Y(_00922_));
 sky130_fd_sc_hd__nand2_4 _06174_ (.A(_00900_),
    .B(_00922_),
    .Y(_00933_));
 sky130_fd_sc_hd__or2_1 _06175_ (.A(_00890_),
    .B(_00933_),
    .X(_00944_));
 sky130_fd_sc_hd__nand2_1 _06176_ (.A(_00933_),
    .B(_00890_),
    .Y(_00955_));
 sky130_fd_sc_hd__a31o_1 _06177_ (.A1(_00944_),
    .A2(_00762_),
    .A3(_00955_),
    .B1(_00783_),
    .X(_00019_));
 sky130_fd_sc_hd__nor2_1 _06178_ (.A(net20),
    .B(_00911_),
    .Y(_00975_));
 sky130_fd_sc_hd__nor2_1 _06179_ (.A(_00610_),
    .B(_00922_),
    .Y(_00986_));
 sky130_fd_sc_hd__nor2_1 _06180_ (.A(_00975_),
    .B(_00986_),
    .Y(_00997_));
 sky130_fd_sc_hd__inv_2 _06181_ (.A(_00997_),
    .Y(_01008_));
 sky130_fd_sc_hd__and3_1 _06182_ (.A(_00933_),
    .B(_00740_),
    .C(_00837_),
    .X(_01019_));
 sky130_fd_sc_hd__nor2_1 _06183_ (.A(_01008_),
    .B(_01019_),
    .Y(_01030_));
 sky130_fd_sc_hd__and2_1 _06184_ (.A(_01019_),
    .B(_01008_),
    .X(_01041_));
 sky130_fd_sc_hd__o21ai_1 _06185_ (.A1(_01030_),
    .A2(_01041_),
    .B1(_00762_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand2_1 _06186_ (.A(_01052_),
    .B(net134),
    .Y(_00020_));
 sky130_fd_sc_hd__or2_1 _06187_ (.A(net21),
    .B(_00986_),
    .X(_01073_));
 sky130_fd_sc_hd__nand2_1 _06188_ (.A(_00986_),
    .B(net21),
    .Y(_01084_));
 sky130_fd_sc_hd__nand2_4 _06189_ (.A(_01073_),
    .B(_01084_),
    .Y(_01095_));
 sky130_fd_sc_hd__inv_2 _06190_ (.A(_01095_),
    .Y(_01106_));
 sky130_fd_sc_hd__or2_1 _06191_ (.A(_01106_),
    .B(_01041_),
    .X(_01117_));
 sky130_fd_sc_hd__nand2_1 _06192_ (.A(_01041_),
    .B(_01106_),
    .Y(_01128_));
 sky130_fd_sc_hd__a31o_1 _06193_ (.A1(_01117_),
    .A2(_00762_),
    .A3(_01128_),
    .B1(_00783_),
    .X(_00021_));
 sky130_fd_sc_hd__or2_2 _06194_ (.A(_00620_),
    .B(_01084_),
    .X(_01149_));
 sky130_fd_sc_hd__nand2_1 _06195_ (.A(_01084_),
    .B(_00620_),
    .Y(_01160_));
 sky130_fd_sc_hd__nand2_4 _06196_ (.A(_01149_),
    .B(_01160_),
    .Y(_01171_));
 sky130_fd_sc_hd__nand2_1 _06197_ (.A(_01041_),
    .B(_01095_),
    .Y(_01182_));
 sky130_fd_sc_hd__or2_1 _06198_ (.A(_01171_),
    .B(_01182_),
    .X(_01193_));
 sky130_fd_sc_hd__nand2_1 _06199_ (.A(_01182_),
    .B(_01171_),
    .Y(_01203_));
 sky130_fd_sc_hd__a31o_1 _06200_ (.A1(_01193_),
    .A2(_00762_),
    .A3(_01203_),
    .B1(_00783_),
    .X(_00022_));
 sky130_fd_sc_hd__xor2_4 _06201_ (.A(_00556_),
    .B(_01149_),
    .X(_01223_));
 sky130_fd_sc_hd__or2b_1 _06202_ (.A(_01182_),
    .B_N(_01171_),
    .X(_01234_));
 sky130_fd_sc_hd__or2_1 _06203_ (.A(_01223_),
    .B(_01234_),
    .X(_01245_));
 sky130_fd_sc_hd__nand2_1 _06204_ (.A(_01234_),
    .B(_01223_),
    .Y(_01256_));
 sky130_fd_sc_hd__a31o_1 _06205_ (.A1(_01245_),
    .A2(_00762_),
    .A3(_01256_),
    .B1(_00783_),
    .X(_00023_));
 sky130_fd_sc_hd__buf_6 _06206_ (.A(net137),
    .X(_01277_));
 sky130_fd_sc_hd__o21ai_1 _06207_ (.A1(_01277_),
    .A2(_01256_),
    .B1(net134),
    .Y(_00025_));
 sky130_fd_sc_hd__inv_2 _06208_ (.A(net142),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _06209_ (.A(net11),
    .B(net16),
    .Y(_01309_));
 sky130_fd_sc_hd__o21ai_4 _06210_ (.A1(net16),
    .A2(_00336_),
    .B1(_01309_),
    .Y(_01320_));
 sky130_fd_sc_hd__mux2_1 _06211_ (.A0(net9),
    .A1(net10),
    .S(_00707_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _06212_ (.A0(net8),
    .A1(net9),
    .S(net113),
    .X(_01342_));
 sky130_fd_sc_hd__buf_6 _06213_ (.A(_01342_),
    .X(_01353_));
 sky130_fd_sc_hd__or2_1 _06214_ (.A(_01331_),
    .B(_01353_),
    .X(_01364_));
 sky130_fd_sc_hd__nor2_1 _06215_ (.A(_01320_),
    .B(_01364_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _06216_ (.A(_00358_),
    .B(_00446_),
    .Y(_01386_));
 sky130_fd_sc_hd__o21ai_2 _06217_ (.A1(net13),
    .A2(_00446_),
    .B1(_01386_),
    .Y(_01397_));
 sky130_fd_sc_hd__a31oi_4 _06218_ (.A1(_00358_),
    .A2(_00369_),
    .A3(_00435_),
    .B1(_00446_),
    .Y(_01408_));
 sky130_fd_sc_hd__o211ai_1 _06219_ (.A1(net14),
    .A2(net15),
    .B1(_00369_),
    .C1(_00685_),
    .Y(_01419_));
 sky130_fd_sc_hd__o21ai_2 _06220_ (.A1(net14),
    .A2(_00446_),
    .B1(_00457_),
    .Y(_01430_));
 sky130_fd_sc_hd__inv_2 _06221_ (.A(_01430_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _06222_ (.A(_01419_),
    .B(_01441_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand3_2 _06223_ (.A(_01430_),
    .B(_01397_),
    .C(net15),
    .Y(_01463_));
 sky130_fd_sc_hd__nand2_1 _06224_ (.A(_01452_),
    .B(_01463_),
    .Y(_01474_));
 sky130_fd_sc_hd__o21ai_1 _06225_ (.A1(_01397_),
    .A2(_01408_),
    .B1(_01474_),
    .Y(_01485_));
 sky130_fd_sc_hd__and4_1 _06226_ (.A(_00685_),
    .B(net14),
    .C(net13),
    .D(net15),
    .X(_01496_));
 sky130_fd_sc_hd__clkinvlp_2 _06227_ (.A(_01496_),
    .Y(_01507_));
 sky130_fd_sc_hd__a31oi_1 _06228_ (.A1(_00358_),
    .A2(_00369_),
    .A3(net15),
    .B1(_00446_),
    .Y(_01518_));
 sky130_fd_sc_hd__o211ai_1 _06229_ (.A1(net14),
    .A2(net13),
    .B1(_00435_),
    .C1(_00685_),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_1 _06230_ (.A(_01518_),
    .B(_01529_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand3_1 _06231_ (.A(_01540_),
    .B(_01452_),
    .C(_01463_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand3_1 _06232_ (.A(_01485_),
    .B(_01507_),
    .C(_01551_),
    .Y(_01562_));
 sky130_fd_sc_hd__nand2_1 _06233_ (.A(net13),
    .B(_00446_),
    .Y(_01573_));
 sky130_fd_sc_hd__o21ai_2 _06234_ (.A1(net16),
    .A2(_00325_),
    .B1(_01573_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _06235_ (.A(_01584_),
    .B(_01320_),
    .Y(_01595_));
 sky130_fd_sc_hd__a211o_1 _06236_ (.A1(_00685_),
    .A2(net13),
    .B1(net14),
    .C1(_00435_),
    .X(_01606_));
 sky130_fd_sc_hd__o21a_1 _06237_ (.A1(_01595_),
    .A2(_01606_),
    .B1(_01507_),
    .X(_01617_));
 sky130_fd_sc_hd__nand2_1 _06238_ (.A(_01562_),
    .B(_01617_),
    .Y(_01628_));
 sky130_fd_sc_hd__buf_6 _06239_ (.A(_01628_),
    .X(_01639_));
 sky130_fd_sc_hd__xor2_1 _06240_ (.A(_01584_),
    .B(_01320_),
    .X(_01650_));
 sky130_fd_sc_hd__inv_2 _06241_ (.A(_01650_),
    .Y(_01661_));
 sky130_fd_sc_hd__nand2_2 _06242_ (.A(_01639_),
    .B(_01661_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand3_1 _06243_ (.A(_01562_),
    .B(_01584_),
    .C(_01617_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand2_2 _06244_ (.A(_01672_),
    .B(_01683_),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _06245_ (.A(_01694_),
    .B(_01408_),
    .Y(_01705_));
 sky130_fd_sc_hd__clkinvlp_2 _06246_ (.A(_01320_),
    .Y(_01716_));
 sky130_fd_sc_hd__inv_4 _06247_ (.A(_01639_),
    .Y(_01727_));
 sky130_fd_sc_hd__nor2_1 _06248_ (.A(_01716_),
    .B(_01727_),
    .Y(_01738_));
 sky130_fd_sc_hd__inv_2 _06249_ (.A(_01738_),
    .Y(_01749_));
 sky130_fd_sc_hd__inv_2 _06250_ (.A(_01408_),
    .Y(_01760_));
 sky130_fd_sc_hd__nand3_1 _06251_ (.A(_01672_),
    .B(_01760_),
    .C(_01683_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand3_1 _06252_ (.A(_01705_),
    .B(_01749_),
    .C(_01770_),
    .Y(_01780_));
 sky130_fd_sc_hd__nand2_1 _06253_ (.A(_01694_),
    .B(_01760_),
    .Y(_01791_));
 sky130_fd_sc_hd__nand3_2 _06254_ (.A(_01672_),
    .B(_01408_),
    .C(_01683_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand3_1 _06255_ (.A(_01791_),
    .B(_01802_),
    .C(_01738_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _06256_ (.A(_01780_),
    .B(_01812_),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_2 _06257_ (.A(_01375_),
    .B(_01823_),
    .Y(_01834_));
 sky130_fd_sc_hd__o21ai_1 _06258_ (.A1(_00358_),
    .A2(_00685_),
    .B1(_01419_),
    .Y(_01845_));
 sky130_fd_sc_hd__inv_2 _06259_ (.A(_01397_),
    .Y(_01856_));
 sky130_fd_sc_hd__inv_2 _06260_ (.A(_01595_),
    .Y(_01865_));
 sky130_fd_sc_hd__nor2_1 _06261_ (.A(_01856_),
    .B(_01865_),
    .Y(_01876_));
 sky130_fd_sc_hd__inv_2 _06262_ (.A(_01876_),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_1 _06263_ (.A(_01865_),
    .B(_01856_),
    .Y(_01898_));
 sky130_fd_sc_hd__and2_1 _06264_ (.A(_01887_),
    .B(_01898_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_1 _06265_ (.A(_01639_),
    .B(_01909_),
    .Y(_01920_));
 sky130_fd_sc_hd__o21ai_2 _06266_ (.A1(_01845_),
    .A2(_01628_),
    .B1(_01920_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _06267_ (.A(net112),
    .B(_00369_),
    .Y(_01942_));
 sky130_fd_sc_hd__or2_1 _06268_ (.A(_01942_),
    .B(_01474_),
    .X(_01953_));
 sky130_fd_sc_hd__nand2_1 _06269_ (.A(_01474_),
    .B(_01942_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _06270_ (.A(_01953_),
    .B(_01964_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _06271_ (.A(_01975_),
    .B(_01876_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand3_1 _06272_ (.A(_01953_),
    .B(_01964_),
    .C(_01887_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand2_1 _06273_ (.A(_01986_),
    .B(_01997_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2_1 _06274_ (.A(_02008_),
    .B(_01639_),
    .Y(_02019_));
 sky130_fd_sc_hd__nand2_1 _06275_ (.A(_02019_),
    .B(_01551_),
    .Y(_02029_));
 sky130_fd_sc_hd__nor2_1 _06276_ (.A(_01931_),
    .B(_02029_),
    .Y(_02040_));
 sky130_fd_sc_hd__inv_2 _06277_ (.A(_02040_),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _06278_ (.A(_02029_),
    .B(_01931_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _06279_ (.A(_02051_),
    .B(_02062_),
    .Y(_02073_));
 sky130_fd_sc_hd__inv_2 _06280_ (.A(_02073_),
    .Y(_02084_));
 sky130_fd_sc_hd__nor2_1 _06281_ (.A(_01802_),
    .B(_01931_),
    .Y(_02095_));
 sky130_fd_sc_hd__nand2_1 _06282_ (.A(_01802_),
    .B(_01931_),
    .Y(_02106_));
 sky130_fd_sc_hd__inv_2 _06283_ (.A(_02106_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _06284_ (.A(_02095_),
    .B(_02117_),
    .Y(_02128_));
 sky130_fd_sc_hd__nand3_2 _06285_ (.A(_01834_),
    .B(_02084_),
    .C(_02128_),
    .Y(_02139_));
 sky130_fd_sc_hd__o21bai_1 _06286_ (.A1(_02095_),
    .A2(_01780_),
    .B1_N(_02117_),
    .Y(_02150_));
 sky130_fd_sc_hd__nand2_1 _06287_ (.A(_02150_),
    .B(_02084_),
    .Y(_02161_));
 sky130_fd_sc_hd__nand3_4 _06288_ (.A(_02139_),
    .B(_02051_),
    .C(_02161_),
    .Y(_02171_));
 sky130_fd_sc_hd__xor2_1 _06289_ (.A(_01331_),
    .B(_01353_),
    .X(_02182_));
 sky130_fd_sc_hd__inv_2 _06290_ (.A(_02182_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand2_1 _06291_ (.A(_02171_),
    .B(_02193_),
    .Y(_02204_));
 sky130_fd_sc_hd__a21oi_2 _06292_ (.A1(_02150_),
    .A2(_02084_),
    .B1(_02040_),
    .Y(_02215_));
 sky130_fd_sc_hd__nand3_1 _06293_ (.A(_02215_),
    .B(_01331_),
    .C(net92),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _06294_ (.A(_02204_),
    .B(_02226_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_1 _06295_ (.A(_02237_),
    .B(_01727_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand3_1 _06296_ (.A(_02215_),
    .B(_01353_),
    .C(net93),
    .Y(_02259_));
 sky130_fd_sc_hd__mux2_1 _06297_ (.A0(net7),
    .A1(net8),
    .S(_00707_),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _06298_ (.A0(net6),
    .A1(net7),
    .S(_00707_),
    .X(_02281_));
 sky130_fd_sc_hd__buf_6 _06299_ (.A(_02281_),
    .X(_02291_));
 sky130_fd_sc_hd__nor2_1 _06300_ (.A(_02270_),
    .B(_02291_),
    .Y(_02302_));
 sky130_fd_sc_hd__nand2_1 _06301_ (.A(_02259_),
    .B(_02302_),
    .Y(_02313_));
 sky130_fd_sc_hd__buf_6 _06302_ (.A(_02171_),
    .X(_02324_));
 sky130_fd_sc_hd__nand2_1 _06303_ (.A(_02324_),
    .B(_01353_),
    .Y(_02335_));
 sky130_fd_sc_hd__nand2_1 _06304_ (.A(_02313_),
    .B(_02335_),
    .Y(_02346_));
 sky130_fd_sc_hd__nand3_2 _06305_ (.A(_02204_),
    .B(_02226_),
    .C(_01639_),
    .Y(_02357_));
 sky130_fd_sc_hd__nand3_2 _06306_ (.A(_02248_),
    .B(_02346_),
    .C(_02357_),
    .Y(_02368_));
 sky130_fd_sc_hd__inv_2 _06307_ (.A(_02368_),
    .Y(_02379_));
 sky130_fd_sc_hd__inv_2 _06308_ (.A(_01375_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand2_1 _06309_ (.A(_01364_),
    .B(_01320_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand2_1 _06310_ (.A(_02390_),
    .B(_02401_),
    .Y(_02412_));
 sky130_fd_sc_hd__inv_2 _06311_ (.A(_02412_),
    .Y(_02423_));
 sky130_fd_sc_hd__nand2_1 _06312_ (.A(_02324_),
    .B(_02423_),
    .Y(_02434_));
 sky130_fd_sc_hd__nand2_1 _06313_ (.A(_01727_),
    .B(_01320_),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _06314_ (.A(_01639_),
    .B(_01716_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _06315_ (.A(_02445_),
    .B(_02456_),
    .Y(_02467_));
 sky130_fd_sc_hd__clkinvlp_2 _06316_ (.A(_02467_),
    .Y(_02478_));
 sky130_fd_sc_hd__nand3_1 _06317_ (.A(_02215_),
    .B(_02478_),
    .C(net92),
    .Y(_02489_));
 sky130_fd_sc_hd__nand3_2 _06318_ (.A(_02434_),
    .B(_02489_),
    .C(_01408_),
    .Y(_02499_));
 sky130_fd_sc_hd__nand2_1 _06319_ (.A(_02324_),
    .B(_02412_),
    .Y(_02510_));
 sky130_fd_sc_hd__nand3_1 _06320_ (.A(_02215_),
    .B(_02467_),
    .C(net92),
    .Y(_02521_));
 sky130_fd_sc_hd__nand3_1 _06321_ (.A(_02510_),
    .B(_02521_),
    .C(_01760_),
    .Y(_02532_));
 sky130_fd_sc_hd__nand2_1 _06322_ (.A(_02499_),
    .B(_02532_),
    .Y(_02543_));
 sky130_fd_sc_hd__inv_2 _06323_ (.A(net119),
    .Y(_02554_));
 sky130_fd_sc_hd__nand2_1 _06324_ (.A(_02543_),
    .B(_02554_),
    .Y(_02565_));
 sky130_fd_sc_hd__nand3_2 _06325_ (.A(_02357_),
    .B(_02499_),
    .C(_02532_),
    .Y(_02576_));
 sky130_fd_sc_hd__nand2_1 _06326_ (.A(_02565_),
    .B(_02576_),
    .Y(_02587_));
 sky130_fd_sc_hd__nor2_2 _06327_ (.A(_02379_),
    .B(_02587_),
    .Y(_02598_));
 sky130_fd_sc_hd__and2_1 _06328_ (.A(_01823_),
    .B(_01375_),
    .X(_02609_));
 sky130_fd_sc_hd__or2_1 _06329_ (.A(_01834_),
    .B(_02609_),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_1 _06330_ (.A(_02171_),
    .B(_02620_),
    .Y(_02631_));
 sky130_fd_sc_hd__o21ai_2 _06331_ (.A1(_01694_),
    .A2(_02171_),
    .B1(_02631_),
    .Y(_02642_));
 sky130_fd_sc_hd__inv_2 _06332_ (.A(_02642_),
    .Y(_02653_));
 sky130_fd_sc_hd__inv_2 _06333_ (.A(_02128_),
    .Y(_02664_));
 sky130_fd_sc_hd__a21boi_1 _06334_ (.A1(_02390_),
    .A2(_01812_),
    .B1_N(_01780_),
    .Y(_02675_));
 sky130_fd_sc_hd__or2_1 _06335_ (.A(_02664_),
    .B(_02675_),
    .X(_02686_));
 sky130_fd_sc_hd__nand2_1 _06336_ (.A(_02675_),
    .B(_02664_),
    .Y(_02697_));
 sky130_fd_sc_hd__nand3_1 _06337_ (.A(_02324_),
    .B(_02686_),
    .C(_02697_),
    .Y(_02708_));
 sky130_fd_sc_hd__o21ai_1 _06338_ (.A1(_01931_),
    .A2(_02324_),
    .B1(_02708_),
    .Y(_02719_));
 sky130_fd_sc_hd__nor2_1 _06339_ (.A(_02653_),
    .B(_02719_),
    .Y(_02730_));
 sky130_fd_sc_hd__nand2_1 _06340_ (.A(_02719_),
    .B(_02653_),
    .Y(_02741_));
 sky130_fd_sc_hd__inv_2 _06341_ (.A(_02741_),
    .Y(_02752_));
 sky130_fd_sc_hd__nor2_1 _06342_ (.A(_02730_),
    .B(_02752_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_1 _06343_ (.A(_02434_),
    .B(_02489_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_2 _06344_ (.A(_02774_),
    .B(_01408_),
    .Y(_02785_));
 sky130_fd_sc_hd__nor2_4 _06345_ (.A(_02642_),
    .B(_02785_),
    .Y(_02796_));
 sky130_fd_sc_hd__nand2_1 _06346_ (.A(_02785_),
    .B(_02642_),
    .Y(_02807_));
 sky130_fd_sc_hd__nor2b_4 _06347_ (.A(_02796_),
    .B_N(_02807_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand3_2 _06348_ (.A(_02598_),
    .B(_02763_),
    .C(_02818_),
    .Y(_02829_));
 sky130_fd_sc_hd__o21ai_2 _06349_ (.A1(_02796_),
    .A2(_02576_),
    .B1(_02807_),
    .Y(_02840_));
 sky130_fd_sc_hd__nand2_1 _06350_ (.A(_02840_),
    .B(_02763_),
    .Y(_02851_));
 sky130_fd_sc_hd__nand3_2 _06351_ (.A(_02829_),
    .B(_02741_),
    .C(_02851_),
    .Y(_02862_));
 sky130_fd_sc_hd__buf_6 _06352_ (.A(_02862_),
    .X(_02873_));
 sky130_fd_sc_hd__xor2_1 _06353_ (.A(_02270_),
    .B(_02291_),
    .X(_02884_));
 sky130_fd_sc_hd__inv_2 _06354_ (.A(_02884_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_1 _06355_ (.A(_02873_),
    .B(_02895_),
    .Y(_02906_));
 sky130_fd_sc_hd__a21oi_1 _06356_ (.A1(_02840_),
    .A2(_02763_),
    .B1(_02752_),
    .Y(_02917_));
 sky130_fd_sc_hd__nand3_2 _06357_ (.A(_02917_),
    .B(_02270_),
    .C(net100),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_2 _06358_ (.A(_02906_),
    .B(_02928_),
    .Y(_02939_));
 sky130_fd_sc_hd__nand2_1 _06359_ (.A(_02939_),
    .B(net107),
    .Y(_02950_));
 sky130_fd_sc_hd__inv_2 _06360_ (.A(net107),
    .Y(_02961_));
 sky130_fd_sc_hd__nand3_1 _06361_ (.A(_02906_),
    .B(_02928_),
    .C(_02961_),
    .Y(_02972_));
 sky130_fd_sc_hd__inv_2 _06362_ (.A(_02291_),
    .Y(_02983_));
 sky130_fd_sc_hd__inv_4 _06363_ (.A(_02862_),
    .Y(_02994_));
 sky130_fd_sc_hd__nor2_1 _06364_ (.A(_02983_),
    .B(_02994_),
    .Y(_03005_));
 sky130_fd_sc_hd__clkinvlp_2 _06365_ (.A(_03005_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand3_1 _06366_ (.A(_02950_),
    .B(_02972_),
    .C(_03015_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand2_1 _06367_ (.A(_02939_),
    .B(_02961_),
    .Y(_03037_));
 sky130_fd_sc_hd__nand3_1 _06368_ (.A(_02906_),
    .B(_02928_),
    .C(net107),
    .Y(_03048_));
 sky130_fd_sc_hd__nand3_1 _06369_ (.A(_03037_),
    .B(_03048_),
    .C(_03005_),
    .Y(_03059_));
 sky130_fd_sc_hd__nand2_1 _06370_ (.A(net5),
    .B(_00707_),
    .Y(_03070_));
 sky130_fd_sc_hd__inv_2 _06371_ (.A(_03070_),
    .Y(_03081_));
 sky130_fd_sc_hd__and2_1 _06372_ (.A(_00685_),
    .B(net4),
    .X(_03092_));
 sky130_fd_sc_hd__or2_1 _06373_ (.A(_03081_),
    .B(_03092_),
    .X(_03103_));
 sky130_fd_sc_hd__buf_6 _06374_ (.A(_03103_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_1 _06375_ (.A0(net5),
    .A1(net6),
    .S(_00707_),
    .X(_03125_));
 sky130_fd_sc_hd__or2_1 _06376_ (.A(_03114_),
    .B(_03125_),
    .X(_03136_));
 sky130_fd_sc_hd__nor2_1 _06377_ (.A(_02291_),
    .B(_03136_),
    .Y(_03147_));
 sky130_fd_sc_hd__inv_2 _06378_ (.A(_03147_),
    .Y(_03158_));
 sky130_fd_sc_hd__nand3_1 _06379_ (.A(_03026_),
    .B(_03059_),
    .C(_03158_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand2_1 _06380_ (.A(_03169_),
    .B(_03026_),
    .Y(_03180_));
 sky130_fd_sc_hd__or2_1 _06381_ (.A(_01353_),
    .B(_02961_),
    .X(_03191_));
 sky130_fd_sc_hd__nand2_1 _06382_ (.A(_03191_),
    .B(_02259_),
    .Y(_03201_));
 sky130_fd_sc_hd__nand2_1 _06383_ (.A(_02994_),
    .B(_03201_),
    .Y(_03212_));
 sky130_fd_sc_hd__xor2_1 _06384_ (.A(_01353_),
    .B(_02302_),
    .X(_03223_));
 sky130_fd_sc_hd__nand2_1 _06385_ (.A(_02873_),
    .B(_03223_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_2 _06386_ (.A(_03212_),
    .B(_03234_),
    .Y(_03245_));
 sky130_fd_sc_hd__buf_6 _06387_ (.A(_01727_),
    .X(_03256_));
 sky130_fd_sc_hd__nand2_1 _06388_ (.A(_03245_),
    .B(_03256_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand3_2 _06389_ (.A(_03212_),
    .B(net108),
    .C(_03234_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand2_1 _06390_ (.A(_03267_),
    .B(_03278_),
    .Y(_03289_));
 sky130_fd_sc_hd__inv_2 _06391_ (.A(_02939_),
    .Y(_03300_));
 sky130_fd_sc_hd__nand3_1 _06392_ (.A(_03289_),
    .B(net107),
    .C(_03300_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand3_1 _06393_ (.A(_03267_),
    .B(_03278_),
    .C(_03048_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _06394_ (.A(_03311_),
    .B(_03322_),
    .Y(_03333_));
 sky130_fd_sc_hd__nand2_1 _06395_ (.A(_03180_),
    .B(_03333_),
    .Y(_03344_));
 sky130_fd_sc_hd__nand2_1 _06396_ (.A(_03289_),
    .B(_03048_),
    .Y(_03355_));
 sky130_fd_sc_hd__nand2_1 _06397_ (.A(_03344_),
    .B(_03355_),
    .Y(_03365_));
 sky130_fd_sc_hd__inv_2 _06398_ (.A(_02598_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _06399_ (.A(_02587_),
    .B(_02379_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_1 _06400_ (.A(_03376_),
    .B(_03387_),
    .Y(_03398_));
 sky130_fd_sc_hd__inv_4 _06401_ (.A(_03398_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand2_1 _06402_ (.A(_02994_),
    .B(_02774_),
    .Y(_03420_));
 sky130_fd_sc_hd__o21ai_2 _06403_ (.A1(_03409_),
    .A2(_02994_),
    .B1(_03420_),
    .Y(_03431_));
 sky130_fd_sc_hd__inv_2 _06404_ (.A(_03431_),
    .Y(_03442_));
 sky130_fd_sc_hd__nand2_1 _06405_ (.A(_03376_),
    .B(_02576_),
    .Y(_03453_));
 sky130_fd_sc_hd__and2_1 _06406_ (.A(_03453_),
    .B(_02818_),
    .X(_03464_));
 sky130_fd_sc_hd__o21ai_1 _06407_ (.A1(_02818_),
    .A2(_03453_),
    .B1(_02873_),
    .Y(_03475_));
 sky130_fd_sc_hd__o22ai_1 _06408_ (.A1(_02642_),
    .A2(_02873_),
    .B1(_03464_),
    .B2(_03475_),
    .Y(_03486_));
 sky130_fd_sc_hd__or2_1 _06409_ (.A(_03442_),
    .B(_03486_),
    .X(_03497_));
 sky130_fd_sc_hd__nand2_1 _06410_ (.A(_03486_),
    .B(_03442_),
    .Y(_03507_));
 sky130_fd_sc_hd__nand2_1 _06411_ (.A(_03497_),
    .B(_03507_),
    .Y(_03518_));
 sky130_fd_sc_hd__a21oi_1 _06412_ (.A1(_02248_),
    .A2(_02357_),
    .B1(_02346_),
    .Y(_03529_));
 sky130_fd_sc_hd__o21ai_1 _06413_ (.A1(_02379_),
    .A2(_03529_),
    .B1(_02873_),
    .Y(_03540_));
 sky130_fd_sc_hd__nand3_1 _06414_ (.A(_02917_),
    .B(_02237_),
    .C(net100),
    .Y(_03551_));
 sky130_fd_sc_hd__nand3_2 _06415_ (.A(_03540_),
    .B(_03551_),
    .C(_01408_),
    .Y(_03562_));
 sky130_fd_sc_hd__nor2_1 _06416_ (.A(_03431_),
    .B(_03562_),
    .Y(_03573_));
 sky130_fd_sc_hd__nand2_2 _06417_ (.A(_03562_),
    .B(_03431_),
    .Y(_03584_));
 sky130_fd_sc_hd__inv_2 _06418_ (.A(_03584_),
    .Y(_03595_));
 sky130_fd_sc_hd__nor2_1 _06419_ (.A(_03573_),
    .B(_03595_),
    .Y(_03606_));
 sky130_fd_sc_hd__nand3b_4 _06420_ (.A_N(_03529_),
    .B(net111),
    .C(_02368_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand3b_1 _06421_ (.A_N(_02237_),
    .B(_02917_),
    .C(net100),
    .Y(_03628_));
 sky130_fd_sc_hd__nand3_2 _06422_ (.A(_03617_),
    .B(_03628_),
    .C(_01408_),
    .Y(_03639_));
 sky130_fd_sc_hd__buf_6 _06423_ (.A(_01760_),
    .X(_03650_));
 sky130_fd_sc_hd__nand3_1 _06424_ (.A(_03540_),
    .B(_03551_),
    .C(_03650_),
    .Y(_03661_));
 sky130_fd_sc_hd__nand3_2 _06425_ (.A(_03639_),
    .B(_03278_),
    .C(_03661_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_1 _06426_ (.A(_03639_),
    .B(_03661_),
    .Y(_03683_));
 sky130_fd_sc_hd__inv_2 _06427_ (.A(_03278_),
    .Y(_03694_));
 sky130_fd_sc_hd__nand2_1 _06428_ (.A(_03683_),
    .B(_03694_),
    .Y(_03705_));
 sky130_fd_sc_hd__nand3_1 _06429_ (.A(_03606_),
    .B(_03672_),
    .C(_03705_),
    .Y(_03716_));
 sky130_fd_sc_hd__nor2_1 _06430_ (.A(_03518_),
    .B(_03716_),
    .Y(_03727_));
 sky130_fd_sc_hd__nand2_2 _06431_ (.A(_03727_),
    .B(_03365_),
    .Y(_03738_));
 sky130_fd_sc_hd__o21ai_2 _06432_ (.A1(_03573_),
    .A2(_03672_),
    .B1(_03584_),
    .Y(_03749_));
 sky130_fd_sc_hd__a21boi_4 _06433_ (.A1(_03749_),
    .A2(_03497_),
    .B1_N(_03507_),
    .Y(_03760_));
 sky130_fd_sc_hd__nand2_4 _06434_ (.A(_03738_),
    .B(_03760_),
    .Y(_03771_));
 sky130_fd_sc_hd__buf_8 _06435_ (.A(_03771_),
    .X(_03782_));
 sky130_fd_sc_hd__a21o_1 _06436_ (.A1(_03026_),
    .A2(_03059_),
    .B1(_03158_),
    .X(_03793_));
 sky130_fd_sc_hd__nand2_1 _06437_ (.A(_03793_),
    .B(_03169_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand2_1 _06438_ (.A(_03782_),
    .B(_03804_),
    .Y(_03815_));
 sky130_fd_sc_hd__nand3_1 _06439_ (.A(_03738_),
    .B(_03760_),
    .C(_03300_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand3_1 _06440_ (.A(_03815_),
    .B(net109),
    .C(_03826_),
    .Y(_03837_));
 sky130_fd_sc_hd__clkinvlp_2 _06441_ (.A(_03804_),
    .Y(_03848_));
 sky130_fd_sc_hd__nand2_1 _06442_ (.A(net94),
    .B(_03848_),
    .Y(_03859_));
 sky130_fd_sc_hd__nand3_1 _06443_ (.A(_03738_),
    .B(_03760_),
    .C(_02939_),
    .Y(_03869_));
 sky130_fd_sc_hd__nand3_2 _06444_ (.A(_03859_),
    .B(_03256_),
    .C(_03869_),
    .Y(_03880_));
 sky130_fd_sc_hd__nand2_1 _06445_ (.A(_03837_),
    .B(_03880_),
    .Y(_03891_));
 sky130_fd_sc_hd__and2_1 _06446_ (.A(_03136_),
    .B(_02291_),
    .X(_03902_));
 sky130_fd_sc_hd__nor2_1 _06447_ (.A(_03147_),
    .B(_03902_),
    .Y(_03913_));
 sky130_fd_sc_hd__inv_2 _06448_ (.A(_03913_),
    .Y(_03924_));
 sky130_fd_sc_hd__nand2_1 _06449_ (.A(_03771_),
    .B(_03924_),
    .Y(_03935_));
 sky130_fd_sc_hd__buf_6 _06450_ (.A(net107),
    .X(_03946_));
 sky130_fd_sc_hd__xor2_1 _06451_ (.A(_02291_),
    .B(net111),
    .X(_03957_));
 sky130_fd_sc_hd__nand3_1 _06452_ (.A(_03738_),
    .B(_03760_),
    .C(_03957_),
    .Y(_03968_));
 sky130_fd_sc_hd__nand3_1 _06453_ (.A(_03935_),
    .B(_03946_),
    .C(_03968_),
    .Y(_03979_));
 sky130_fd_sc_hd__inv_2 _06454_ (.A(_03979_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand2_1 _06455_ (.A(_03891_),
    .B(_03990_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand3_2 _06456_ (.A(_03979_),
    .B(_03837_),
    .C(_03880_),
    .Y(_04012_));
 sky130_fd_sc_hd__nand2_2 _06457_ (.A(_04001_),
    .B(_04012_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2_1 _06458_ (.A(_03935_),
    .B(_03968_),
    .Y(_04034_));
 sky130_fd_sc_hd__nand2_1 _06459_ (.A(_04034_),
    .B(_03946_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand3_1 _06460_ (.A(_03935_),
    .B(_02961_),
    .C(_03968_),
    .Y(_04056_));
 sky130_fd_sc_hd__nand2_1 _06461_ (.A(_04045_),
    .B(_04056_),
    .Y(_04067_));
 sky130_fd_sc_hd__xor2_1 _06462_ (.A(_03114_),
    .B(_03125_),
    .X(_04078_));
 sky130_fd_sc_hd__inv_2 _06463_ (.A(_04078_),
    .Y(_04089_));
 sky130_fd_sc_hd__nand2_1 _06464_ (.A(_03771_),
    .B(_04089_),
    .Y(_04100_));
 sky130_fd_sc_hd__nand3_2 _06465_ (.A(net116),
    .B(_03760_),
    .C(_03125_),
    .Y(_04111_));
 sky130_fd_sc_hd__nand3_2 _06466_ (.A(_04100_),
    .B(net111),
    .C(_04111_),
    .Y(_04122_));
 sky130_fd_sc_hd__inv_2 _06467_ (.A(_04122_),
    .Y(_04133_));
 sky130_fd_sc_hd__nand2_1 _06468_ (.A(_04067_),
    .B(_04133_),
    .Y(_04144_));
 sky130_fd_sc_hd__nand3_2 _06469_ (.A(_04045_),
    .B(_04122_),
    .C(_04056_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand2_1 _06470_ (.A(_04144_),
    .B(_04155_),
    .Y(_04166_));
 sky130_fd_sc_hd__nor2_2 _06471_ (.A(_04023_),
    .B(_04166_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_2 _06472_ (.A(_04100_),
    .B(_04111_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _06473_ (.A(_04188_),
    .B(net111),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _06474_ (.A(net94),
    .B(_03114_),
    .Y(_04210_));
 sky130_fd_sc_hd__buf_6 _06475_ (.A(_02994_),
    .X(_04220_));
 sky130_fd_sc_hd__nand3_1 _06476_ (.A(_04100_),
    .B(_04220_),
    .C(_04111_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand3_1 _06477_ (.A(_04199_),
    .B(_04210_),
    .C(_04231_),
    .Y(_04242_));
 sky130_fd_sc_hd__nand2_1 _06478_ (.A(_04188_),
    .B(_04220_),
    .Y(_04253_));
 sky130_fd_sc_hd__inv_2 _06479_ (.A(_04210_),
    .Y(_04264_));
 sky130_fd_sc_hd__nand3_1 _06480_ (.A(_04253_),
    .B(_04122_),
    .C(_04264_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand2_1 _06481_ (.A(_04242_),
    .B(_04275_),
    .Y(_04286_));
 sky130_fd_sc_hd__nor2_1 _06482_ (.A(_03114_),
    .B(_04286_),
    .Y(_04297_));
 sky130_fd_sc_hd__mux2_1 _06483_ (.A0(net2),
    .A1(net3),
    .S(_00707_),
    .X(_04308_));
 sky130_fd_sc_hd__buf_6 _06484_ (.A(_04308_),
    .X(_04319_));
 sky130_fd_sc_hd__mux2_4 _06485_ (.A0(net32),
    .A1(net2),
    .S(_00707_),
    .X(_04330_));
 sky130_fd_sc_hd__mux2_2 _06486_ (.A0(net3),
    .A1(net4),
    .S(_00707_),
    .X(_04341_));
 sky130_fd_sc_hd__mux2_1 _06487_ (.A0(net31),
    .A1(net32),
    .S(_00707_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_4 _06488_ (.A(_04352_),
    .X(_04363_));
 sky130_fd_sc_hd__mux2_4 _06489_ (.A0(net30),
    .A1(net31),
    .S(_00718_),
    .X(_04374_));
 sky130_fd_sc_hd__inv_2 _06490_ (.A(_04330_),
    .Y(_04385_));
 sky130_fd_sc_hd__inv_2 _06491_ (.A(_04319_),
    .Y(_04396_));
 sky130_fd_sc_hd__nand2_1 _06492_ (.A(_04396_),
    .B(_04330_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand2_1 _06493_ (.A(_04385_),
    .B(_04319_),
    .Y(_04418_));
 sky130_fd_sc_hd__a21oi_1 _06494_ (.A1(_04407_),
    .A2(_04418_),
    .B1(_04341_),
    .Y(_04429_));
 sky130_fd_sc_hd__o211a_1 _06495_ (.A1(_04363_),
    .A2(_04374_),
    .B1(_04385_),
    .C1(_04429_),
    .X(_04440_));
 sky130_fd_sc_hd__a211o_1 _06496_ (.A1(_04319_),
    .A2(_04330_),
    .B1(_04341_),
    .C1(_04440_),
    .X(_04451_));
 sky130_fd_sc_hd__nand3_1 _06497_ (.A(_04177_),
    .B(_04297_),
    .C(_04451_),
    .Y(_04462_));
 sky130_fd_sc_hd__o21a_1 _06498_ (.A1(_04155_),
    .A2(_04023_),
    .B1(_04012_),
    .X(_04473_));
 sky130_fd_sc_hd__inv_6 _06499_ (.A(_03771_),
    .Y(_04484_));
 sky130_fd_sc_hd__a22o_1 _06500_ (.A1(_03114_),
    .A2(_04484_),
    .B1(_04199_),
    .B2(_04231_),
    .X(_04495_));
 sky130_fd_sc_hd__nand2_1 _06501_ (.A(_04177_),
    .B(_04495_),
    .Y(_04506_));
 sky130_fd_sc_hd__nand3_1 _06502_ (.A(_04462_),
    .B(_04473_),
    .C(_04506_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand2_1 _06503_ (.A(_03705_),
    .B(_03672_),
    .Y(_04528_));
 sky130_fd_sc_hd__a21o_1 _06504_ (.A1(_03344_),
    .A2(_03355_),
    .B1(_04528_),
    .X(_04539_));
 sky130_fd_sc_hd__a21bo_1 _06505_ (.A1(_04539_),
    .A2(_03672_),
    .B1_N(_03606_),
    .X(_04550_));
 sky130_fd_sc_hd__nand3b_1 _06506_ (.A_N(_03606_),
    .B(_04539_),
    .C(_03672_),
    .Y(_04561_));
 sky130_fd_sc_hd__nand3_1 _06507_ (.A(_04550_),
    .B(_04561_),
    .C(_03782_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand2_1 _06508_ (.A(_04484_),
    .B(_03442_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _06509_ (.A(_04572_),
    .B(_04583_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2b_1 _06510_ (.A_N(_03365_),
    .B(_04528_),
    .Y(_04605_));
 sky130_fd_sc_hd__nand2_1 _06511_ (.A(_04605_),
    .B(_04539_),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _06512_ (.A(_04616_),
    .B(net94),
    .Y(_04627_));
 sky130_fd_sc_hd__nand2_1 _06513_ (.A(_03617_),
    .B(_03628_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand2_1 _06514_ (.A(_04484_),
    .B(_04638_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_2 _06515_ (.A(_04627_),
    .B(_04649_),
    .Y(_04660_));
 sky130_fd_sc_hd__inv_2 _06516_ (.A(_04660_),
    .Y(_04670_));
 sky130_fd_sc_hd__nand2_1 _06517_ (.A(_04594_),
    .B(_04670_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand3_2 _06518_ (.A(_04572_),
    .B(_04583_),
    .C(_04660_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand2_1 _06519_ (.A(_04681_),
    .B(_04692_),
    .Y(_04703_));
 sky130_fd_sc_hd__nand3_1 _06520_ (.A(_03859_),
    .B(net109),
    .C(_03869_),
    .Y(_04714_));
 sky130_fd_sc_hd__or2_1 _06521_ (.A(_03333_),
    .B(_03180_),
    .X(_04725_));
 sky130_fd_sc_hd__nand2_1 _06522_ (.A(_04725_),
    .B(_03344_),
    .Y(_04736_));
 sky130_fd_sc_hd__nand2_1 _06523_ (.A(_03771_),
    .B(_04736_),
    .Y(_04747_));
 sky130_fd_sc_hd__o21ai_4 _06524_ (.A1(_03245_),
    .A2(net94),
    .B1(_04747_),
    .Y(_04758_));
 sky130_fd_sc_hd__inv_2 _06525_ (.A(_04758_),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_1 _06526_ (.A(_04769_),
    .B(_03650_),
    .Y(_04780_));
 sky130_fd_sc_hd__buf_6 _06527_ (.A(_01408_),
    .X(_04791_));
 sky130_fd_sc_hd__nand2_2 _06528_ (.A(_04758_),
    .B(_04791_),
    .Y(_04802_));
 sky130_fd_sc_hd__nand3b_1 _06529_ (.A_N(_04714_),
    .B(_04780_),
    .C(_04802_),
    .Y(_04813_));
 sky130_fd_sc_hd__nand3_1 _06530_ (.A(_04660_),
    .B(_04791_),
    .C(_04758_),
    .Y(_04824_));
 sky130_fd_sc_hd__nand2_1 _06531_ (.A(_04670_),
    .B(_04802_),
    .Y(_04835_));
 sky130_fd_sc_hd__nand2_1 _06532_ (.A(_04824_),
    .B(_04835_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_1 _06533_ (.A(_04769_),
    .B(_04791_),
    .Y(_04857_));
 sky130_fd_sc_hd__nand2_1 _06534_ (.A(_04758_),
    .B(_03650_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand3_2 _06535_ (.A(_04857_),
    .B(_04714_),
    .C(_04868_),
    .Y(_04879_));
 sky130_fd_sc_hd__nand3_1 _06536_ (.A(_04813_),
    .B(_04846_),
    .C(_04879_),
    .Y(_04890_));
 sky130_fd_sc_hd__nor2_2 _06537_ (.A(_04703_),
    .B(_04890_),
    .Y(_04901_));
 sky130_fd_sc_hd__nand2_1 _06538_ (.A(_04517_),
    .B(_04901_),
    .Y(_04912_));
 sky130_fd_sc_hd__nor2_1 _06539_ (.A(_04660_),
    .B(_04802_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _06540_ (.A(_04802_),
    .B(_04660_),
    .Y(_04934_));
 sky130_fd_sc_hd__o21ai_1 _06541_ (.A1(_04923_),
    .A2(_04879_),
    .B1(_04934_),
    .Y(_04945_));
 sky130_fd_sc_hd__a21boi_4 _06542_ (.A1(_04945_),
    .A2(_04692_),
    .B1_N(_04681_),
    .Y(_04956_));
 sky130_fd_sc_hd__nand2_1 _06543_ (.A(_04385_),
    .B(_04363_),
    .Y(_04967_));
 sky130_fd_sc_hd__inv_2 _06544_ (.A(_04363_),
    .Y(_04978_));
 sky130_fd_sc_hd__nand2_1 _06545_ (.A(_04978_),
    .B(_04330_),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_1 _06546_ (.A(_04967_),
    .B(_04989_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _06547_ (.A(_04978_),
    .B(_04374_),
    .Y(_05011_));
 sky130_fd_sc_hd__inv_2 _06548_ (.A(_04374_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand2_1 _06549_ (.A(_05022_),
    .B(_04363_),
    .Y(_05033_));
 sky130_fd_sc_hd__nand2_1 _06550_ (.A(_05011_),
    .B(_05033_),
    .Y(_05044_));
 sky130_fd_sc_hd__or3b_1 _06551_ (.A(_05000_),
    .B(_05044_),
    .C_N(_04429_),
    .X(_05055_));
 sky130_fd_sc_hd__nand2_1 _06552_ (.A(_04177_),
    .B(_04297_),
    .Y(_05066_));
 sky130_fd_sc_hd__nor2_1 _06553_ (.A(_05055_),
    .B(_05066_),
    .Y(_05077_));
 sky130_fd_sc_hd__nand3_2 _06554_ (.A(_05077_),
    .B(_05022_),
    .C(_04901_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand3_4 _06555_ (.A(_04912_),
    .B(_04956_),
    .C(_05088_),
    .Y(_05098_));
 sky130_fd_sc_hd__inv_4 _06556_ (.A(_05098_),
    .Y(_05109_));
 sky130_fd_sc_hd__buf_6 _06557_ (.A(_05109_),
    .X(_05119_));
 sky130_fd_sc_hd__buf_6 _06558_ (.A(_05119_),
    .X(_05130_));
 sky130_fd_sc_hd__buf_6 _06559_ (.A(_05130_),
    .X(_05140_));
 sky130_fd_sc_hd__xor2_1 _06560_ (.A(_04341_),
    .B(_04319_),
    .X(_05151_));
 sky130_fd_sc_hd__nand2_1 _06561_ (.A(_05098_),
    .B(_05151_),
    .Y(_05161_));
 sky130_fd_sc_hd__inv_2 _06562_ (.A(_04341_),
    .Y(_05172_));
 sky130_fd_sc_hd__nand2_1 _06563_ (.A(_05172_),
    .B(_04396_),
    .Y(_05183_));
 sky130_fd_sc_hd__or2_1 _06564_ (.A(_03114_),
    .B(_05183_),
    .X(_05193_));
 sky130_fd_sc_hd__nand3_1 _06565_ (.A(_04242_),
    .B(_04275_),
    .C(_05193_),
    .Y(_05204_));
 sky130_fd_sc_hd__nand2_1 _06566_ (.A(_05204_),
    .B(_04242_),
    .Y(_05214_));
 sky130_fd_sc_hd__inv_2 _06567_ (.A(_04166_),
    .Y(_05225_));
 sky130_fd_sc_hd__nand2_1 _06568_ (.A(_05214_),
    .B(_05225_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_1 _06569_ (.A(_05236_),
    .B(_04155_),
    .Y(_05246_));
 sky130_fd_sc_hd__inv_2 _06570_ (.A(_04023_),
    .Y(_05257_));
 sky130_fd_sc_hd__nand2_1 _06571_ (.A(_05246_),
    .B(_05257_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand2_1 _06572_ (.A(_05267_),
    .B(_04012_),
    .Y(_05278_));
 sky130_fd_sc_hd__nand2_2 _06573_ (.A(_05278_),
    .B(_04901_),
    .Y(_05288_));
 sky130_fd_sc_hd__nand3_1 _06574_ (.A(_05288_),
    .B(_05172_),
    .C(net99),
    .Y(_05299_));
 sky130_fd_sc_hd__nand2_2 _06575_ (.A(_05161_),
    .B(_05299_),
    .Y(_05310_));
 sky130_fd_sc_hd__nand2_2 _06576_ (.A(_05310_),
    .B(_03782_),
    .Y(_05320_));
 sky130_fd_sc_hd__nand3_1 _06577_ (.A(_05161_),
    .B(_05299_),
    .C(_04484_),
    .Y(_05331_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(_05320_),
    .B(_05331_),
    .Y(_05341_));
 sky130_fd_sc_hd__nand2_1 _06579_ (.A(_05098_),
    .B(_04319_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_1 _06580_ (.A(_05341_),
    .B(_05352_),
    .Y(_05363_));
 sky130_fd_sc_hd__inv_2 _06581_ (.A(_05352_),
    .Y(_05373_));
 sky130_fd_sc_hd__nand3_1 _06582_ (.A(_05320_),
    .B(_05331_),
    .C(_05373_),
    .Y(_05384_));
 sky130_fd_sc_hd__nand2_2 _06583_ (.A(_05363_),
    .B(_05384_),
    .Y(_05394_));
 sky130_fd_sc_hd__buf_8 _06584_ (.A(_05098_),
    .X(_05405_));
 sky130_fd_sc_hd__nand2_1 _06585_ (.A(_05183_),
    .B(_03114_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand2_1 _06586_ (.A(_05193_),
    .B(_05415_),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_2 _06587_ (.A(_05405_),
    .B(_05426_),
    .Y(_05436_));
 sky130_fd_sc_hd__xor2_1 _06588_ (.A(_03114_),
    .B(_03782_),
    .X(_05447_));
 sky130_fd_sc_hd__nand3_1 _06589_ (.A(_05288_),
    .B(_04956_),
    .C(_05447_),
    .Y(_05457_));
 sky130_fd_sc_hd__nand2_2 _06590_ (.A(_05436_),
    .B(_05457_),
    .Y(_05468_));
 sky130_fd_sc_hd__buf_8 _06591_ (.A(net111),
    .X(_05479_));
 sky130_fd_sc_hd__nand2_1 _06592_ (.A(_05468_),
    .B(_05479_),
    .Y(_05489_));
 sky130_fd_sc_hd__nand3_1 _06593_ (.A(_05436_),
    .B(_05457_),
    .C(_04220_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_1 _06594_ (.A(_05489_),
    .B(_05500_),
    .Y(_05510_));
 sky130_fd_sc_hd__inv_2 _06595_ (.A(_05320_),
    .Y(_05521_));
 sky130_fd_sc_hd__nand2_1 _06596_ (.A(_05510_),
    .B(_05521_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _06597_ (.A(_05468_),
    .B(_04220_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand3_2 _06598_ (.A(_05436_),
    .B(_05457_),
    .C(_05479_),
    .Y(_05553_));
 sky130_fd_sc_hd__nand2_1 _06599_ (.A(_05542_),
    .B(_05553_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2_1 _06600_ (.A(_05563_),
    .B(_05320_),
    .Y(_05574_));
 sky130_fd_sc_hd__nand2_1 _06601_ (.A(_05532_),
    .B(_05574_),
    .Y(_05584_));
 sky130_fd_sc_hd__nor2_1 _06602_ (.A(_05394_),
    .B(_05584_),
    .Y(_05595_));
 sky130_fd_sc_hd__nand3b_1 _06603_ (.A_N(_04034_),
    .B(_05288_),
    .C(_04956_),
    .Y(_05606_));
 sky130_fd_sc_hd__or2_1 _06604_ (.A(_05225_),
    .B(_05214_),
    .X(_05616_));
 sky130_fd_sc_hd__nand2_1 _06605_ (.A(_05616_),
    .B(_05236_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand2_1 _06606_ (.A(_05405_),
    .B(_05627_),
    .Y(_05637_));
 sky130_fd_sc_hd__buf_6 _06607_ (.A(net110),
    .X(_05648_));
 sky130_fd_sc_hd__nand3_1 _06608_ (.A(_05606_),
    .B(_05637_),
    .C(_05648_),
    .Y(_05659_));
 sky130_fd_sc_hd__inv_2 _06609_ (.A(_05627_),
    .Y(_05670_));
 sky130_fd_sc_hd__nand2_1 _06610_ (.A(_05405_),
    .B(_05670_),
    .Y(_05681_));
 sky130_fd_sc_hd__nand3_1 _06611_ (.A(_05288_),
    .B(_04956_),
    .C(_04034_),
    .Y(_05692_));
 sky130_fd_sc_hd__nand3_1 _06612_ (.A(_05681_),
    .B(_05692_),
    .C(_03256_),
    .Y(_05703_));
 sky130_fd_sc_hd__nand2_1 _06613_ (.A(_05659_),
    .B(_05703_),
    .Y(_05714_));
 sky130_fd_sc_hd__or2b_1 _06614_ (.A(_05193_),
    .B_N(_04286_),
    .X(_05725_));
 sky130_fd_sc_hd__nand2_1 _06615_ (.A(_05725_),
    .B(_05204_),
    .Y(_05736_));
 sky130_fd_sc_hd__inv_2 _06616_ (.A(_05736_),
    .Y(_05743_));
 sky130_fd_sc_hd__nand2_1 _06617_ (.A(_05098_),
    .B(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand3_2 _06618_ (.A(_05288_),
    .B(_04956_),
    .C(_04188_),
    .Y(_05745_));
 sky130_fd_sc_hd__nand3_1 _06619_ (.A(_05744_),
    .B(_05745_),
    .C(_03946_),
    .Y(_05746_));
 sky130_fd_sc_hd__inv_2 _06620_ (.A(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__nand2_1 _06621_ (.A(_05714_),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand3_2 _06622_ (.A(_05659_),
    .B(_05746_),
    .C(_05703_),
    .Y(_05749_));
 sky130_fd_sc_hd__nand2_2 _06623_ (.A(_05749_),
    .B(_05748_),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_2 _06624_ (.A(_05744_),
    .B(_05745_),
    .Y(_05751_));
 sky130_fd_sc_hd__nand2_1 _06625_ (.A(_05751_),
    .B(_03946_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand3_1 _06626_ (.A(_05744_),
    .B(_05745_),
    .C(_02961_),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2_1 _06627_ (.A(_05752_),
    .B(_05753_),
    .Y(_05754_));
 sky130_fd_sc_hd__inv_2 _06628_ (.A(_05553_),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _06629_ (.A(_05754_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__nand3_2 _06630_ (.A(_05752_),
    .B(_05553_),
    .C(_05753_),
    .Y(_05757_));
 sky130_fd_sc_hd__nand2_1 _06631_ (.A(_05756_),
    .B(_05757_),
    .Y(_05758_));
 sky130_fd_sc_hd__nor2_2 _06632_ (.A(_05758_),
    .B(_05750_),
    .Y(_05759_));
 sky130_fd_sc_hd__mux2_1 _06633_ (.A0(net29),
    .A1(net30),
    .S(_00718_),
    .X(_05760_));
 sky130_fd_sc_hd__buf_6 _06634_ (.A(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__inv_1 _06635_ (.A(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand2_1 _06636_ (.A(_05022_),
    .B(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2_1 _06637_ (.A(_05763_),
    .B(_04363_),
    .Y(_05764_));
 sky130_fd_sc_hd__or3b_1 _06638_ (.A(_04319_),
    .B(_04330_),
    .C_N(_05764_),
    .X(_05765_));
 sky130_fd_sc_hd__nand3_1 _06639_ (.A(_05595_),
    .B(_05759_),
    .C(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__nand2_1 _06640_ (.A(_05563_),
    .B(_05521_),
    .Y(_05767_));
 sky130_fd_sc_hd__nand2_1 _06641_ (.A(_05510_),
    .B(_05320_),
    .Y(_05768_));
 sky130_fd_sc_hd__nand2_1 _06642_ (.A(_05767_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__inv_2 _06643_ (.A(_05363_),
    .Y(_05770_));
 sky130_fd_sc_hd__nand2_1 _06644_ (.A(_05769_),
    .B(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _06645_ (.A(_05771_),
    .B(_05574_),
    .Y(_05772_));
 sky130_fd_sc_hd__nand2_1 _06646_ (.A(_05772_),
    .B(_05759_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21a_1 _06647_ (.A1(_05757_),
    .A2(_05750_),
    .B1(_05749_),
    .X(_05774_));
 sky130_fd_sc_hd__nand3_1 _06648_ (.A(_05766_),
    .B(_05773_),
    .C(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__or2_1 _06649_ (.A(_05257_),
    .B(_05246_),
    .X(_05776_));
 sky130_fd_sc_hd__nand3_1 _06650_ (.A(_05098_),
    .B(_05267_),
    .C(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_1 _06651_ (.A(_03859_),
    .B(_03869_),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_1 _06652_ (.A(_05109_),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_1 _06653_ (.A(_05777_),
    .B(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__inv_2 _06654_ (.A(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_2 _06655_ (.A(_05781_),
    .B(_04791_),
    .Y(_05782_));
 sky130_fd_sc_hd__nand2_1 _06656_ (.A(_04813_),
    .B(_04879_),
    .Y(_05783_));
 sky130_fd_sc_hd__inv_2 _06657_ (.A(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__or2_1 _06658_ (.A(_05784_),
    .B(_05278_),
    .X(_05785_));
 sky130_fd_sc_hd__nand2_1 _06659_ (.A(_05278_),
    .B(_05784_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand2_1 _06660_ (.A(_05785_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__nand2_1 _06661_ (.A(_05787_),
    .B(_05405_),
    .Y(_05788_));
 sky130_fd_sc_hd__nand2_1 _06662_ (.A(_05109_),
    .B(_04758_),
    .Y(_05789_));
 sky130_fd_sc_hd__nand2_1 _06663_ (.A(_05788_),
    .B(_05789_),
    .Y(_05790_));
 sky130_fd_sc_hd__inv_2 _06664_ (.A(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__nand2_1 _06665_ (.A(_05782_),
    .B(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hd__nand3_1 _06666_ (.A(_05790_),
    .B(_05781_),
    .C(_04791_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_1 _06667_ (.A(_05792_),
    .B(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__nand2_1 _06668_ (.A(_05780_),
    .B(_03650_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand2_1 _06669_ (.A(_05782_),
    .B(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__nand2_1 _06670_ (.A(_05606_),
    .B(_05637_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand2_1 _06671_ (.A(_05797_),
    .B(_05648_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_1 _06672_ (.A(_05796_),
    .B(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__nand3b_1 _06673_ (.A_N(_05798_),
    .B(_05782_),
    .C(_05795_),
    .Y(_05800_));
 sky130_fd_sc_hd__nand3_1 _06674_ (.A(_05794_),
    .B(_05799_),
    .C(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__nand2_1 _06675_ (.A(_05786_),
    .B(_04879_),
    .Y(_05802_));
 sky130_fd_sc_hd__or2_1 _06676_ (.A(_04846_),
    .B(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__nand2_1 _06677_ (.A(_05802_),
    .B(_04846_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand3_1 _06678_ (.A(_05803_),
    .B(_05804_),
    .C(_05405_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_1 _06679_ (.A1(_04660_),
    .A2(_05405_),
    .B1(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__or2_1 _06680_ (.A(_05791_),
    .B(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__nand2_1 _06681_ (.A(_05806_),
    .B(_05791_),
    .Y(_05808_));
 sky130_fd_sc_hd__nand2_1 _06682_ (.A(_05807_),
    .B(_05808_),
    .Y(_05809_));
 sky130_fd_sc_hd__nor2_2 _06683_ (.A(_05809_),
    .B(_05801_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand2_1 _06684_ (.A(_05775_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__xor2_2 _06685_ (.A(_04374_),
    .B(_05761_),
    .X(_05812_));
 sky130_fd_sc_hd__a2111o_1 _06686_ (.A1(_05011_),
    .A2(_05033_),
    .B1(_04319_),
    .C1(_04330_),
    .D1(_05812_),
    .X(_05813_));
 sky130_fd_sc_hd__nand2_1 _06687_ (.A(_05595_),
    .B(_05759_),
    .Y(_05814_));
 sky130_fd_sc_hd__nor2_1 _06688_ (.A(_05813_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__nand3_2 _06689_ (.A(_05810_),
    .B(_05815_),
    .C(_05762_),
    .Y(_05816_));
 sky130_fd_sc_hd__nor2_1 _06690_ (.A(_05790_),
    .B(_05782_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _06691_ (.A(_05782_),
    .B(_05790_),
    .Y(_05818_));
 sky130_fd_sc_hd__o21ai_1 _06692_ (.A1(_05817_),
    .A2(_05799_),
    .B1(_05818_),
    .Y(_05819_));
 sky130_fd_sc_hd__a21boi_2 _06693_ (.A1(_05819_),
    .A2(_05807_),
    .B1_N(_05808_),
    .Y(_05820_));
 sky130_fd_sc_hd__nand3_4 _06694_ (.A(_05811_),
    .B(_05816_),
    .C(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__buf_6 _06695_ (.A(_05821_),
    .X(_05822_));
 sky130_fd_sc_hd__nand2_1 _06696_ (.A(_04385_),
    .B(_04978_),
    .Y(_05823_));
 sky130_fd_sc_hd__nor2_1 _06697_ (.A(_04319_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__inv_2 _06698_ (.A(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(_05823_),
    .B(_04319_),
    .Y(_05826_));
 sky130_fd_sc_hd__nand2_1 _06700_ (.A(_05825_),
    .B(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__inv_2 _06701_ (.A(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__nand2_1 _06702_ (.A(_05822_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__inv_2 _06703_ (.A(_05394_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand3_1 _06704_ (.A(_05830_),
    .B(_05769_),
    .C(_05825_),
    .Y(_05831_));
 sky130_fd_sc_hd__a21boi_1 _06705_ (.A1(_05770_),
    .A2(_05532_),
    .B1_N(_05574_),
    .Y(_05832_));
 sky130_fd_sc_hd__nand2_1 _06706_ (.A(_05831_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__clkinvlp_2 _06707_ (.A(_05750_),
    .Y(_05834_));
 sky130_fd_sc_hd__inv_2 _06708_ (.A(_05758_),
    .Y(_05835_));
 sky130_fd_sc_hd__nand3_1 _06709_ (.A(_05833_),
    .B(_05834_),
    .C(_05835_),
    .Y(_05836_));
 sky130_fd_sc_hd__nand2_1 _06710_ (.A(_05836_),
    .B(_05774_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_4 _06711_ (.A(_05837_),
    .B(_05810_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_1 _06712_ (.A(_05109_),
    .B(_04319_),
    .Y(_05839_));
 sky130_fd_sc_hd__nand2_1 _06713_ (.A(_05405_),
    .B(_04396_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(_05839_),
    .B(_05840_),
    .Y(_05841_));
 sky130_fd_sc_hd__inv_2 _06715_ (.A(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__nand3_1 _06716_ (.A(_05838_),
    .B(net96),
    .C(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__nand3_1 _06717_ (.A(_05829_),
    .B(_05843_),
    .C(_03782_),
    .Y(_05844_));
 sky130_fd_sc_hd__nand2_1 _06718_ (.A(_05821_),
    .B(_05827_),
    .Y(_05845_));
 sky130_fd_sc_hd__nand3_1 _06719_ (.A(_05838_),
    .B(net103),
    .C(_05841_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand3_1 _06720_ (.A(_05845_),
    .B(_05846_),
    .C(_04484_),
    .Y(_05847_));
 sky130_fd_sc_hd__nand2_1 _06721_ (.A(_05844_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__inv_2 _06722_ (.A(_05000_),
    .Y(_05849_));
 sky130_fd_sc_hd__nand2_1 _06723_ (.A(_05821_),
    .B(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hd__nand3_2 _06724_ (.A(_05838_),
    .B(_04330_),
    .C(net103),
    .Y(_05851_));
 sky130_fd_sc_hd__nand3_2 _06725_ (.A(_05850_),
    .B(_05851_),
    .C(_05405_),
    .Y(_05852_));
 sky130_fd_sc_hd__inv_2 _06726_ (.A(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__nand2_1 _06727_ (.A(_05848_),
    .B(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__nand3_2 _06728_ (.A(_05852_),
    .B(_05844_),
    .C(_05847_),
    .Y(_05855_));
 sky130_fd_sc_hd__nand2_1 _06729_ (.A(_05854_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__inv_2 _06730_ (.A(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__nand2_1 _06731_ (.A(_05830_),
    .B(_05825_),
    .Y(_05858_));
 sky130_fd_sc_hd__nand2_1 _06732_ (.A(_05394_),
    .B(_05824_),
    .Y(_05859_));
 sky130_fd_sc_hd__nand2_1 _06733_ (.A(_05858_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__inv_2 _06734_ (.A(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__nand2_1 _06735_ (.A(_05821_),
    .B(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__inv_2 _06736_ (.A(_05310_),
    .Y(_05863_));
 sky130_fd_sc_hd__nand3_1 _06737_ (.A(_05838_),
    .B(net103),
    .C(_05863_),
    .Y(_05864_));
 sky130_fd_sc_hd__nand2_1 _06738_ (.A(_05862_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__nand2_1 _06739_ (.A(_05865_),
    .B(_05479_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand3_1 _06740_ (.A(_05862_),
    .B(_05864_),
    .C(_04220_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand2_1 _06741_ (.A(_05866_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__nand2_2 _06742_ (.A(_05845_),
    .B(_05846_),
    .Y(_05869_));
 sky130_fd_sc_hd__inv_2 _06743_ (.A(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__nand2_1 _06744_ (.A(_05870_),
    .B(_03782_),
    .Y(_05871_));
 sky130_fd_sc_hd__nand2_1 _06745_ (.A(_05868_),
    .B(_05871_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand3_2 _06746_ (.A(_05862_),
    .B(_05864_),
    .C(_05479_),
    .Y(_05873_));
 sky130_fd_sc_hd__nand2_1 _06747_ (.A(_05822_),
    .B(_05860_),
    .Y(_05874_));
 sky130_fd_sc_hd__nand3_1 _06748_ (.A(_05838_),
    .B(net96),
    .C(_05310_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand3_1 _06749_ (.A(_05874_),
    .B(_05875_),
    .C(_04220_),
    .Y(_05876_));
 sky130_fd_sc_hd__nand2_1 _06750_ (.A(_05873_),
    .B(_05876_),
    .Y(_05877_));
 sky130_fd_sc_hd__nor2_1 _06751_ (.A(_04484_),
    .B(_05869_),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_1 _06752_ (.A(_05877_),
    .B(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__nand2_1 _06753_ (.A(_05872_),
    .B(_05879_),
    .Y(_05880_));
 sky130_fd_sc_hd__nand2_1 _06754_ (.A(_05857_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__nand2_1 _06755_ (.A(_05858_),
    .B(_05363_),
    .Y(_05882_));
 sky130_fd_sc_hd__xor2_1 _06756_ (.A(_05584_),
    .B(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__inv_2 _06757_ (.A(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand2_1 _06758_ (.A(_05821_),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__nand3_2 _06759_ (.A(_05838_),
    .B(net103),
    .C(_05468_),
    .Y(_05886_));
 sky130_fd_sc_hd__nand2_1 _06760_ (.A(_05885_),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__nand2_1 _06761_ (.A(_05887_),
    .B(_03946_),
    .Y(_05888_));
 sky130_fd_sc_hd__nand3_1 _06762_ (.A(_05885_),
    .B(_05886_),
    .C(_02961_),
    .Y(_05889_));
 sky130_fd_sc_hd__nand2_1 _06763_ (.A(_05888_),
    .B(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__inv_2 _06764_ (.A(_05873_),
    .Y(_05891_));
 sky130_fd_sc_hd__nand2_1 _06765_ (.A(_05890_),
    .B(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__nand3_1 _06766_ (.A(_05888_),
    .B(_05873_),
    .C(_05889_),
    .Y(_05893_));
 sky130_fd_sc_hd__nand2_2 _06767_ (.A(_05892_),
    .B(_05893_),
    .Y(_05894_));
 sky130_fd_sc_hd__inv_2 _06768_ (.A(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__nand3_2 _06769_ (.A(_05885_),
    .B(_05886_),
    .C(_03946_),
    .Y(_05896_));
 sky130_fd_sc_hd__inv_2 _06770_ (.A(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__or2_1 _06771_ (.A(_05835_),
    .B(_05833_),
    .X(_05898_));
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(_05833_),
    .B(_05835_),
    .Y(_05899_));
 sky130_fd_sc_hd__nand2_1 _06773_ (.A(_05898_),
    .B(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(net115),
    .B(_05900_),
    .Y(_05901_));
 sky130_fd_sc_hd__inv_2 _06775_ (.A(_05751_),
    .Y(_05902_));
 sky130_fd_sc_hd__nand3_1 _06776_ (.A(_05838_),
    .B(net96),
    .C(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__nand3_2 _06777_ (.A(_05901_),
    .B(_05903_),
    .C(_05648_),
    .Y(_05904_));
 sky130_fd_sc_hd__clkinvlp_2 _06778_ (.A(_05900_),
    .Y(_05905_));
 sky130_fd_sc_hd__nand2_1 _06779_ (.A(_05822_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand3_1 _06780_ (.A(_05838_),
    .B(net96),
    .C(_05751_),
    .Y(_05907_));
 sky130_fd_sc_hd__nand3_1 _06781_ (.A(_05906_),
    .B(_05907_),
    .C(_03256_),
    .Y(_05908_));
 sky130_fd_sc_hd__nand3_1 _06782_ (.A(_05897_),
    .B(_05904_),
    .C(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(_05904_),
    .B(_05908_),
    .Y(_05910_));
 sky130_fd_sc_hd__nand2_1 _06784_ (.A(_05910_),
    .B(_05896_),
    .Y(_05911_));
 sky130_fd_sc_hd__nand2_1 _06785_ (.A(_05909_),
    .B(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__nand2_1 _06786_ (.A(_05895_),
    .B(_05912_),
    .Y(_05913_));
 sky130_fd_sc_hd__nor2_1 _06787_ (.A(_05881_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__mux2_1 _06788_ (.A0(net28),
    .A1(net29),
    .S(_00718_),
    .X(_05915_));
 sky130_fd_sc_hd__buf_6 _06789_ (.A(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__inv_1 _06790_ (.A(_05916_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand2_1 _06791_ (.A(_05762_),
    .B(_05916_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand2_1 _06792_ (.A(_05917_),
    .B(_05761_),
    .Y(_05919_));
 sky130_fd_sc_hd__a21o_1 _06793_ (.A1(_05918_),
    .A2(_05919_),
    .B1(_04374_),
    .X(_05920_));
 sky130_fd_sc_hd__nand2_1 _06794_ (.A(_05850_),
    .B(_05851_),
    .Y(_05921_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(_05921_),
    .B(_05405_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand3_1 _06796_ (.A(_05850_),
    .B(_05851_),
    .C(_05119_),
    .Y(_05923_));
 sky130_fd_sc_hd__nand2_1 _06797_ (.A(_05822_),
    .B(_04363_),
    .Y(_05924_));
 sky130_fd_sc_hd__inv_2 _06798_ (.A(_05924_),
    .Y(_05925_));
 sky130_fd_sc_hd__nand3_1 _06799_ (.A(_05922_),
    .B(_05923_),
    .C(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__nand2_1 _06800_ (.A(_05921_),
    .B(_05119_),
    .Y(_05927_));
 sky130_fd_sc_hd__nand3_1 _06801_ (.A(_05927_),
    .B(_05852_),
    .C(_05924_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _06802_ (.A(_05926_),
    .B(_05928_),
    .Y(_05929_));
 sky130_fd_sc_hd__nand3b_2 _06803_ (.A_N(_05920_),
    .B(_05929_),
    .C(_04978_),
    .Y(_05930_));
 sky130_fd_sc_hd__inv_2 _06804_ (.A(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__nand3_1 _06805_ (.A(_05914_),
    .B(_05917_),
    .C(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__nor2_1 _06806_ (.A(_05871_),
    .B(_05877_),
    .Y(_05933_));
 sky130_fd_sc_hd__nand2_1 _06807_ (.A(_05877_),
    .B(_05871_),
    .Y(_05934_));
 sky130_fd_sc_hd__o21ai_1 _06808_ (.A1(_05855_),
    .A2(_05933_),
    .B1(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__nand2_1 _06809_ (.A(_05910_),
    .B(_05897_),
    .Y(_05936_));
 sky130_fd_sc_hd__nand3_1 _06810_ (.A(_05896_),
    .B(_05904_),
    .C(_05908_),
    .Y(_05937_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(_05936_),
    .B(_05937_),
    .Y(_05938_));
 sky130_fd_sc_hd__nor2_2 _06812_ (.A(_05938_),
    .B(_05894_),
    .Y(_05939_));
 sky130_fd_sc_hd__nand2_1 _06813_ (.A(_05906_),
    .B(_05907_),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_1 _06814_ (.A(_05940_),
    .B(_03256_),
    .Y(_05941_));
 sky130_fd_sc_hd__nand3_1 _06815_ (.A(_05906_),
    .B(_05907_),
    .C(_05648_),
    .Y(_05942_));
 sky130_fd_sc_hd__nand2_1 _06816_ (.A(_05941_),
    .B(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__nor2_1 _06817_ (.A(_05896_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__o21ai_1 _06818_ (.A1(_05893_),
    .A2(_05944_),
    .B1(_05937_),
    .Y(_05945_));
 sky130_fd_sc_hd__a21oi_2 _06819_ (.A1(_05935_),
    .A2(_05939_),
    .B1(_05945_),
    .Y(_05946_));
 sky130_fd_sc_hd__a21o_1 _06820_ (.A1(_05761_),
    .A2(_05916_),
    .B1(_04374_),
    .X(_05947_));
 sky130_fd_sc_hd__nand3_1 _06821_ (.A(_05929_),
    .B(_04978_),
    .C(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__nand2_1 _06822_ (.A(_05922_),
    .B(_05923_),
    .Y(_05949_));
 sky130_fd_sc_hd__o21a_1 _06823_ (.A1(_04978_),
    .A2(net115),
    .B1(_05949_),
    .X(_05950_));
 sky130_fd_sc_hd__nand2_1 _06824_ (.A(_05948_),
    .B(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand2_1 _06825_ (.A(_05914_),
    .B(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__nand3_2 _06826_ (.A(_05932_),
    .B(_05946_),
    .C(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__nand2_1 _06827_ (.A(_05799_),
    .B(_05800_),
    .Y(_05954_));
 sky130_fd_sc_hd__a21o_1 _06828_ (.A1(_05836_),
    .A2(_05774_),
    .B1(_05954_),
    .X(_05955_));
 sky130_fd_sc_hd__nand2_1 _06829_ (.A(_05955_),
    .B(_05799_),
    .Y(_05956_));
 sky130_fd_sc_hd__or2_1 _06830_ (.A(_05794_),
    .B(_05956_),
    .X(_05957_));
 sky130_fd_sc_hd__nand2_1 _06831_ (.A(_05956_),
    .B(_05794_),
    .Y(_05958_));
 sky130_fd_sc_hd__nand3_1 _06832_ (.A(_05957_),
    .B(_05958_),
    .C(net115),
    .Y(_05959_));
 sky130_fd_sc_hd__inv_6 _06833_ (.A(_05821_),
    .Y(_05960_));
 sky130_fd_sc_hd__nand2_1 _06834_ (.A(_05960_),
    .B(_05791_),
    .Y(_05961_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_05959_),
    .B(_05961_),
    .Y(_05962_));
 sky130_fd_sc_hd__or2b_1 _06836_ (.A(_05837_),
    .B_N(_05954_),
    .X(_05963_));
 sky130_fd_sc_hd__nand2_1 _06837_ (.A(_05963_),
    .B(_05955_),
    .Y(_05964_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_05960_),
    .B(_05780_),
    .Y(_05965_));
 sky130_fd_sc_hd__o21ai_2 _06839_ (.A1(_05960_),
    .A2(_05964_),
    .B1(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(_05962_),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__inv_2 _06841_ (.A(_05966_),
    .Y(_05968_));
 sky130_fd_sc_hd__nand3_2 _06842_ (.A(_05959_),
    .B(_05961_),
    .C(_05968_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2_1 _06843_ (.A(_05967_),
    .B(_05969_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand3_1 _06844_ (.A(_05899_),
    .B(_05834_),
    .C(_05757_),
    .Y(_05971_));
 sky130_fd_sc_hd__a21o_1 _06845_ (.A1(_05899_),
    .A2(_05757_),
    .B1(_05834_),
    .X(_05972_));
 sky130_fd_sc_hd__nand3_1 _06846_ (.A(_05822_),
    .B(_05971_),
    .C(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand2_1 _06847_ (.A(_05960_),
    .B(_05797_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand2_1 _06848_ (.A(_05973_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__nand2_2 _06849_ (.A(_05975_),
    .B(_04791_),
    .Y(_05976_));
 sky130_fd_sc_hd__xnor2_1 _06850_ (.A(_05966_),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__inv_2 _06851_ (.A(_05975_),
    .Y(_05978_));
 sky130_fd_sc_hd__nand2_1 _06852_ (.A(_05978_),
    .B(_03650_),
    .Y(_05979_));
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(_05979_),
    .B(_05976_),
    .Y(_05980_));
 sky130_fd_sc_hd__nand2_1 _06854_ (.A(_05980_),
    .B(_05942_),
    .Y(_05981_));
 sky130_fd_sc_hd__nand3b_1 _06855_ (.A_N(_05942_),
    .B(_05979_),
    .C(_05976_),
    .Y(_05982_));
 sky130_fd_sc_hd__nand3_1 _06856_ (.A(_05977_),
    .B(_05981_),
    .C(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__nor2_2 _06857_ (.A(_05970_),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__nand2_2 _06858_ (.A(_05953_),
    .B(_05984_),
    .Y(_05985_));
 sky130_fd_sc_hd__nor2_1 _06859_ (.A(_05976_),
    .B(_05968_),
    .Y(_05986_));
 sky130_fd_sc_hd__nand2_1 _06860_ (.A(_05968_),
    .B(_05976_),
    .Y(_05987_));
 sky130_fd_sc_hd__o21ai_1 _06861_ (.A1(_05986_),
    .A2(_05981_),
    .B1(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__a21boi_4 _06862_ (.A1(_05988_),
    .A2(_05969_),
    .B1_N(_05967_),
    .Y(_05989_));
 sky130_fd_sc_hd__nand3_1 _06863_ (.A(_05985_),
    .B(_05022_),
    .C(_05989_),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(_05946_),
    .B(_05952_),
    .Y(_05991_));
 sky130_fd_sc_hd__nand2_1 _06865_ (.A(_05991_),
    .B(_05984_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(_05868_),
    .B(_05878_),
    .Y(_05993_));
 sky130_fd_sc_hd__nand2_1 _06867_ (.A(_05993_),
    .B(_05934_),
    .Y(_05994_));
 sky130_fd_sc_hd__nor2_1 _06868_ (.A(_05856_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2_1 _06869_ (.A(_05995_),
    .B(_05939_),
    .Y(_05996_));
 sky130_fd_sc_hd__nor2_1 _06870_ (.A(_05930_),
    .B(_05996_),
    .Y(_05997_));
 sky130_fd_sc_hd__nand3_2 _06871_ (.A(_05984_),
    .B(_05997_),
    .C(_05917_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand3_4 _06872_ (.A(_05992_),
    .B(_05998_),
    .C(_05989_),
    .Y(_05999_));
 sky130_fd_sc_hd__nand2_1 _06873_ (.A(_05999_),
    .B(_05812_),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2_1 _06874_ (.A(_05990_),
    .B(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__buf_8 _06875_ (.A(net115),
    .X(_06002_));
 sky130_fd_sc_hd__nand2_2 _06876_ (.A(_06001_),
    .B(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand3_1 _06877_ (.A(_05990_),
    .B(_06000_),
    .C(_05960_),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2_1 _06878_ (.A(_06003_),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__nand2_1 _06879_ (.A(net91),
    .B(_05761_),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(_06005_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__inv_2 _06881_ (.A(_06006_),
    .Y(_06008_));
 sky130_fd_sc_hd__nand3_1 _06882_ (.A(_06003_),
    .B(_06004_),
    .C(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2_1 _06883_ (.A(_06007_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__inv_2 _06884_ (.A(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__inv_2 _06885_ (.A(_06003_),
    .Y(_06012_));
 sky130_fd_sc_hd__xor2_1 _06886_ (.A(_04363_),
    .B(net115),
    .X(_06013_));
 sky130_fd_sc_hd__nand3_1 _06887_ (.A(_05985_),
    .B(_06013_),
    .C(net87),
    .Y(_06014_));
 sky130_fd_sc_hd__nor2_1 _06888_ (.A(_04363_),
    .B(_05763_),
    .Y(_06015_));
 sky130_fd_sc_hd__inv_2 _06889_ (.A(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__nand2_1 _06890_ (.A(_06016_),
    .B(_05764_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand2_1 _06891_ (.A(_05999_),
    .B(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__nand2_1 _06892_ (.A(_06014_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__buf_6 _06893_ (.A(_05405_),
    .X(_06020_));
 sky130_fd_sc_hd__nand2_1 _06894_ (.A(_06019_),
    .B(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__nand3_1 _06895_ (.A(_06014_),
    .B(_06018_),
    .C(_05119_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand3_1 _06896_ (.A(_06012_),
    .B(_06021_),
    .C(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__nand2_1 _06897_ (.A(_06021_),
    .B(_06022_),
    .Y(_06024_));
 sky130_fd_sc_hd__nand2_1 _06898_ (.A(_06024_),
    .B(_06003_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2_1 _06899_ (.A(_06023_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__nor2_1 _06900_ (.A(_05761_),
    .B(_05916_),
    .Y(_06027_));
 sky130_fd_sc_hd__inv_2 _06901_ (.A(_06027_),
    .Y(_06028_));
 sky130_fd_sc_hd__nand3_1 _06902_ (.A(_06011_),
    .B(_06026_),
    .C(_06028_),
    .Y(_06029_));
 sky130_fd_sc_hd__inv_2 _06903_ (.A(_06007_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(_06024_),
    .B(_06012_),
    .Y(_06031_));
 sky130_fd_sc_hd__nor2_1 _06905_ (.A(_06012_),
    .B(_06024_),
    .Y(_06032_));
 sky130_fd_sc_hd__a21oi_1 _06906_ (.A1(_06030_),
    .A2(_06031_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__nand2_1 _06907_ (.A(_06029_),
    .B(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__nand3b_1 _06908_ (.A_N(_05921_),
    .B(net89),
    .C(net88),
    .Y(_06035_));
 sky130_fd_sc_hd__clkbuf_8 _06909_ (.A(_05999_),
    .X(_06036_));
 sky130_fd_sc_hd__or2_1 _06910_ (.A(_06016_),
    .B(_05929_),
    .X(_06037_));
 sky130_fd_sc_hd__nand2_1 _06911_ (.A(_05929_),
    .B(_06016_),
    .Y(_06038_));
 sky130_fd_sc_hd__nand2_1 _06912_ (.A(_06037_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_1 _06913_ (.A(_06036_),
    .B(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__nand3_1 _06914_ (.A(_06035_),
    .B(_06040_),
    .C(_03782_),
    .Y(_06041_));
 sky130_fd_sc_hd__nand3_1 _06915_ (.A(net89),
    .B(_05921_),
    .C(net87),
    .Y(_06042_));
 sky130_fd_sc_hd__inv_2 _06916_ (.A(_06039_),
    .Y(_06043_));
 sky130_fd_sc_hd__nand2_1 _06917_ (.A(_05999_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__buf_6 _06918_ (.A(_04484_),
    .X(_06045_));
 sky130_fd_sc_hd__nand3_1 _06919_ (.A(_06042_),
    .B(_06044_),
    .C(_06045_),
    .Y(_06046_));
 sky130_fd_sc_hd__nand2_1 _06920_ (.A(_06041_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__nand3_1 _06921_ (.A(_06014_),
    .B(_06018_),
    .C(_06020_),
    .Y(_06048_));
 sky130_fd_sc_hd__inv_2 _06922_ (.A(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand2_1 _06923_ (.A(_06047_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand3_2 _06924_ (.A(_06041_),
    .B(_06048_),
    .C(_06046_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand2_1 _06925_ (.A(_06050_),
    .B(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__nand3_2 _06926_ (.A(_05985_),
    .B(_05869_),
    .C(net117),
    .Y(_06053_));
 sky130_fd_sc_hd__o21ai_2 _06927_ (.A1(_05925_),
    .A2(_05949_),
    .B1(_06038_),
    .Y(_06054_));
 sky130_fd_sc_hd__or2_1 _06928_ (.A(_05857_),
    .B(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__nand2_1 _06929_ (.A(_06054_),
    .B(_05857_),
    .Y(_06056_));
 sky130_fd_sc_hd__nand2_1 _06930_ (.A(_06055_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__inv_2 _06931_ (.A(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_2 _06932_ (.A(net91),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_2 _06933_ (.A(_06059_),
    .B(_06053_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _06934_ (.A(_06060_),
    .B(_05479_),
    .Y(_06061_));
 sky130_fd_sc_hd__nand3_1 _06935_ (.A(_06053_),
    .B(_06059_),
    .C(_04220_),
    .Y(_06062_));
 sky130_fd_sc_hd__nand2_1 _06936_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__nand2_2 _06937_ (.A(_06042_),
    .B(_06044_),
    .Y(_06064_));
 sky130_fd_sc_hd__nor2_1 _06938_ (.A(_06045_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_1 _06939_ (.A(_06063_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__nand3_2 _06940_ (.A(_06053_),
    .B(_06059_),
    .C(_05479_),
    .Y(_06067_));
 sky130_fd_sc_hd__nand3_1 _06941_ (.A(net89),
    .B(_05870_),
    .C(net117),
    .Y(_06068_));
 sky130_fd_sc_hd__nand2_1 _06942_ (.A(net91),
    .B(_06057_),
    .Y(_06069_));
 sky130_fd_sc_hd__nand3_1 _06943_ (.A(_06068_),
    .B(_06069_),
    .C(_04220_),
    .Y(_06070_));
 sky130_fd_sc_hd__nand2_1 _06944_ (.A(_06067_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__inv_2 _06945_ (.A(_06064_),
    .Y(_06072_));
 sky130_fd_sc_hd__nand2_1 _06946_ (.A(_06072_),
    .B(_03782_),
    .Y(_06073_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(_06071_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__nand2_1 _06948_ (.A(_06066_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__nor2_2 _06949_ (.A(_06052_),
    .B(_06075_),
    .Y(_06076_));
 sky130_fd_sc_hd__clkinvlp_2 _06950_ (.A(_05887_),
    .Y(_06077_));
 sky130_fd_sc_hd__nand3_1 _06951_ (.A(net89),
    .B(_06077_),
    .C(net117),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2_1 _06952_ (.A(_06054_),
    .B(_05995_),
    .Y(_06079_));
 sky130_fd_sc_hd__inv_2 _06953_ (.A(_05935_),
    .Y(_06080_));
 sky130_fd_sc_hd__nand2_1 _06954_ (.A(_06079_),
    .B(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__nand2_1 _06955_ (.A(_06081_),
    .B(_05895_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand3_1 _06956_ (.A(_06079_),
    .B(_05894_),
    .C(_06080_),
    .Y(_06083_));
 sky130_fd_sc_hd__nand2_1 _06957_ (.A(_06082_),
    .B(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__nand2_1 _06958_ (.A(net91),
    .B(_06084_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand3_1 _06959_ (.A(_06078_),
    .B(_06085_),
    .C(_05648_),
    .Y(_06086_));
 sky130_fd_sc_hd__nand3_1 _06960_ (.A(_05985_),
    .B(_05887_),
    .C(net117),
    .Y(_06087_));
 sky130_fd_sc_hd__clkinvlp_2 _06961_ (.A(_06084_),
    .Y(_06088_));
 sky130_fd_sc_hd__nand2_1 _06962_ (.A(net91),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__nand3_1 _06963_ (.A(_06087_),
    .B(_06089_),
    .C(_03256_),
    .Y(_06090_));
 sky130_fd_sc_hd__nand2_1 _06964_ (.A(_06086_),
    .B(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__nand3_2 _06965_ (.A(_05985_),
    .B(_05865_),
    .C(net117),
    .Y(_06092_));
 sky130_fd_sc_hd__nand2_1 _06966_ (.A(_06056_),
    .B(_05855_),
    .Y(_06093_));
 sky130_fd_sc_hd__nand2_1 _06967_ (.A(_06093_),
    .B(_05880_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand3_1 _06968_ (.A(_06056_),
    .B(_05994_),
    .C(_05855_),
    .Y(_06095_));
 sky130_fd_sc_hd__nand2_1 _06969_ (.A(_06094_),
    .B(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__inv_2 _06970_ (.A(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__nand2_1 _06971_ (.A(_05999_),
    .B(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand3_2 _06972_ (.A(_06092_),
    .B(_06098_),
    .C(_03946_),
    .Y(_06099_));
 sky130_fd_sc_hd__inv_2 _06973_ (.A(_06099_),
    .Y(_06100_));
 sky130_fd_sc_hd__nand2_1 _06974_ (.A(_06091_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__nand3_1 _06975_ (.A(_06099_),
    .B(_06086_),
    .C(_06090_),
    .Y(_06102_));
 sky130_fd_sc_hd__nand2_1 _06976_ (.A(_06101_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__nand2_1 _06977_ (.A(_06092_),
    .B(_06098_),
    .Y(_06104_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(_06104_),
    .B(_03946_),
    .Y(_06105_));
 sky130_fd_sc_hd__clkbuf_8 _06979_ (.A(_02961_),
    .X(_06106_));
 sky130_fd_sc_hd__nand3_1 _06980_ (.A(_06092_),
    .B(_06098_),
    .C(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__nand2_1 _06981_ (.A(_06105_),
    .B(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__clkinvlp_2 _06982_ (.A(_06067_),
    .Y(_06109_));
 sky130_fd_sc_hd__nand2_1 _06983_ (.A(_06108_),
    .B(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__nand3_2 _06984_ (.A(_06105_),
    .B(_06067_),
    .C(_06107_),
    .Y(_06111_));
 sky130_fd_sc_hd__nand2_1 _06985_ (.A(_06110_),
    .B(_06111_),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_2 _06986_ (.A(_06103_),
    .B(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand2_2 _06987_ (.A(_06076_),
    .B(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__inv_2 _06988_ (.A(_06114_),
    .Y(_06115_));
 sky130_fd_sc_hd__nand2_1 _06989_ (.A(_06034_),
    .B(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__nor2_1 _06990_ (.A(_06073_),
    .B(_06071_),
    .Y(_00035_));
 sky130_fd_sc_hd__o21ai_2 _06991_ (.A1(_06051_),
    .A2(_00035_),
    .B1(_06074_),
    .Y(_00036_));
 sky130_fd_sc_hd__inv_2 _06992_ (.A(_06101_),
    .Y(_00037_));
 sky130_fd_sc_hd__o21ai_1 _06993_ (.A1(_06111_),
    .A2(_00037_),
    .B1(_06102_),
    .Y(_00038_));
 sky130_fd_sc_hd__a21oi_1 _06994_ (.A1(_00036_),
    .A2(_06113_),
    .B1(_00038_),
    .Y(_00039_));
 sky130_fd_sc_hd__nand2_1 _06995_ (.A(_06116_),
    .B(_00039_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _06996_ (.A(_05981_),
    .B(_05982_),
    .Y(_00041_));
 sky130_fd_sc_hd__nand2b_1 _06997_ (.A_N(_00041_),
    .B(_05953_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand2_1 _06998_ (.A(_00042_),
    .B(_05981_),
    .Y(_00043_));
 sky130_fd_sc_hd__or2_1 _06999_ (.A(_05977_),
    .B(_00043_),
    .X(_00044_));
 sky130_fd_sc_hd__nand2_1 _07000_ (.A(_00043_),
    .B(_05977_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand2_1 _07001_ (.A(_00044_),
    .B(_00045_),
    .Y(_00046_));
 sky130_fd_sc_hd__nand2_1 _07002_ (.A(_00046_),
    .B(_06036_),
    .Y(_00047_));
 sky130_fd_sc_hd__nand2_1 _07003_ (.A(_00047_),
    .B(_05969_),
    .Y(_00048_));
 sky130_fd_sc_hd__inv_6 _07004_ (.A(_06036_),
    .Y(_00049_));
 sky130_fd_sc_hd__or2b_1 _07005_ (.A(_05953_),
    .B_N(_00041_),
    .X(_00050_));
 sky130_fd_sc_hd__nand2_1 _07006_ (.A(_00050_),
    .B(_00042_),
    .Y(_00051_));
 sky130_fd_sc_hd__nand2_1 _07007_ (.A(_00049_),
    .B(_05978_),
    .Y(_00052_));
 sky130_fd_sc_hd__o21ai_2 _07008_ (.A1(_00049_),
    .A2(_00051_),
    .B1(_00052_),
    .Y(_00053_));
 sky130_fd_sc_hd__inv_2 _07009_ (.A(_00053_),
    .Y(_00054_));
 sky130_fd_sc_hd__nand2_1 _07010_ (.A(_00048_),
    .B(_00054_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand3_1 _07011_ (.A(_00047_),
    .B(_05969_),
    .C(_00053_),
    .Y(_00056_));
 sky130_fd_sc_hd__nand2_1 _07012_ (.A(_00055_),
    .B(_00056_),
    .Y(_00057_));
 sky130_fd_sc_hd__nand2_1 _07013_ (.A(_06082_),
    .B(_05893_),
    .Y(_00058_));
 sky130_fd_sc_hd__or2_1 _07014_ (.A(_05912_),
    .B(_00058_),
    .X(_00059_));
 sky130_fd_sc_hd__nand2_1 _07015_ (.A(_00058_),
    .B(_05912_),
    .Y(_00060_));
 sky130_fd_sc_hd__nand3_1 _07016_ (.A(_00059_),
    .B(_00060_),
    .C(_06036_),
    .Y(_00061_));
 sky130_fd_sc_hd__nand2_1 _07017_ (.A(_00049_),
    .B(_05940_),
    .Y(_00062_));
 sky130_fd_sc_hd__nand2_1 _07018_ (.A(_00061_),
    .B(_00062_),
    .Y(_00063_));
 sky130_fd_sc_hd__inv_2 _07019_ (.A(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__nand3_1 _07020_ (.A(_00054_),
    .B(_04791_),
    .C(_00064_),
    .Y(_00065_));
 sky130_fd_sc_hd__nand2_1 _07021_ (.A(_00064_),
    .B(_04791_),
    .Y(_00066_));
 sky130_fd_sc_hd__nand2_1 _07022_ (.A(_00066_),
    .B(_00053_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_1 _07023_ (.A(_00065_),
    .B(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_1 _07024_ (.A(_00063_),
    .B(_04791_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand3_1 _07025_ (.A(_00061_),
    .B(_03650_),
    .C(_00062_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_1 _07026_ (.A(_00069_),
    .B(_00070_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand2_1 _07027_ (.A(_06078_),
    .B(_06085_),
    .Y(_00072_));
 sky130_fd_sc_hd__nand3_1 _07028_ (.A(_00071_),
    .B(_05648_),
    .C(_00072_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand3_1 _07029_ (.A(_06087_),
    .B(_06089_),
    .C(_05648_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand3_2 _07030_ (.A(_00069_),
    .B(_00074_),
    .C(_00070_),
    .Y(_00075_));
 sky130_fd_sc_hd__nand3_1 _07031_ (.A(_00068_),
    .B(_00073_),
    .C(_00075_),
    .Y(_00076_));
 sky130_fd_sc_hd__nor2_2 _07032_ (.A(_00076_),
    .B(_00057_),
    .Y(_00077_));
 sky130_fd_sc_hd__nand2_1 _07033_ (.A(_00040_),
    .B(_00077_),
    .Y(_00078_));
 sky130_fd_sc_hd__nor2_1 _07034_ (.A(_00054_),
    .B(_00066_),
    .Y(_00079_));
 sky130_fd_sc_hd__nand2_1 _07035_ (.A(_00066_),
    .B(_00054_),
    .Y(_00080_));
 sky130_fd_sc_hd__o21ai_1 _07036_ (.A1(_00075_),
    .A2(_00079_),
    .B1(_00080_),
    .Y(_00081_));
 sky130_fd_sc_hd__a21boi_4 _07037_ (.A1(_00081_),
    .A2(_00055_),
    .B1_N(_00056_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand3_1 _07038_ (.A(_06011_),
    .B(_06026_),
    .C(_06027_),
    .Y(_00083_));
 sky130_fd_sc_hd__nor2_2 _07039_ (.A(_00083_),
    .B(_06114_),
    .Y(_00084_));
 sky130_fd_sc_hd__mux2_1 _07040_ (.A0(net27),
    .A1(net28),
    .S(_00718_),
    .X(_00085_));
 sky130_fd_sc_hd__buf_6 _07041_ (.A(_00085_),
    .X(_00086_));
 sky130_fd_sc_hd__nand3_2 _07042_ (.A(_00077_),
    .B(_00084_),
    .C(_00086_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand3_4 _07043_ (.A(_00078_),
    .B(_00082_),
    .C(_00087_),
    .Y(_00088_));
 sky130_fd_sc_hd__buf_8 _07044_ (.A(_00088_),
    .X(_00089_));
 sky130_fd_sc_hd__inv_6 _07045_ (.A(_00089_),
    .Y(_00090_));
 sky130_fd_sc_hd__clkbuf_8 _07046_ (.A(_00090_),
    .X(_00091_));
 sky130_fd_sc_hd__buf_6 _07047_ (.A(_00091_),
    .X(_00092_));
 sky130_fd_sc_hd__nand2_1 _07048_ (.A(_00084_),
    .B(_00086_),
    .Y(_00093_));
 sky130_fd_sc_hd__nand3_1 _07049_ (.A(_00093_),
    .B(_00039_),
    .C(_06116_),
    .Y(_00094_));
 sky130_fd_sc_hd__nand2_2 _07050_ (.A(_00094_),
    .B(_00077_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand3_1 _07051_ (.A(_00095_),
    .B(_00082_),
    .C(_06064_),
    .Y(_00096_));
 sky130_fd_sc_hd__inv_2 _07052_ (.A(_06052_),
    .Y(_00097_));
 sky130_fd_sc_hd__inv_2 _07053_ (.A(_00086_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_1 _07054_ (.A(_06027_),
    .B(_00098_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand3_1 _07055_ (.A(_06007_),
    .B(_06009_),
    .C(_00099_),
    .Y(_00100_));
 sky130_fd_sc_hd__nand2_1 _07056_ (.A(_00100_),
    .B(_06007_),
    .Y(_00101_));
 sky130_fd_sc_hd__nand2_1 _07057_ (.A(_00101_),
    .B(_06026_),
    .Y(_00102_));
 sky130_fd_sc_hd__inv_2 _07058_ (.A(_06032_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_1 _07059_ (.A(_00102_),
    .B(_00103_),
    .Y(_00104_));
 sky130_fd_sc_hd__or2_1 _07060_ (.A(_00097_),
    .B(_00104_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2_1 _07061_ (.A(_00104_),
    .B(_00097_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_1 _07062_ (.A(_00105_),
    .B(_00106_),
    .Y(_00107_));
 sky130_fd_sc_hd__inv_2 _07063_ (.A(_00107_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_1 _07064_ (.A(_00088_),
    .B(_00108_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand3_2 _07065_ (.A(_00096_),
    .B(_00109_),
    .C(_05479_),
    .Y(_00110_));
 sky130_fd_sc_hd__buf_6 _07066_ (.A(_00095_),
    .X(_00111_));
 sky130_fd_sc_hd__buf_6 _07067_ (.A(_00082_),
    .X(_00112_));
 sky130_fd_sc_hd__nand3_1 _07068_ (.A(_00111_),
    .B(_00112_),
    .C(_06072_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_1 _07069_ (.A(_00089_),
    .B(_00107_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand3_2 _07070_ (.A(_00113_),
    .B(_00114_),
    .C(_04220_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_2 _07071_ (.A(_00115_),
    .B(_00110_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand3_1 _07072_ (.A(_00111_),
    .B(_00112_),
    .C(_06019_),
    .Y(_00117_));
 sky130_fd_sc_hd__or2_1 _07073_ (.A(_06026_),
    .B(_00101_),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_1 _07074_ (.A(_00118_),
    .B(_00102_),
    .Y(_00119_));
 sky130_fd_sc_hd__inv_2 _07075_ (.A(_00119_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_2 _07076_ (.A(net106),
    .B(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand3_4 _07077_ (.A(_00117_),
    .B(_00121_),
    .C(_03782_),
    .Y(_00122_));
 sky130_fd_sc_hd__inv_2 _07078_ (.A(_00122_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _07079_ (.A(_00116_),
    .B(_00123_),
    .Y(_00124_));
 sky130_fd_sc_hd__nand3_1 _07080_ (.A(_00110_),
    .B(_00122_),
    .C(_00115_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _07081_ (.A(_00124_),
    .B(_00125_),
    .Y(_00126_));
 sky130_fd_sc_hd__inv_2 _07082_ (.A(_06019_),
    .Y(_00127_));
 sky130_fd_sc_hd__nand3_1 _07083_ (.A(_00111_),
    .B(_00112_),
    .C(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _07084_ (.A(_00089_),
    .B(_00119_),
    .Y(_00129_));
 sky130_fd_sc_hd__nand3_1 _07085_ (.A(_00128_),
    .B(_00129_),
    .C(_06045_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _07086_ (.A(_00122_),
    .B(_00130_),
    .Y(_00131_));
 sky130_fd_sc_hd__inv_2 _07087_ (.A(_06001_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand3_2 _07088_ (.A(_00111_),
    .B(_00112_),
    .C(_00132_),
    .Y(_00133_));
 sky130_fd_sc_hd__or2_1 _07089_ (.A(_00099_),
    .B(_06011_),
    .X(_00134_));
 sky130_fd_sc_hd__nand2_1 _07090_ (.A(_00134_),
    .B(_00100_),
    .Y(_00135_));
 sky130_fd_sc_hd__inv_2 _07091_ (.A(_00135_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand2_2 _07092_ (.A(net106),
    .B(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__nand3_2 _07093_ (.A(_00133_),
    .B(_00137_),
    .C(_06020_),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2_2 _07094_ (.A(_00131_),
    .B(_00138_),
    .Y(_00139_));
 sky130_fd_sc_hd__nand3b_1 _07095_ (.A_N(_00138_),
    .B(_00122_),
    .C(_00130_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand3_1 _07096_ (.A(_00126_),
    .B(_00139_),
    .C(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__nand3b_1 _07097_ (.A_N(_06104_),
    .B(_00111_),
    .C(_00112_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand2_1 _07098_ (.A(_00104_),
    .B(_06076_),
    .Y(_00143_));
 sky130_fd_sc_hd__inv_2 _07099_ (.A(_00036_),
    .Y(_00144_));
 sky130_fd_sc_hd__nand2_1 _07100_ (.A(_00143_),
    .B(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _07101_ (.A(_06112_),
    .Y(_00146_));
 sky130_fd_sc_hd__nand2_1 _07102_ (.A(_00145_),
    .B(_00146_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand3_1 _07103_ (.A(_00143_),
    .B(_06112_),
    .C(_00144_),
    .Y(_00148_));
 sky130_fd_sc_hd__nand2_1 _07104_ (.A(_00147_),
    .B(_00148_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand2_1 _07105_ (.A(_00089_),
    .B(_00149_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand3_1 _07106_ (.A(_00142_),
    .B(_05648_),
    .C(_00150_),
    .Y(_00151_));
 sky130_fd_sc_hd__clkinvlp_2 _07107_ (.A(_00149_),
    .Y(_00152_));
 sky130_fd_sc_hd__nand2_2 _07108_ (.A(_00152_),
    .B(_00088_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand3_2 _07109_ (.A(_00111_),
    .B(_00112_),
    .C(_06104_),
    .Y(_00154_));
 sky130_fd_sc_hd__nand3_1 _07110_ (.A(_00153_),
    .B(_00154_),
    .C(_03256_),
    .Y(_00155_));
 sky130_fd_sc_hd__nand2_1 _07111_ (.A(_00151_),
    .B(_00155_),
    .Y(_00156_));
 sky130_fd_sc_hd__nand2_1 _07112_ (.A(_00106_),
    .B(_06051_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand2_1 _07113_ (.A(_06063_),
    .B(_06073_),
    .Y(_00158_));
 sky130_fd_sc_hd__nand2_1 _07114_ (.A(_06071_),
    .B(_06065_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(_00158_),
    .B(_00159_),
    .Y(_00160_));
 sky130_fd_sc_hd__nand2_1 _07116_ (.A(_00157_),
    .B(_00160_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand3_1 _07117_ (.A(_00106_),
    .B(_06075_),
    .C(_06051_),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _07118_ (.A(_00161_),
    .B(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__inv_2 _07119_ (.A(_00163_),
    .Y(_00164_));
 sky130_fd_sc_hd__nand2_1 _07120_ (.A(_00164_),
    .B(_00088_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand3_2 _07121_ (.A(_00111_),
    .B(_00112_),
    .C(_06060_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand3_1 _07122_ (.A(_00165_),
    .B(_00166_),
    .C(_03946_),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _07123_ (.A(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _07124_ (.A(_00156_),
    .B(_00168_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand3_1 _07125_ (.A(_00167_),
    .B(_00151_),
    .C(_00155_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_2 _07126_ (.A(_00169_),
    .B(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _07127_ (.A(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__nand3_1 _07128_ (.A(_00165_),
    .B(_00166_),
    .C(_06106_),
    .Y(_00173_));
 sky130_fd_sc_hd__inv_2 _07129_ (.A(_06060_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand3_1 _07130_ (.A(_00111_),
    .B(_00112_),
    .C(_00174_),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _07131_ (.A(net106),
    .B(_00163_),
    .Y(_00176_));
 sky130_fd_sc_hd__clkbuf_8 _07132_ (.A(_03946_),
    .X(_00177_));
 sky130_fd_sc_hd__nand3_2 _07133_ (.A(_00175_),
    .B(_00176_),
    .C(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _07134_ (.A(_00173_),
    .B(_00178_),
    .Y(_00179_));
 sky130_fd_sc_hd__inv_2 _07135_ (.A(_00110_),
    .Y(_00180_));
 sky130_fd_sc_hd__nand2_1 _07136_ (.A(_00179_),
    .B(_00180_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand3_2 _07137_ (.A(_00173_),
    .B(_00110_),
    .C(_00178_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_2 _07138_ (.A(_00181_),
    .B(_00182_),
    .Y(_00183_));
 sky130_fd_sc_hd__inv_2 _07139_ (.A(_00183_),
    .Y(_00184_));
 sky130_fd_sc_hd__nand2_1 _07140_ (.A(_00172_),
    .B(_00184_),
    .Y(_00185_));
 sky130_fd_sc_hd__nor2_2 _07141_ (.A(_00141_),
    .B(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _07142_ (.A(_00089_),
    .B(_00086_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand3_2 _07143_ (.A(_00095_),
    .B(_05916_),
    .C(_00082_),
    .Y(_00188_));
 sky130_fd_sc_hd__xor2_1 _07144_ (.A(_05916_),
    .B(_00086_),
    .X(_00189_));
 sky130_fd_sc_hd__inv_2 _07145_ (.A(_00189_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_2 _07146_ (.A(_00088_),
    .B(_00190_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_2 _07147_ (.A(_00188_),
    .B(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _07148_ (.A(_00192_),
    .B(_06036_),
    .Y(_00193_));
 sky130_fd_sc_hd__buf_6 _07149_ (.A(_00049_),
    .X(_00194_));
 sky130_fd_sc_hd__nand3_1 _07150_ (.A(_00188_),
    .B(_00191_),
    .C(_00194_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand3b_1 _07151_ (.A_N(_00187_),
    .B(_00193_),
    .C(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _07152_ (.A(_00192_),
    .B(_00194_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand3_4 _07153_ (.A(_00188_),
    .B(_00191_),
    .C(_06036_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand3_1 _07154_ (.A(_00197_),
    .B(_00198_),
    .C(_00187_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _07155_ (.A(_00196_),
    .B(_00199_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _07156_ (.A(_00200_),
    .B(_00098_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _07157_ (.A(_00049_),
    .B(_05761_),
    .Y(_00202_));
 sky130_fd_sc_hd__nand2_1 _07158_ (.A(_06036_),
    .B(_05762_),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _07159_ (.A(_00202_),
    .B(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__inv_2 _07160_ (.A(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand3_1 _07161_ (.A(_00111_),
    .B(_00112_),
    .C(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__o21ai_1 _07162_ (.A1(_05916_),
    .A2(_00086_),
    .B1(_05761_),
    .Y(_00207_));
 sky130_fd_sc_hd__and2_1 _07163_ (.A(_00207_),
    .B(_00099_),
    .X(_00208_));
 sky130_fd_sc_hd__nand2_1 _07164_ (.A(_00089_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand3_2 _07165_ (.A(_00206_),
    .B(_00209_),
    .C(_06002_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand3_1 _07166_ (.A(_00111_),
    .B(_00112_),
    .C(_00204_),
    .Y(_00211_));
 sky130_fd_sc_hd__inv_2 _07167_ (.A(_00208_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _07168_ (.A(net106),
    .B(_00212_),
    .Y(_00213_));
 sky130_fd_sc_hd__buf_6 _07169_ (.A(_05960_),
    .X(_00214_));
 sky130_fd_sc_hd__nand3_2 _07170_ (.A(_00211_),
    .B(_00213_),
    .C(_00214_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _07171_ (.A(_00210_),
    .B(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _07172_ (.A(_00198_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _07173_ (.A(_00216_),
    .B(_00217_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand3_4 _07174_ (.A(_00198_),
    .B(_00210_),
    .C(_00215_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _07175_ (.A(_00218_),
    .B(_00219_),
    .Y(_00220_));
 sky130_fd_sc_hd__inv_2 _07176_ (.A(_00220_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_2 _07177_ (.A(_00133_),
    .B(_00137_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _07178_ (.A(_00222_),
    .B(_06020_),
    .Y(_00223_));
 sky130_fd_sc_hd__nand3_1 _07179_ (.A(_00133_),
    .B(_00137_),
    .C(_05119_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_1 _07180_ (.A(_00223_),
    .B(_00224_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_2 _07181_ (.A(_00211_),
    .B(_00213_),
    .Y(_00226_));
 sky130_fd_sc_hd__nor2_4 _07182_ (.A(_00214_),
    .B(_00226_),
    .Y(_00227_));
 sky130_fd_sc_hd__inv_2 _07183_ (.A(_00227_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _07184_ (.A(_00225_),
    .B(_00228_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _07185_ (.A(_00222_),
    .B(_05119_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _07186_ (.A(_00230_),
    .B(_00138_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _07187_ (.A(_00231_),
    .B(_00227_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _07188_ (.A(_00229_),
    .B(_00232_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(_00221_),
    .B(_00233_),
    .Y(_00234_));
 sky130_fd_sc_hd__nor2_1 _07190_ (.A(_00201_),
    .B(_00234_),
    .Y(_00235_));
 sky130_fd_sc_hd__mux2_1 _07191_ (.A0(net23),
    .A1(net26),
    .S(_00718_),
    .X(_00236_));
 sky130_fd_sc_hd__buf_6 _07192_ (.A(_00236_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_2 _07193_ (.A0(net26),
    .A1(net27),
    .S(_00718_),
    .X(_00238_));
 sky130_fd_sc_hd__nor2_1 _07194_ (.A(_00237_),
    .B(_00238_),
    .Y(_00239_));
 sky130_fd_sc_hd__clkinvlp_2 _07195_ (.A(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand3_1 _07196_ (.A(_00186_),
    .B(_00235_),
    .C(_00240_),
    .Y(_00241_));
 sky130_fd_sc_hd__nor2_1 _07197_ (.A(_00122_),
    .B(_00116_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _07198_ (.A(_00116_),
    .B(_00122_),
    .Y(_00243_));
 sky130_fd_sc_hd__o21ai_2 _07199_ (.A1(_00139_),
    .A2(_00242_),
    .B1(_00243_),
    .Y(_00244_));
 sky130_fd_sc_hd__nor2_2 _07200_ (.A(_00183_),
    .B(_00171_),
    .Y(_00245_));
 sky130_fd_sc_hd__inv_2 _07201_ (.A(_00169_),
    .Y(_00246_));
 sky130_fd_sc_hd__o21ai_1 _07202_ (.A1(_00182_),
    .A2(_00246_),
    .B1(_00170_),
    .Y(_00247_));
 sky130_fd_sc_hd__a21oi_2 _07203_ (.A1(_00244_),
    .A2(_00245_),
    .B1(_00247_),
    .Y(_00248_));
 sky130_fd_sc_hd__buf_6 _07204_ (.A(_00089_),
    .X(_00249_));
 sky130_fd_sc_hd__o211ai_1 _07205_ (.A1(_00098_),
    .A2(_00249_),
    .B1(_00198_),
    .C1(_00197_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand3_1 _07206_ (.A(_00221_),
    .B(_00233_),
    .C(_00250_),
    .Y(_00251_));
 sky130_fd_sc_hd__inv_2 _07207_ (.A(_00219_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _07208_ (.A(_00225_),
    .B(_00227_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _07209_ (.A(_00231_),
    .B(_00228_),
    .Y(_00254_));
 sky130_fd_sc_hd__a21boi_1 _07210_ (.A1(_00252_),
    .A2(_00253_),
    .B1_N(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _07211_ (.A(_00251_),
    .B(_00255_),
    .Y(_00256_));
 sky130_fd_sc_hd__nand2_1 _07212_ (.A(_00186_),
    .B(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand3_2 _07213_ (.A(_00241_),
    .B(_00248_),
    .C(_00257_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _07214_ (.A(_00073_),
    .B(_00075_),
    .Y(_00259_));
 sky130_fd_sc_hd__or2b_4 _07215_ (.A(_00259_),
    .B_N(_00094_),
    .X(_00260_));
 sky130_fd_sc_hd__a21bo_1 _07216_ (.A1(_00260_),
    .A2(_00075_),
    .B1_N(_00068_),
    .X(_00261_));
 sky130_fd_sc_hd__nand3b_1 _07217_ (.A_N(_00068_),
    .B(_00260_),
    .C(_00075_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand3_1 _07218_ (.A(_00261_),
    .B(_00262_),
    .C(_00249_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _07219_ (.A(_00090_),
    .B(_00053_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _07220_ (.A(_00263_),
    .B(_00264_),
    .Y(_00265_));
 sky130_fd_sc_hd__or2b_1 _07221_ (.A(_00094_),
    .B_N(_00259_),
    .X(_00266_));
 sky130_fd_sc_hd__nand2_1 _07222_ (.A(_00266_),
    .B(_00260_),
    .Y(_00267_));
 sky130_fd_sc_hd__nand2_1 _07223_ (.A(_00267_),
    .B(_00089_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _07224_ (.A(_00090_),
    .B(_00064_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_2 _07225_ (.A(_00268_),
    .B(_00269_),
    .Y(_00270_));
 sky130_fd_sc_hd__inv_2 _07226_ (.A(_00270_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _07227_ (.A(_00265_),
    .B(_00271_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand3_1 _07228_ (.A(_00263_),
    .B(_00264_),
    .C(_00270_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _07229_ (.A(_00272_),
    .B(_00273_),
    .Y(_00274_));
 sky130_fd_sc_hd__nor2_1 _07230_ (.A(_06099_),
    .B(_06091_),
    .Y(_00275_));
 sky130_fd_sc_hd__and2_1 _07231_ (.A(_06091_),
    .B(_06099_),
    .X(_00276_));
 sky130_fd_sc_hd__o211ai_2 _07232_ (.A1(_00275_),
    .A2(_00276_),
    .B1(_06111_),
    .C1(_00147_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _07233_ (.A(_00147_),
    .B(_06111_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(_00278_),
    .B(_06103_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand3_2 _07235_ (.A(_00277_),
    .B(_00089_),
    .C(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _07236_ (.A(_00090_),
    .B(_00072_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_2 _07237_ (.A(_00280_),
    .B(_00281_),
    .Y(_00282_));
 sky130_fd_sc_hd__buf_6 _07238_ (.A(_04791_),
    .X(_00283_));
 sky130_fd_sc_hd__nand2_2 _07239_ (.A(_00282_),
    .B(_00283_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _07240_ (.A(_00284_),
    .B(_00271_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand3_1 _07241_ (.A(_00282_),
    .B(_00270_),
    .C(_00283_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(_00285_),
    .B(_00286_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand3_1 _07243_ (.A(_00280_),
    .B(_03650_),
    .C(_00281_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand2_1 _07244_ (.A(_00284_),
    .B(_00288_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand3_1 _07245_ (.A(_00153_),
    .B(_00154_),
    .C(_05648_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_2 _07246_ (.A(_00289_),
    .B(_00290_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand3b_1 _07247_ (.A_N(_00290_),
    .B(_00284_),
    .C(_00288_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand3_1 _07248_ (.A(_00287_),
    .B(_00291_),
    .C(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__nor2_2 _07249_ (.A(_00274_),
    .B(_00293_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_4 _07250_ (.A(_00258_),
    .B(_00294_),
    .Y(_00295_));
 sky130_fd_sc_hd__nor2_1 _07251_ (.A(_00270_),
    .B(_00284_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _07252_ (.A(_00284_),
    .B(_00270_),
    .Y(_00297_));
 sky130_fd_sc_hd__o21ai_1 _07253_ (.A1(_00296_),
    .A2(_00291_),
    .B1(_00297_),
    .Y(_00298_));
 sky130_fd_sc_hd__a21boi_2 _07254_ (.A1(_00298_),
    .A2(_00273_),
    .B1_N(_00272_),
    .Y(_00299_));
 sky130_fd_sc_hd__clkbuf_4 _07255_ (.A(_00299_),
    .X(_00300_));
 sky130_fd_sc_hd__nand3_2 _07256_ (.A(_00295_),
    .B(_00300_),
    .C(_00238_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _07257_ (.A(_00257_),
    .B(_00248_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _07258_ (.A(_00302_),
    .B(_00294_),
    .Y(_00303_));
 sky130_fd_sc_hd__inv_2 _07259_ (.A(_00201_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(_00254_),
    .B(_00253_),
    .Y(_00305_));
 sky130_fd_sc_hd__nor2_1 _07261_ (.A(_00220_),
    .B(_00305_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _07262_ (.A(_00304_),
    .B(_00306_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand3_1 _07263_ (.A(_00123_),
    .B(_00110_),
    .C(_00115_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _07264_ (.A(_00308_),
    .B(_00243_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand2_1 _07265_ (.A(_00140_),
    .B(_00139_),
    .Y(_00310_));
 sky130_fd_sc_hd__nor2_2 _07266_ (.A(_00309_),
    .B(_00310_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(_00311_),
    .B(_00245_),
    .Y(_00312_));
 sky130_fd_sc_hd__nor2_1 _07268_ (.A(_00307_),
    .B(_00312_),
    .Y(_00313_));
 sky130_fd_sc_hd__nand3_2 _07269_ (.A(_00313_),
    .B(_00294_),
    .C(_00240_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand3_4 _07270_ (.A(_00303_),
    .B(_00299_),
    .C(_00314_),
    .Y(_00315_));
 sky130_fd_sc_hd__buf_6 _07271_ (.A(_00315_),
    .X(_00316_));
 sky130_fd_sc_hd__nand2_1 _07272_ (.A(_00237_),
    .B(_00238_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _07273_ (.A(_00240_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_2 _07274_ (.A(_00316_),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_2 _07275_ (.A(_00319_),
    .B(_00301_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _07276_ (.A(_00320_),
    .B(_00249_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand3_1 _07277_ (.A(_00301_),
    .B(_00319_),
    .C(_00090_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _07278_ (.A(_00316_),
    .B(_00237_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand3_2 _07279_ (.A(_00321_),
    .B(_00322_),
    .C(_00323_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand3_2 _07280_ (.A(_00301_),
    .B(_00319_),
    .C(_00249_),
    .Y(_00326_));
 sky130_fd_sc_hd__nor2_1 _07281_ (.A(_00098_),
    .B(_00089_),
    .Y(_00327_));
 sky130_fd_sc_hd__clkinvlp_2 _07282_ (.A(_00327_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _07283_ (.A(_00249_),
    .B(_00098_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _07284_ (.A(_00328_),
    .B(_00329_),
    .Y(_00330_));
 sky130_fd_sc_hd__nand3_2 _07285_ (.A(net122),
    .B(_00300_),
    .C(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__nor2_1 _07286_ (.A(_00086_),
    .B(_00239_),
    .Y(_00332_));
 sky130_fd_sc_hd__inv_2 _07287_ (.A(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _07288_ (.A(_00239_),
    .B(_00086_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _07289_ (.A(_00333_),
    .B(_00334_),
    .Y(_00335_));
 sky130_fd_sc_hd__inv_2 _07290_ (.A(_00335_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_2 _07291_ (.A(_00316_),
    .B(_00337_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand3_4 _07292_ (.A(_00331_),
    .B(_00338_),
    .C(_06036_),
    .Y(_00339_));
 sky130_fd_sc_hd__clkinvlp_2 _07293_ (.A(_00330_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand3_1 _07294_ (.A(net122),
    .B(_00300_),
    .C(_00340_),
    .Y(_00341_));
 sky130_fd_sc_hd__buf_6 _07295_ (.A(_00315_),
    .X(_00342_));
 sky130_fd_sc_hd__nand2_1 _07296_ (.A(_00342_),
    .B(_00335_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand3_1 _07297_ (.A(_00341_),
    .B(_00343_),
    .C(_00194_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_2 _07298_ (.A(_00339_),
    .B(_00344_),
    .Y(_00345_));
 sky130_fd_sc_hd__nor2_2 _07299_ (.A(_00326_),
    .B(_00345_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _07300_ (.A(_00345_),
    .B(_00326_),
    .Y(_00348_));
 sky130_fd_sc_hd__o21ai_2 _07301_ (.A1(_00324_),
    .A2(_00346_),
    .B1(_00348_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand3_2 _07302_ (.A(_00295_),
    .B(_00300_),
    .C(_00192_),
    .Y(_00350_));
 sky130_fd_sc_hd__nor2_1 _07303_ (.A(_00332_),
    .B(_00327_),
    .Y(_00351_));
 sky130_fd_sc_hd__a21o_1 _07304_ (.A1(_00197_),
    .A2(_00198_),
    .B1(_00351_),
    .X(_00352_));
 sky130_fd_sc_hd__nand3_2 _07305_ (.A(_00197_),
    .B(_00198_),
    .C(_00351_),
    .Y(_00353_));
 sky130_fd_sc_hd__nand2_1 _07306_ (.A(_00352_),
    .B(_00353_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_2 _07307_ (.A(_00316_),
    .B(_00354_),
    .Y(_00355_));
 sky130_fd_sc_hd__nand2_2 _07308_ (.A(_00355_),
    .B(_00350_),
    .Y(_00356_));
 sky130_fd_sc_hd__nor2_2 _07309_ (.A(_00214_),
    .B(_00356_),
    .Y(_00357_));
 sky130_fd_sc_hd__nand3_1 _07310_ (.A(_00295_),
    .B(_00300_),
    .C(_00226_),
    .Y(_00359_));
 sky130_fd_sc_hd__or2_1 _07311_ (.A(_00353_),
    .B(_00221_),
    .X(_00360_));
 sky130_fd_sc_hd__nand3_1 _07312_ (.A(_00218_),
    .B(_00219_),
    .C(_00353_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_1 _07313_ (.A(_00360_),
    .B(_00361_),
    .Y(_00362_));
 sky130_fd_sc_hd__inv_2 _07314_ (.A(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_2 _07315_ (.A(_00316_),
    .B(_00363_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand3_4 _07316_ (.A(_00359_),
    .B(_00364_),
    .C(_06020_),
    .Y(_00365_));
 sky130_fd_sc_hd__nand3b_1 _07317_ (.A_N(_00226_),
    .B(net122),
    .C(_00300_),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _07318_ (.A(_00342_),
    .B(_00362_),
    .Y(_00367_));
 sky130_fd_sc_hd__nand3_1 _07319_ (.A(_00366_),
    .B(_00367_),
    .C(_05119_),
    .Y(_00368_));
 sky130_fd_sc_hd__nand3_2 _07320_ (.A(_00357_),
    .B(_00365_),
    .C(_00368_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand3_1 _07321_ (.A(_00366_),
    .B(_00367_),
    .C(_06020_),
    .Y(_00371_));
 sky130_fd_sc_hd__nand3_2 _07322_ (.A(_00350_),
    .B(_00355_),
    .C(_06002_),
    .Y(_00372_));
 sky130_fd_sc_hd__nand3_1 _07323_ (.A(_00359_),
    .B(_00364_),
    .C(_05119_),
    .Y(_00373_));
 sky130_fd_sc_hd__nand3_1 _07324_ (.A(_00371_),
    .B(_00372_),
    .C(_00373_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_2 _07325_ (.A(_00370_),
    .B(_00374_),
    .Y(_00375_));
 sky130_fd_sc_hd__inv_2 _07326_ (.A(_00339_),
    .Y(_00376_));
 sky130_fd_sc_hd__nand3b_1 _07327_ (.A_N(_00192_),
    .B(_00295_),
    .C(_00300_),
    .Y(_00377_));
 sky130_fd_sc_hd__inv_2 _07328_ (.A(_00354_),
    .Y(_00378_));
 sky130_fd_sc_hd__nand2_1 _07329_ (.A(_00342_),
    .B(_00378_),
    .Y(_00379_));
 sky130_fd_sc_hd__nand3_1 _07330_ (.A(_00377_),
    .B(_00379_),
    .C(_00214_),
    .Y(_00381_));
 sky130_fd_sc_hd__nand3_1 _07331_ (.A(_00376_),
    .B(_00372_),
    .C(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__nand2_1 _07332_ (.A(_00381_),
    .B(_00372_),
    .Y(_00383_));
 sky130_fd_sc_hd__nand2_2 _07333_ (.A(_00383_),
    .B(_00339_),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_2 _07334_ (.A(_00382_),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__nor2_4 _07335_ (.A(_00375_),
    .B(_00385_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _07336_ (.A(_00349_),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__inv_2 _07337_ (.A(_00384_),
    .Y(_00388_));
 sky130_fd_sc_hd__a21boi_2 _07338_ (.A1(_00388_),
    .A2(_00370_),
    .B1_N(_00374_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _07339_ (.A(_00387_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _07340_ (.A(_00096_),
    .B(_00109_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand3b_1 _07341_ (.A_N(_00392_),
    .B(net122),
    .C(_00300_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _07342_ (.A(_00361_),
    .B(_00219_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(_00394_),
    .B(_00233_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_2 _07344_ (.A(_00395_),
    .B(_00254_),
    .Y(_00396_));
 sky130_fd_sc_hd__inv_2 _07345_ (.A(_00310_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _07346_ (.A(_00396_),
    .B(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _07347_ (.A(_00398_),
    .B(_00139_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _07348_ (.A(_00399_),
    .B(_00126_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand3_1 _07349_ (.A(_00398_),
    .B(_00309_),
    .C(_00139_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _07350_ (.A(_00400_),
    .B(_00401_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _07351_ (.A(_00316_),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__nand3_1 _07352_ (.A(_00393_),
    .B(_00177_),
    .C(_00404_),
    .Y(_00405_));
 sky130_fd_sc_hd__inv_2 _07353_ (.A(_00403_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _07354_ (.A(_00406_),
    .B(_00316_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand3_2 _07355_ (.A(net122),
    .B(_00300_),
    .C(_00392_),
    .Y(_00408_));
 sky130_fd_sc_hd__nand3_1 _07356_ (.A(_00407_),
    .B(_00408_),
    .C(_06106_),
    .Y(_00409_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(_00405_),
    .B(_00409_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _07358_ (.A(_00117_),
    .B(_00121_),
    .Y(_00411_));
 sky130_fd_sc_hd__nand3_1 _07359_ (.A(_00295_),
    .B(_00300_),
    .C(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__or2_1 _07360_ (.A(_00397_),
    .B(_00396_),
    .X(_00414_));
 sky130_fd_sc_hd__nand2_1 _07361_ (.A(_00414_),
    .B(_00398_),
    .Y(_00415_));
 sky130_fd_sc_hd__inv_2 _07362_ (.A(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__nand2_1 _07363_ (.A(_00315_),
    .B(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand3_2 _07364_ (.A(_00412_),
    .B(_00417_),
    .C(_05479_),
    .Y(_00418_));
 sky130_fd_sc_hd__inv_2 _07365_ (.A(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _07366_ (.A(_00410_),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand3_2 _07367_ (.A(_00405_),
    .B(_00409_),
    .C(_00418_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_2 _07368_ (.A(_00420_),
    .B(_00421_),
    .Y(_00422_));
 sky130_fd_sc_hd__inv_2 _07369_ (.A(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__clkinv_4 _07370_ (.A(_00315_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _07371_ (.A(_00165_),
    .B(_00166_),
    .Y(_00426_));
 sky130_fd_sc_hd__nand2_1 _07372_ (.A(_00425_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _07373_ (.A(_00396_),
    .B(_00311_),
    .Y(_00428_));
 sky130_fd_sc_hd__inv_2 _07374_ (.A(_00244_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _07375_ (.A(_00428_),
    .B(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(_00430_),
    .B(_00184_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand3_1 _07377_ (.A(_00428_),
    .B(_00429_),
    .C(_00183_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _07378_ (.A(_00431_),
    .B(_00432_),
    .Y(_00433_));
 sky130_fd_sc_hd__clkinvlp_2 _07379_ (.A(_00433_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _07380_ (.A(_00434_),
    .B(_00342_),
    .Y(_00436_));
 sky130_fd_sc_hd__buf_6 _07381_ (.A(_05648_),
    .X(_00437_));
 sky130_fd_sc_hd__nand3_2 _07382_ (.A(_00427_),
    .B(_00436_),
    .C(_00437_),
    .Y(_00438_));
 sky130_fd_sc_hd__inv_2 _07383_ (.A(_00426_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _07384_ (.A(_00425_),
    .B(_00439_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _07385_ (.A(_00342_),
    .B(_00433_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand3_1 _07386_ (.A(_00440_),
    .B(_00441_),
    .C(_03256_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_2 _07387_ (.A(_00438_),
    .B(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand3_2 _07388_ (.A(_00407_),
    .B(_00408_),
    .C(_00177_),
    .Y(_00444_));
 sky130_fd_sc_hd__inv_2 _07389_ (.A(_00444_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _07390_ (.A(_00443_),
    .B(_00445_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand3_1 _07391_ (.A(_00427_),
    .B(_00436_),
    .C(_03256_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand3_1 _07392_ (.A(_00440_),
    .B(_00441_),
    .C(_00437_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _07393_ (.A(_00448_),
    .B(_00449_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _07394_ (.A(_00450_),
    .B(_00444_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(_00447_),
    .B(_00451_),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _07396_ (.A(_00423_),
    .B(_00452_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(_00412_),
    .B(_00417_),
    .Y(_00454_));
 sky130_fd_sc_hd__buf_8 _07398_ (.A(_04220_),
    .X(_00455_));
 sky130_fd_sc_hd__nand2_1 _07399_ (.A(_00454_),
    .B(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _07400_ (.A(_00456_),
    .B(_00418_),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _07401_ (.A(_00425_),
    .B(_00222_),
    .Y(_00459_));
 sky130_fd_sc_hd__clkbuf_8 _07402_ (.A(_03782_),
    .X(_00460_));
 sky130_fd_sc_hd__or2_1 _07403_ (.A(_00233_),
    .B(_00394_),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _07404_ (.A(_00461_),
    .B(_00395_),
    .X(_00462_));
 sky130_fd_sc_hd__nand2_2 _07405_ (.A(_00316_),
    .B(_00462_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand3_4 _07406_ (.A(_00459_),
    .B(_00460_),
    .C(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__inv_2 _07407_ (.A(_00464_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(_00458_),
    .B(_00465_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand3_1 _07409_ (.A(_00464_),
    .B(_00456_),
    .C(_00418_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _07410_ (.A(_00466_),
    .B(_00467_),
    .Y(_00469_));
 sky130_fd_sc_hd__clkinvlp_2 _07411_ (.A(_00222_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _07412_ (.A(_00425_),
    .B(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__inv_2 _07413_ (.A(_00462_),
    .Y(_00472_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(_00342_),
    .B(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand3_1 _07415_ (.A(_00471_),
    .B(_06045_),
    .C(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _07416_ (.A(_00464_),
    .B(_00474_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_4 _07417_ (.A(_00475_),
    .B(_00365_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand3b_1 _07418_ (.A_N(_00365_),
    .B(_00464_),
    .C(_00474_),
    .Y(_00477_));
 sky130_fd_sc_hd__nand3_1 _07419_ (.A(_00469_),
    .B(_00476_),
    .C(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__nor2_2 _07420_ (.A(_00453_),
    .B(_00478_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_2 _07421_ (.A(_00390_),
    .B(_00480_),
    .Y(_00481_));
 sky130_fd_sc_hd__inv_2 _07422_ (.A(_00476_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _07423_ (.A(_00469_),
    .B(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _07424_ (.A(_00458_),
    .B(_00464_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _07425_ (.A(_00483_),
    .B(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(_00443_),
    .B(_00444_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _07427_ (.A(_00450_),
    .B(_00445_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _07428_ (.A(_00486_),
    .B(_00487_),
    .Y(_00488_));
 sky130_fd_sc_hd__nor2_2 _07429_ (.A(_00422_),
    .B(_00488_),
    .Y(_00489_));
 sky130_fd_sc_hd__nor2_1 _07430_ (.A(_00444_),
    .B(_00443_),
    .Y(_00491_));
 sky130_fd_sc_hd__o21ai_1 _07431_ (.A1(_00421_),
    .A2(_00491_),
    .B1(_00486_),
    .Y(_00492_));
 sky130_fd_sc_hd__a21oi_2 _07432_ (.A1(_00485_),
    .A2(_00489_),
    .B1(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _07433_ (.A(_00481_),
    .B(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__a21o_1 _07434_ (.A1(_00431_),
    .A2(_00182_),
    .B1(_00171_),
    .X(_00495_));
 sky130_fd_sc_hd__nand3_1 _07435_ (.A(_00431_),
    .B(_00171_),
    .C(_00182_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand3_1 _07436_ (.A(_00495_),
    .B(_00316_),
    .C(_00496_),
    .Y(_00497_));
 sky130_fd_sc_hd__a21o_1 _07437_ (.A1(_00154_),
    .A2(_00153_),
    .B1(_00316_),
    .X(_00498_));
 sky130_fd_sc_hd__nand2_1 _07438_ (.A(_00497_),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__inv_2 _07439_ (.A(_00499_),
    .Y(_00500_));
 sky130_fd_sc_hd__inv_2 _07440_ (.A(_00282_),
    .Y(_00502_));
 sky130_fd_sc_hd__a21o_1 _07441_ (.A1(_00291_),
    .A2(_00292_),
    .B1(_00258_),
    .X(_00503_));
 sky130_fd_sc_hd__nand3_1 _07442_ (.A(_00258_),
    .B(_00291_),
    .C(_00292_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _07443_ (.A(_00503_),
    .B(_00504_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _07444_ (.A(_00505_),
    .B(_00342_),
    .Y(_00506_));
 sky130_fd_sc_hd__o21ai_2 _07445_ (.A1(_00502_),
    .A2(_00342_),
    .B1(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand3_1 _07446_ (.A(_00500_),
    .B(_00283_),
    .C(_00507_),
    .Y(_00508_));
 sky130_fd_sc_hd__inv_2 _07447_ (.A(_00507_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand3_1 _07448_ (.A(_00497_),
    .B(_00283_),
    .C(_00498_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _07449_ (.A(_00509_),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _07450_ (.A(_00508_),
    .B(_00511_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(_00499_),
    .B(_00283_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand3_1 _07452_ (.A(_00497_),
    .B(_03650_),
    .C(_00498_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _07453_ (.A(_00514_),
    .B(_00515_),
    .Y(_00516_));
 sky130_fd_sc_hd__inv_2 _07454_ (.A(_00438_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _07455_ (.A(_00516_),
    .B(_00517_),
    .Y(_00518_));
 sky130_fd_sc_hd__nand3_2 _07456_ (.A(_00514_),
    .B(_00438_),
    .C(_00515_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand3_1 _07457_ (.A(_00513_),
    .B(_00518_),
    .C(_00519_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _07458_ (.A(_00504_),
    .B(_00291_),
    .Y(_00521_));
 sky130_fd_sc_hd__or2_1 _07459_ (.A(_00287_),
    .B(_00521_),
    .X(_00522_));
 sky130_fd_sc_hd__nand2_1 _07460_ (.A(_00521_),
    .B(_00287_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand3_1 _07461_ (.A(_00522_),
    .B(_00524_),
    .C(_00342_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _07462_ (.A(_00425_),
    .B(_00271_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _07463_ (.A(_00525_),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__or2_1 _07464_ (.A(_00509_),
    .B(_00527_),
    .X(_00528_));
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(_00527_),
    .B(_00509_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _07466_ (.A(_00528_),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__nor2_2 _07467_ (.A(_00520_),
    .B(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _07468_ (.A(_00494_),
    .B(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__inv_2 _07469_ (.A(_00519_),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2_1 _07470_ (.A(_00513_),
    .B(_00533_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _07471_ (.A(_00510_),
    .B(_00507_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _07472_ (.A(_00535_),
    .B(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__a21boi_4 _07473_ (.A1(_00537_),
    .A2(_00528_),
    .B1_N(_00529_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _07474_ (.A(_00320_),
    .B(_00091_),
    .Y(_00539_));
 sky130_fd_sc_hd__inv_2 _07475_ (.A(_00323_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand3_1 _07476_ (.A(_00539_),
    .B(_00326_),
    .C(_00540_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_2 _07477_ (.A(_00324_),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_2 _07478_ (.A(_00331_),
    .B(_00338_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _07479_ (.A(_00543_),
    .B(_06036_),
    .Y(_00544_));
 sky130_fd_sc_hd__nand3_1 _07480_ (.A(_00331_),
    .B(_00338_),
    .C(_00194_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _07481_ (.A(_00544_),
    .B(_00546_),
    .Y(_00547_));
 sky130_fd_sc_hd__inv_2 _07482_ (.A(_00326_),
    .Y(_00548_));
 sky130_fd_sc_hd__nand2_1 _07483_ (.A(_00547_),
    .B(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _07484_ (.A(_00549_),
    .B(_00348_),
    .Y(_00550_));
 sky130_fd_sc_hd__nor2_2 _07485_ (.A(_00542_),
    .B(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _07486_ (.A(_00386_),
    .B(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand3_1 _07487_ (.A(_00465_),
    .B(_00418_),
    .C(_00456_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_1 _07488_ (.A(_00553_),
    .B(_00484_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _07489_ (.A(_00477_),
    .B(_00476_),
    .Y(_00555_));
 sky130_fd_sc_hd__nor2_1 _07490_ (.A(_00554_),
    .B(_00555_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _07491_ (.A(_00557_),
    .B(_00489_),
    .Y(_00558_));
 sky130_fd_sc_hd__nor2_1 _07492_ (.A(_00552_),
    .B(_00558_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _07493_ (.A(_00685_),
    .B(_00578_),
    .Y(_00560_));
 sky130_fd_sc_hd__o21a_1 _07494_ (.A1(net23),
    .A2(_00685_),
    .B1(_00560_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _07495_ (.A0(_00567_),
    .A1(_00578_),
    .S(_00718_),
    .X(_00562_));
 sky130_fd_sc_hd__inv_2 _07496_ (.A(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__or2_1 _07497_ (.A(_00561_),
    .B(_00563_),
    .X(_00564_));
 sky130_fd_sc_hd__nor2_1 _07498_ (.A(_00237_),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__inv_2 _07499_ (.A(_00565_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand3_2 _07500_ (.A(_00531_),
    .B(_00559_),
    .C(_00566_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand3_4 _07501_ (.A(_00532_),
    .B(_00538_),
    .C(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _07502_ (.A(_00563_),
    .B(_00561_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _07503_ (.A(_00564_),
    .B(_00570_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _07504_ (.A(net90),
    .B(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__inv_2 _07505_ (.A(_00542_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _07506_ (.A(_00547_),
    .B(_00326_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _07507_ (.A(_00345_),
    .B(_00548_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _07508_ (.A(_00574_),
    .B(_00575_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _07509_ (.A(_00573_),
    .B(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand3_1 _07510_ (.A(_00357_),
    .B(_00371_),
    .C(_00373_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand3_1 _07511_ (.A(_00368_),
    .B(_00365_),
    .C(_00372_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_1 _07512_ (.A(_00579_),
    .B(_00580_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand3_1 _07513_ (.A(_00581_),
    .B(_00384_),
    .C(_00382_),
    .Y(_00582_));
 sky130_fd_sc_hd__nor2_1 _07514_ (.A(_00577_),
    .B(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand3_2 _07515_ (.A(_00480_),
    .B(_00583_),
    .C(_00566_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand3_4 _07516_ (.A(_00584_),
    .B(_00481_),
    .C(_00493_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_4 _07517_ (.A(_00585_),
    .B(_00531_),
    .Y(_00586_));
 sky130_fd_sc_hd__buf_6 _07518_ (.A(_00586_),
    .X(_00587_));
 sky130_fd_sc_hd__buf_6 _07519_ (.A(_00538_),
    .X(_00588_));
 sky130_fd_sc_hd__nand3_2 _07520_ (.A(_00587_),
    .B(_00561_),
    .C(_00588_),
    .Y(_00590_));
 sky130_fd_sc_hd__buf_12 _07521_ (.A(_00342_),
    .X(\sq.out[15] ));
 sky130_fd_sc_hd__nand3_2 _07522_ (.A(_00572_),
    .B(_00590_),
    .C(\sq.out[15] ),
    .Y(_00591_));
 sky130_fd_sc_hd__buf_12 _07523_ (.A(_00569_),
    .X(_00592_));
 sky130_fd_sc_hd__nand2_1 _07524_ (.A(_00564_),
    .B(_00237_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _07525_ (.A(_00566_),
    .B(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__clkinvlp_2 _07526_ (.A(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _07527_ (.A(_00592_),
    .B(_00595_),
    .Y(_00596_));
 sky130_fd_sc_hd__xor2_1 _07528_ (.A(_00237_),
    .B(\sq.out[15] ),
    .X(_00597_));
 sky130_fd_sc_hd__clkinvlp_2 _07529_ (.A(_00597_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand3_1 _07530_ (.A(_00587_),
    .B(_00588_),
    .C(_00598_),
    .Y(_00600_));
 sky130_fd_sc_hd__nand3_1 _07531_ (.A(_00596_),
    .B(_00600_),
    .C(_00249_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _07532_ (.A(net90),
    .B(_00594_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand3_1 _07533_ (.A(_00586_),
    .B(_00538_),
    .C(_00597_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand3_1 _07534_ (.A(_00602_),
    .B(_00603_),
    .C(_00091_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand3_1 _07535_ (.A(_00591_),
    .B(_00601_),
    .C(_00604_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_2 _07536_ (.A(_00602_),
    .B(_00603_),
    .Y(_00606_));
 sky130_fd_sc_hd__inv_2 _07537_ (.A(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _07538_ (.A(_00607_),
    .B(_00249_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _07539_ (.A(_00573_),
    .B(_00566_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _07540_ (.A(_00542_),
    .B(_00565_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _07541_ (.A(_00609_),
    .B(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__inv_2 _07542_ (.A(_00612_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _07543_ (.A(net90),
    .B(_00613_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand3_2 _07544_ (.A(_00587_),
    .B(_00588_),
    .C(_00320_),
    .Y(_00615_));
 sky130_fd_sc_hd__buf_12 _07545_ (.A(_06036_),
    .X(\sq.out[17] ));
 sky130_fd_sc_hd__nand3_2 _07546_ (.A(_00614_),
    .B(_00615_),
    .C(\sq.out[17] ),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _07547_ (.A(net120),
    .B(_00612_),
    .Y(_00617_));
 sky130_fd_sc_hd__inv_2 _07548_ (.A(_00320_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand3_1 _07549_ (.A(_00587_),
    .B(_00588_),
    .C(_00618_),
    .Y(_00619_));
 sky130_fd_sc_hd__nand3_1 _07550_ (.A(_00617_),
    .B(_00619_),
    .C(_00194_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(_00616_),
    .B(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__nor2_1 _07552_ (.A(_00608_),
    .B(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _07553_ (.A(_00622_),
    .B(_00608_),
    .Y(_00624_));
 sky130_fd_sc_hd__o21ai_2 _07554_ (.A1(_00605_),
    .A2(_00623_),
    .B1(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__inv_2 _07555_ (.A(_00385_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _07556_ (.A(_00551_),
    .B(_00566_),
    .Y(_00627_));
 sky130_fd_sc_hd__inv_2 _07557_ (.A(_00349_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _07558_ (.A(_00627_),
    .B(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__or2_1 _07559_ (.A(_00626_),
    .B(_00629_),
    .X(_00630_));
 sky130_fd_sc_hd__nand2_1 _07560_ (.A(_00629_),
    .B(_00626_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _07561_ (.A(_00630_),
    .B(_00632_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _07562_ (.A(_00592_),
    .B(_00633_),
    .Y(_00634_));
 sky130_fd_sc_hd__inv_2 _07563_ (.A(_00356_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand3_1 _07564_ (.A(_00587_),
    .B(_00588_),
    .C(_00635_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand3_1 _07565_ (.A(_00634_),
    .B(_00636_),
    .C(_06020_),
    .Y(_00637_));
 sky130_fd_sc_hd__inv_2 _07566_ (.A(_00633_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _07567_ (.A(_00569_),
    .B(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand3_2 _07568_ (.A(_00587_),
    .B(_00588_),
    .C(_00356_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand3_2 _07569_ (.A(_00639_),
    .B(_00640_),
    .C(_05119_),
    .Y(_00641_));
 sky130_fd_sc_hd__nand2_1 _07570_ (.A(_00637_),
    .B(_00641_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _07571_ (.A(_00609_),
    .B(_00324_),
    .Y(_00644_));
 sky130_fd_sc_hd__xor2_1 _07572_ (.A(_00576_),
    .B(_00644_),
    .X(_00645_));
 sky130_fd_sc_hd__nand2_1 _07573_ (.A(_00569_),
    .B(_00645_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand3_2 _07574_ (.A(_00587_),
    .B(_00588_),
    .C(_00543_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand3_1 _07575_ (.A(_00646_),
    .B(_00647_),
    .C(_06002_),
    .Y(_00648_));
 sky130_fd_sc_hd__inv_2 _07576_ (.A(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand2_1 _07577_ (.A(_00643_),
    .B(_00649_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand3_1 _07578_ (.A(_00648_),
    .B(_00637_),
    .C(_00641_),
    .Y(_00651_));
 sky130_fd_sc_hd__nand2_2 _07579_ (.A(_00650_),
    .B(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__nand2_2 _07580_ (.A(_00646_),
    .B(_00647_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _07581_ (.A(_00654_),
    .B(_06002_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand3_1 _07582_ (.A(_00646_),
    .B(_00647_),
    .C(_00214_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand2_1 _07583_ (.A(_00655_),
    .B(_00656_),
    .Y(_00657_));
 sky130_fd_sc_hd__inv_2 _07584_ (.A(_00616_),
    .Y(_00658_));
 sky130_fd_sc_hd__nand2_1 _07585_ (.A(_00657_),
    .B(_00658_),
    .Y(_00659_));
 sky130_fd_sc_hd__nand3_2 _07586_ (.A(_00655_),
    .B(_00616_),
    .C(_00656_),
    .Y(_00660_));
 sky130_fd_sc_hd__nand2_2 _07587_ (.A(_00659_),
    .B(_00660_),
    .Y(_00661_));
 sky130_fd_sc_hd__nor2_2 _07588_ (.A(_00652_),
    .B(_00661_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _07589_ (.A(_00625_),
    .B(_00662_),
    .Y(_00663_));
 sky130_fd_sc_hd__inv_2 _07590_ (.A(_00660_),
    .Y(_00665_));
 sky130_fd_sc_hd__a21boi_1 _07591_ (.A1(_00665_),
    .A2(_00650_),
    .B1_N(_00651_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _07592_ (.A(_00663_),
    .B(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _07593_ (.A(_00632_),
    .B(_00384_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand2_1 _07594_ (.A(_00668_),
    .B(_00581_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand3_1 _07595_ (.A(_00632_),
    .B(_00375_),
    .C(_00384_),
    .Y(_00670_));
 sky130_fd_sc_hd__nand2_1 _07596_ (.A(_00669_),
    .B(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__inv_2 _07597_ (.A(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(_00569_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand2_1 _07599_ (.A(_00359_),
    .B(_00364_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand3_1 _07600_ (.A(_00586_),
    .B(_00538_),
    .C(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand2_2 _07601_ (.A(_00673_),
    .B(_00675_),
    .Y(_00676_));
 sky130_fd_sc_hd__nand2_1 _07602_ (.A(_00676_),
    .B(_00460_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand3_1 _07603_ (.A(_00673_),
    .B(_00675_),
    .C(_06045_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand2_1 _07604_ (.A(_00677_),
    .B(_00678_),
    .Y(_00679_));
 sky130_fd_sc_hd__nand3_2 _07605_ (.A(_00639_),
    .B(_00640_),
    .C(_06020_),
    .Y(_00680_));
 sky130_fd_sc_hd__inv_2 _07606_ (.A(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__nand2_1 _07607_ (.A(_00679_),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__nand3_2 _07608_ (.A(_00677_),
    .B(_00680_),
    .C(_00678_),
    .Y(_00683_));
 sky130_fd_sc_hd__nand2_1 _07609_ (.A(_00682_),
    .B(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__inv_2 _07610_ (.A(_00684_),
    .Y(_00686_));
 sky130_fd_sc_hd__nor2_1 _07611_ (.A(_06045_),
    .B(_00676_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand3_1 _07612_ (.A(_00386_),
    .B(_00551_),
    .C(_00566_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand3b_1 _07613_ (.A_N(_00390_),
    .B(_00555_),
    .C(_00688_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand3_1 _07614_ (.A(_00688_),
    .B(_00389_),
    .C(_00387_),
    .Y(_00690_));
 sky130_fd_sc_hd__inv_2 _07615_ (.A(_00555_),
    .Y(_00691_));
 sky130_fd_sc_hd__nand2_1 _07616_ (.A(_00690_),
    .B(_00691_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _07617_ (.A(_00689_),
    .B(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__inv_2 _07618_ (.A(_00693_),
    .Y(_00694_));
 sky130_fd_sc_hd__nand2_1 _07619_ (.A(net90),
    .B(_00694_),
    .Y(_00695_));
 sky130_fd_sc_hd__nand2_1 _07620_ (.A(_00459_),
    .B(_00463_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand3_1 _07621_ (.A(_00586_),
    .B(_00538_),
    .C(_00697_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand3_2 _07622_ (.A(_00695_),
    .B(_00698_),
    .C(_05479_),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _07623_ (.A(_00592_),
    .B(_00693_),
    .Y(_00700_));
 sky130_fd_sc_hd__inv_2 _07624_ (.A(_00697_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand3_1 _07625_ (.A(_00587_),
    .B(_00588_),
    .C(_00701_),
    .Y(_00702_));
 sky130_fd_sc_hd__nand3_1 _07626_ (.A(_00700_),
    .B(_00702_),
    .C(_00455_),
    .Y(_00703_));
 sky130_fd_sc_hd__nand3_1 _07627_ (.A(_00687_),
    .B(_00699_),
    .C(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__nand2_1 _07628_ (.A(_00699_),
    .B(_00703_),
    .Y(_00705_));
 sky130_fd_sc_hd__inv_2 _07629_ (.A(_00676_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _07630_ (.A(_00706_),
    .B(_00460_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _07631_ (.A(_00705_),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _07632_ (.A(_00704_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__inv_2 _07633_ (.A(_00710_),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _07634_ (.A(_00686_),
    .B(_00711_),
    .Y(_00712_));
 sky130_fd_sc_hd__nand2_1 _07635_ (.A(_00692_),
    .B(_00476_),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_1 _07636_ (.A(_00713_),
    .B(_00469_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand3_1 _07637_ (.A(_00692_),
    .B(_00554_),
    .C(_00476_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand2_1 _07638_ (.A(_00714_),
    .B(_00715_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2_1 _07639_ (.A(_00716_),
    .B(_00569_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand3b_1 _07640_ (.A_N(_00454_),
    .B(_00587_),
    .C(_00588_),
    .Y(_00719_));
 sky130_fd_sc_hd__nand2_2 _07641_ (.A(_00717_),
    .B(_00719_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand2_2 _07642_ (.A(_00720_),
    .B(_00177_),
    .Y(_00721_));
 sky130_fd_sc_hd__inv_2 _07643_ (.A(_00699_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand3_1 _07644_ (.A(_00717_),
    .B(_06106_),
    .C(_00719_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand3_1 _07645_ (.A(_00721_),
    .B(_00722_),
    .C(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _07646_ (.A(_00720_),
    .B(_06106_),
    .Y(_00725_));
 sky130_fd_sc_hd__nand3_1 _07647_ (.A(_00717_),
    .B(_00177_),
    .C(_00719_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand3_1 _07648_ (.A(_00725_),
    .B(_00726_),
    .C(_00699_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand2_2 _07649_ (.A(_00724_),
    .B(_00727_),
    .Y(_00728_));
 sky130_fd_sc_hd__inv_2 _07650_ (.A(_00728_),
    .Y(_00730_));
 sky130_fd_sc_hd__nand2_1 _07651_ (.A(_00690_),
    .B(_00557_),
    .Y(_00731_));
 sky130_fd_sc_hd__inv_2 _07652_ (.A(_00485_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand2_1 _07653_ (.A(_00731_),
    .B(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand2_1 _07654_ (.A(_00733_),
    .B(_00423_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand3_1 _07655_ (.A(_00731_),
    .B(_00422_),
    .C(_00732_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(_00734_),
    .B(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand2_1 _07657_ (.A(_00736_),
    .B(_00592_),
    .Y(_00737_));
 sky130_fd_sc_hd__nand2_1 _07658_ (.A(_00407_),
    .B(_00408_),
    .Y(_00738_));
 sky130_fd_sc_hd__nand3b_1 _07659_ (.A_N(_00738_),
    .B(_00587_),
    .C(_00588_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _07660_ (.A(_00737_),
    .B(_00739_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(_00741_),
    .B(_00437_),
    .Y(_00742_));
 sky130_fd_sc_hd__clkbuf_8 _07662_ (.A(_03256_),
    .X(_00743_));
 sky130_fd_sc_hd__nand3_1 _07663_ (.A(_00737_),
    .B(_00743_),
    .C(_00739_),
    .Y(_00744_));
 sky130_fd_sc_hd__nand2_1 _07664_ (.A(_00742_),
    .B(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__inv_2 _07665_ (.A(_00721_),
    .Y(_00746_));
 sky130_fd_sc_hd__nand2_1 _07666_ (.A(_00745_),
    .B(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hd__nand3_1 _07667_ (.A(net120),
    .B(_00734_),
    .C(_00735_),
    .Y(_00748_));
 sky130_fd_sc_hd__inv_12 _07668_ (.A(net120),
    .Y(_00749_));
 sky130_fd_sc_hd__nand2_1 _07669_ (.A(_00749_),
    .B(_00738_),
    .Y(_00750_));
 sky130_fd_sc_hd__nand3_1 _07670_ (.A(_00748_),
    .B(_00750_),
    .C(_00743_),
    .Y(_00752_));
 sky130_fd_sc_hd__nand3_1 _07671_ (.A(_00737_),
    .B(_00437_),
    .C(_00739_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _07672_ (.A(_00752_),
    .B(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(_00754_),
    .B(_00721_),
    .Y(_00755_));
 sky130_fd_sc_hd__nand2_1 _07674_ (.A(_00747_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__nand2_1 _07675_ (.A(_00730_),
    .B(_00756_),
    .Y(_00757_));
 sky130_fd_sc_hd__nor2_1 _07676_ (.A(_00712_),
    .B(_00757_),
    .Y(_00758_));
 sky130_fd_sc_hd__nand2_1 _07677_ (.A(_00667_),
    .B(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__nand2_1 _07678_ (.A(_00745_),
    .B(_00721_),
    .Y(_00760_));
 sky130_fd_sc_hd__nand2_1 _07679_ (.A(_00754_),
    .B(_00746_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2_1 _07680_ (.A(_00760_),
    .B(_00761_),
    .Y(_00763_));
 sky130_fd_sc_hd__nor2_2 _07681_ (.A(_00728_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__nor2_1 _07682_ (.A(_00708_),
    .B(_00705_),
    .Y(_00765_));
 sky130_fd_sc_hd__o21ai_1 _07683_ (.A1(_00683_),
    .A2(_00765_),
    .B1(_00709_),
    .Y(_00766_));
 sky130_fd_sc_hd__nor2_1 _07684_ (.A(_00721_),
    .B(_00745_),
    .Y(_00767_));
 sky130_fd_sc_hd__o21ai_1 _07685_ (.A1(_00727_),
    .A2(_00767_),
    .B1(_00760_),
    .Y(_00768_));
 sky130_fd_sc_hd__a21oi_2 _07686_ (.A1(_00764_),
    .A2(_00766_),
    .B1(_00768_),
    .Y(_00769_));
 sky130_fd_sc_hd__nand2_1 _07687_ (.A(_00759_),
    .B(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hd__a21o_1 _07688_ (.A1(_00585_),
    .A2(_00518_),
    .B1(_00533_),
    .X(_00771_));
 sky130_fd_sc_hd__or2_1 _07689_ (.A(_00513_),
    .B(_00771_),
    .X(_00772_));
 sky130_fd_sc_hd__buf_8 _07690_ (.A(net120),
    .X(\sq.out[14] ));
 sky130_fd_sc_hd__nand2_1 _07691_ (.A(_00771_),
    .B(_00513_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand3_1 _07692_ (.A(_00772_),
    .B(\sq.out[14] ),
    .C(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__nand2_1 _07693_ (.A(_00749_),
    .B(_00509_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(_00518_),
    .B(_00519_),
    .Y(_00777_));
 sky130_fd_sc_hd__xor2_1 _07695_ (.A(_00777_),
    .B(_00585_),
    .X(_00778_));
 sky130_fd_sc_hd__inv_4 _07696_ (.A(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(_00749_),
    .B(_00500_),
    .Y(_00780_));
 sky130_fd_sc_hd__o21ai_4 _07698_ (.A1(_00749_),
    .A2(_00779_),
    .B1(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hd__a21o_1 _07699_ (.A1(_00775_),
    .A2(_00776_),
    .B1(_00781_),
    .X(_00782_));
 sky130_fd_sc_hd__nand3_2 _07700_ (.A(_00775_),
    .B(_00776_),
    .C(_00781_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_1 _07701_ (.A(_00782_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand2_1 _07702_ (.A(_00734_),
    .B(_00421_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(_00786_),
    .B(_00452_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand3_1 _07704_ (.A(_00734_),
    .B(_00488_),
    .C(_00421_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand3_4 _07705_ (.A(_00787_),
    .B(_00788_),
    .C(net120),
    .Y(_00789_));
 sky130_fd_sc_hd__a21o_1 _07706_ (.A1(_00427_),
    .A2(_00436_),
    .B1(_00592_),
    .X(_00790_));
 sky130_fd_sc_hd__nand3_4 _07707_ (.A(_00789_),
    .B(_00283_),
    .C(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__inv_2 _07708_ (.A(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__nand2_1 _07709_ (.A(_00792_),
    .B(_00781_),
    .Y(_00793_));
 sky130_fd_sc_hd__inv_2 _07710_ (.A(_00781_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand2_1 _07711_ (.A(_00794_),
    .B(_00791_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand2_1 _07712_ (.A(_00793_),
    .B(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand2_2 _07713_ (.A(_00789_),
    .B(_00790_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _07714_ (.A(_00797_),
    .B(_03650_),
    .Y(_00798_));
 sky130_fd_sc_hd__nand2_1 _07715_ (.A(_00798_),
    .B(_00791_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_1 _07716_ (.A(_00799_),
    .B(_00742_),
    .Y(_00800_));
 sky130_fd_sc_hd__nand3b_1 _07717_ (.A_N(_00742_),
    .B(_00798_),
    .C(_00791_),
    .Y(_00801_));
 sky130_fd_sc_hd__nand3_1 _07718_ (.A(_00796_),
    .B(_00800_),
    .C(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__nor2_2 _07719_ (.A(_00785_),
    .B(_00802_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand2_1 _07720_ (.A(_00770_),
    .B(_00803_),
    .Y(_00805_));
 sky130_fd_sc_hd__nor2_1 _07721_ (.A(_00781_),
    .B(_00791_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand2_1 _07722_ (.A(_00791_),
    .B(_00781_),
    .Y(_00807_));
 sky130_fd_sc_hd__o21ai_1 _07723_ (.A1(_00806_),
    .A2(_00800_),
    .B1(_00807_),
    .Y(_00808_));
 sky130_fd_sc_hd__a21boi_4 _07724_ (.A1(_00808_),
    .A2(_00784_),
    .B1_N(_00782_),
    .Y(_00809_));
 sky130_fd_sc_hd__nand2_1 _07725_ (.A(_00601_),
    .B(_00604_),
    .Y(_00810_));
 sky130_fd_sc_hd__inv_2 _07726_ (.A(_00591_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(_00810_),
    .B(_00811_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _07728_ (.A(_00812_),
    .B(_00605_),
    .Y(_00813_));
 sky130_fd_sc_hd__inv_2 _07729_ (.A(_00608_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _07730_ (.A(_00614_),
    .B(_00615_),
    .Y(_00816_));
 sky130_fd_sc_hd__nand2_1 _07731_ (.A(_00816_),
    .B(\sq.out[17] ),
    .Y(_00817_));
 sky130_fd_sc_hd__nand3_1 _07732_ (.A(_00614_),
    .B(_00615_),
    .C(_00194_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_00817_),
    .B(_00818_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _07734_ (.A(_00814_),
    .B(_00819_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand2_2 _07735_ (.A(_00820_),
    .B(_00624_),
    .Y(_00821_));
 sky130_fd_sc_hd__nor2_2 _07736_ (.A(_00813_),
    .B(_00821_),
    .Y(_00822_));
 sky130_fd_sc_hd__nand2_2 _07737_ (.A(_00822_),
    .B(_00662_),
    .Y(_00823_));
 sky130_fd_sc_hd__nor2_1 _07738_ (.A(_00710_),
    .B(_00684_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_1 _07739_ (.A(_00764_),
    .B(_00824_),
    .Y(_00825_));
 sky130_fd_sc_hd__nor2_1 _07740_ (.A(_00823_),
    .B(_00825_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_4 _07741_ (.A(_00718_),
    .B(net1),
    .Y(_00828_));
 sky130_fd_sc_hd__inv_2 _07742_ (.A(_00828_),
    .Y(_00829_));
 sky130_fd_sc_hd__nor2_1 _07743_ (.A(_00829_),
    .B(_00563_),
    .Y(_00830_));
 sky130_fd_sc_hd__a21o_1 _07744_ (.A1(net90),
    .A2(_00563_),
    .B1(_00830_),
    .X(_00831_));
 sky130_fd_sc_hd__inv_2 _07745_ (.A(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand2_2 _07746_ (.A(_00572_),
    .B(_00590_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_00833_),
    .B(_00425_),
    .Y(_00834_));
 sky130_fd_sc_hd__nand2_1 _07748_ (.A(_00834_),
    .B(_00591_),
    .Y(_00835_));
 sky130_fd_sc_hd__or2_1 _07749_ (.A(_00832_),
    .B(_00835_),
    .X(_00836_));
 sky130_fd_sc_hd__buf_6 _07750_ (.A(_00836_),
    .X(_00838_));
 sky130_fd_sc_hd__nand3_2 _07751_ (.A(_00803_),
    .B(_00827_),
    .C(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__nand3_4 _07752_ (.A(_00805_),
    .B(_00809_),
    .C(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__buf_6 _07753_ (.A(_00840_),
    .X(_00841_));
 sky130_fd_sc_hd__inv_6 _07754_ (.A(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__buf_6 _07755_ (.A(_00842_),
    .X(_00843_));
 sky130_fd_sc_hd__buf_4 _07756_ (.A(_00843_),
    .X(_00844_));
 sky130_fd_sc_hd__buf_12 _07757_ (.A(_00841_),
    .X(_00845_));
 sky130_fd_sc_hd__buf_8 _07758_ (.A(_00845_),
    .X(\sq.out[13] ));
 sky130_fd_sc_hd__inv_2 _07759_ (.A(_00823_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand3_1 _07760_ (.A(_00758_),
    .B(_00846_),
    .C(_00838_),
    .Y(_00848_));
 sky130_fd_sc_hd__nand3_2 _07761_ (.A(_00848_),
    .B(_00769_),
    .C(_00759_),
    .Y(_00849_));
 sky130_fd_sc_hd__nand2_2 _07762_ (.A(_00849_),
    .B(_00803_),
    .Y(_00850_));
 sky130_fd_sc_hd__buf_6 _07763_ (.A(_00850_),
    .X(_00851_));
 sky130_fd_sc_hd__buf_6 _07764_ (.A(_00809_),
    .X(_00852_));
 sky130_fd_sc_hd__nand2_1 _07765_ (.A(_00639_),
    .B(_00640_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand3_1 _07766_ (.A(_00851_),
    .B(_00852_),
    .C(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__nand2_1 _07767_ (.A(_00822_),
    .B(_00838_),
    .Y(_00855_));
 sky130_fd_sc_hd__inv_2 _07768_ (.A(_00625_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(_00855_),
    .B(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _07770_ (.A(_00661_),
    .Y(_00859_));
 sky130_fd_sc_hd__nand2_1 _07771_ (.A(_00857_),
    .B(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__nand2_1 _07772_ (.A(_00860_),
    .B(_00660_),
    .Y(_00861_));
 sky130_fd_sc_hd__inv_2 _07773_ (.A(_00652_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _07774_ (.A(_00861_),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__nand3_1 _07775_ (.A(_00860_),
    .B(_00652_),
    .C(_00660_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2_1 _07776_ (.A(_00863_),
    .B(_00864_),
    .Y(_00865_));
 sky130_fd_sc_hd__inv_2 _07777_ (.A(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__nand2_1 _07778_ (.A(_00866_),
    .B(_00841_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2_1 _07779_ (.A(_00854_),
    .B(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _07780_ (.A(_00868_),
    .B(_00460_),
    .Y(_00870_));
 sky130_fd_sc_hd__nand3_1 _07781_ (.A(_00854_),
    .B(_00867_),
    .C(_06045_),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_1 _07782_ (.A(_00870_),
    .B(_00871_),
    .Y(_00872_));
 sky130_fd_sc_hd__nand3_1 _07783_ (.A(_00851_),
    .B(_00852_),
    .C(_00654_),
    .Y(_00873_));
 sky130_fd_sc_hd__or2_1 _07784_ (.A(_00859_),
    .B(_00857_),
    .X(_00874_));
 sky130_fd_sc_hd__nand2_1 _07785_ (.A(_00874_),
    .B(_00860_),
    .Y(_00875_));
 sky130_fd_sc_hd__inv_2 _07786_ (.A(_00875_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand2_1 _07787_ (.A(_00841_),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand3_1 _07788_ (.A(_00873_),
    .B(_00877_),
    .C(_06020_),
    .Y(_00878_));
 sky130_fd_sc_hd__inv_2 _07789_ (.A(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _07790_ (.A(_00872_),
    .B(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand3_2 _07791_ (.A(_00870_),
    .B(_00871_),
    .C(_00878_),
    .Y(_00881_));
 sky130_fd_sc_hd__nand2_1 _07792_ (.A(_00880_),
    .B(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__inv_2 _07793_ (.A(_00882_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand3_1 _07794_ (.A(_00851_),
    .B(_00852_),
    .C(_00676_),
    .Y(_00884_));
 sky130_fd_sc_hd__nand3_1 _07795_ (.A(_00822_),
    .B(_00662_),
    .C(_00838_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand3b_1 _07796_ (.A_N(_00667_),
    .B(_00684_),
    .C(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand3_1 _07797_ (.A(_00885_),
    .B(_00666_),
    .C(_00663_),
    .Y(_00887_));
 sky130_fd_sc_hd__nand2_1 _07798_ (.A(_00887_),
    .B(_00686_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(_00886_),
    .B(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__inv_2 _07800_ (.A(_00889_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_1 _07801_ (.A(net104),
    .B(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__buf_12 _07802_ (.A(_05479_),
    .X(\sq.out[21] ));
 sky130_fd_sc_hd__nand3_2 _07803_ (.A(_00884_),
    .B(_00892_),
    .C(\sq.out[21] ),
    .Y(_00893_));
 sky130_fd_sc_hd__nand3_1 _07804_ (.A(_00851_),
    .B(_00852_),
    .C(_00706_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(net104),
    .B(_00889_),
    .Y(_00895_));
 sky130_fd_sc_hd__nand3_1 _07806_ (.A(_00894_),
    .B(_00895_),
    .C(_00455_),
    .Y(_00896_));
 sky130_fd_sc_hd__nand2_2 _07807_ (.A(_00893_),
    .B(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__inv_2 _07808_ (.A(_00897_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand3_2 _07809_ (.A(_00854_),
    .B(_00867_),
    .C(_00460_),
    .Y(_00899_));
 sky130_fd_sc_hd__nand2_1 _07810_ (.A(_00898_),
    .B(_00899_),
    .Y(_00901_));
 sky130_fd_sc_hd__inv_2 _07811_ (.A(_00899_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(_00897_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand2_1 _07813_ (.A(_00901_),
    .B(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_1 _07814_ (.A(_00883_),
    .B(_00904_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(_00888_),
    .B(_00683_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand2_1 _07816_ (.A(_00906_),
    .B(_00711_),
    .Y(_00907_));
 sky130_fd_sc_hd__nand3_1 _07817_ (.A(_00888_),
    .B(_00710_),
    .C(_00683_),
    .Y(_00908_));
 sky130_fd_sc_hd__nand3_1 _07818_ (.A(_00845_),
    .B(_00907_),
    .C(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand2_1 _07819_ (.A(_00695_),
    .B(_00698_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand2_1 _07820_ (.A(_00842_),
    .B(_00910_),
    .Y(_00912_));
 sky130_fd_sc_hd__nand3_1 _07821_ (.A(_00909_),
    .B(_00912_),
    .C(_06106_),
    .Y(_00913_));
 sky130_fd_sc_hd__nand2_1 _07822_ (.A(_00907_),
    .B(_00908_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _07823_ (.A(_00914_),
    .B(net104),
    .Y(_00915_));
 sky130_fd_sc_hd__nand3b_1 _07824_ (.A_N(_00910_),
    .B(_00851_),
    .C(_00852_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand3_1 _07825_ (.A(_00915_),
    .B(_00916_),
    .C(_00177_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_1 _07826_ (.A(_00913_),
    .B(_00917_),
    .Y(_00918_));
 sky130_fd_sc_hd__clkinvlp_2 _07827_ (.A(_00893_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand2_1 _07828_ (.A(_00918_),
    .B(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__nand3_2 _07829_ (.A(_00913_),
    .B(_00917_),
    .C(_00893_),
    .Y(_00921_));
 sky130_fd_sc_hd__nand2_2 _07830_ (.A(_00920_),
    .B(_00921_),
    .Y(_00923_));
 sky130_fd_sc_hd__inv_2 _07831_ (.A(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand2_1 _07832_ (.A(_00887_),
    .B(_00824_),
    .Y(_00925_));
 sky130_fd_sc_hd__inv_2 _07833_ (.A(_00766_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_1 _07834_ (.A(_00925_),
    .B(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand2_1 _07835_ (.A(_00927_),
    .B(_00730_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand3_1 _07836_ (.A(_00925_),
    .B(_00728_),
    .C(_00926_),
    .Y(_00929_));
 sky130_fd_sc_hd__nand2_1 _07837_ (.A(_00928_),
    .B(_00929_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _07838_ (.A(_00930_),
    .B(_00845_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _07839_ (.A(_00842_),
    .B(_00720_),
    .Y(_00932_));
 sky130_fd_sc_hd__nand2_2 _07840_ (.A(_00931_),
    .B(_00932_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand2_2 _07841_ (.A(_00934_),
    .B(_00437_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand3_1 _07842_ (.A(_00931_),
    .B(_00932_),
    .C(_00743_),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(_00935_),
    .B(_00936_),
    .Y(_00937_));
 sky130_fd_sc_hd__nand2_1 _07844_ (.A(_00915_),
    .B(_00916_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_2 _07845_ (.A(_00938_),
    .B(_00177_),
    .Y(_00939_));
 sky130_fd_sc_hd__inv_2 _07846_ (.A(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _07847_ (.A(_00937_),
    .B(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand3_1 _07848_ (.A(_00931_),
    .B(_00932_),
    .C(_00437_),
    .Y(_00942_));
 sky130_fd_sc_hd__nand3_1 _07849_ (.A(_00845_),
    .B(_00928_),
    .C(_00929_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand3b_1 _07850_ (.A_N(_00720_),
    .B(_00851_),
    .C(_00852_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand3_1 _07851_ (.A(_00943_),
    .B(_00945_),
    .C(_00743_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _07852_ (.A(_00942_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _07853_ (.A(_00947_),
    .B(_00939_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _07854_ (.A(_00941_),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_1 _07855_ (.A(_00924_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__nor2_1 _07856_ (.A(_00905_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__inv_2 _07857_ (.A(_00654_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand3_1 _07858_ (.A(_00851_),
    .B(_00852_),
    .C(_00952_),
    .Y(_00953_));
 sky130_fd_sc_hd__nand2_1 _07859_ (.A(_00845_),
    .B(_00875_),
    .Y(_00954_));
 sky130_fd_sc_hd__buf_12 _07860_ (.A(_06020_),
    .X(\sq.out[19] ));
 sky130_fd_sc_hd__nand3_1 _07861_ (.A(_00953_),
    .B(_00954_),
    .C(\sq.out[19] ),
    .Y(_00956_));
 sky130_fd_sc_hd__nand3_1 _07862_ (.A(_00873_),
    .B(_00877_),
    .C(_05119_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_1 _07863_ (.A(_00956_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__nand3_1 _07864_ (.A(_00850_),
    .B(_00809_),
    .C(_00816_),
    .Y(_00959_));
 sky130_fd_sc_hd__a21boi_1 _07865_ (.A1(_00838_),
    .A2(_00812_),
    .B1_N(_00605_),
    .Y(_00960_));
 sky130_fd_sc_hd__xor2_1 _07866_ (.A(_00821_),
    .B(_00960_),
    .X(_00961_));
 sky130_fd_sc_hd__nand2_1 _07867_ (.A(_00840_),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__nand3_2 _07868_ (.A(_00959_),
    .B(_00962_),
    .C(_06002_),
    .Y(_00963_));
 sky130_fd_sc_hd__inv_2 _07869_ (.A(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__nand2_1 _07870_ (.A(_00958_),
    .B(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand3_1 _07871_ (.A(_00963_),
    .B(_00956_),
    .C(_00957_),
    .Y(_00966_));
 sky130_fd_sc_hd__nand2_1 _07872_ (.A(_00965_),
    .B(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand2_1 _07873_ (.A(_00959_),
    .B(_00962_),
    .Y(_00968_));
 sky130_fd_sc_hd__nand2_1 _07874_ (.A(_00968_),
    .B(_00214_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_1 _07875_ (.A(_00969_),
    .B(_00963_),
    .Y(_00970_));
 sky130_fd_sc_hd__nand3_2 _07876_ (.A(_00851_),
    .B(_00852_),
    .C(_00606_),
    .Y(_00971_));
 sky130_fd_sc_hd__xor2_2 _07877_ (.A(_00813_),
    .B(_00838_),
    .X(_00972_));
 sky130_fd_sc_hd__inv_2 _07878_ (.A(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__nand2_1 _07879_ (.A(_00841_),
    .B(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand3_1 _07880_ (.A(_00971_),
    .B(_00974_),
    .C(\sq.out[17] ),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_1 _07881_ (.A(_00970_),
    .B(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_2 _07882_ (.A(_00971_),
    .B(_00974_),
    .Y(_00978_));
 sky130_fd_sc_hd__nor2_1 _07883_ (.A(_00194_),
    .B(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__nand3_1 _07884_ (.A(_00979_),
    .B(_00969_),
    .C(_00963_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _07885_ (.A(_00977_),
    .B(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__nor2_2 _07886_ (.A(_00981_),
    .B(_00967_),
    .Y(_00982_));
 sky130_fd_sc_hd__inv_2 _07887_ (.A(_00833_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand3_1 _07888_ (.A(_00851_),
    .B(_00852_),
    .C(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _07889_ (.A(_00835_),
    .B(_00832_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _07890_ (.A(_00838_),
    .B(_00985_),
    .Y(_00987_));
 sky130_fd_sc_hd__inv_2 _07891_ (.A(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _07892_ (.A(net104),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__nand3_1 _07893_ (.A(_00984_),
    .B(_00989_),
    .C(_00249_),
    .Y(_00990_));
 sky130_fd_sc_hd__nand3_2 _07894_ (.A(_00850_),
    .B(_00809_),
    .C(_00833_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand2_2 _07895_ (.A(_00840_),
    .B(_00987_),
    .Y(_00992_));
 sky130_fd_sc_hd__nand3_1 _07896_ (.A(_00991_),
    .B(_00992_),
    .C(_00091_),
    .Y(_00993_));
 sky130_fd_sc_hd__nand2_1 _07897_ (.A(_00990_),
    .B(_00993_),
    .Y(_00994_));
 sky130_fd_sc_hd__xor2_1 _07898_ (.A(_00563_),
    .B(\sq.out[14] ),
    .X(_00995_));
 sky130_fd_sc_hd__inv_2 _07899_ (.A(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hd__nand3_1 _07900_ (.A(_00850_),
    .B(_00809_),
    .C(_00996_),
    .Y(_00998_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(_00563_),
    .B(_00829_),
    .Y(_00999_));
 sky130_fd_sc_hd__and2b_1 _07902_ (.A_N(_00830_),
    .B(_00999_),
    .X(_01000_));
 sky130_fd_sc_hd__nand2_1 _07903_ (.A(_00840_),
    .B(_01000_),
    .Y(_01001_));
 sky130_fd_sc_hd__nand2_2 _07904_ (.A(_00998_),
    .B(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__nand2_1 _07905_ (.A(_01002_),
    .B(\sq.out[15] ),
    .Y(_01003_));
 sky130_fd_sc_hd__inv_2 _07906_ (.A(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__nand2_1 _07907_ (.A(_00994_),
    .B(_01004_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand3_1 _07908_ (.A(_01003_),
    .B(_00990_),
    .C(_00993_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand2_1 _07909_ (.A(_01005_),
    .B(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_1 _07910_ (.A(_00978_),
    .B(\sq.out[17] ),
    .Y(_01009_));
 sky130_fd_sc_hd__nand3_1 _07911_ (.A(_00971_),
    .B(_00974_),
    .C(_00194_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_1 _07912_ (.A(_01009_),
    .B(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand3_2 _07913_ (.A(_00991_),
    .B(_00992_),
    .C(_00249_),
    .Y(_01012_));
 sky130_fd_sc_hd__inv_2 _07914_ (.A(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _07915_ (.A(_01011_),
    .B(_01013_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand3_1 _07916_ (.A(_00851_),
    .B(_00852_),
    .C(_00607_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _07917_ (.A(net104),
    .B(_00972_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand3_1 _07918_ (.A(_01015_),
    .B(_01016_),
    .C(_00194_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _07919_ (.A(_00976_),
    .B(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _07920_ (.A(_01018_),
    .B(_01012_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_1 _07921_ (.A(_01014_),
    .B(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hd__nor2_2 _07922_ (.A(_01021_),
    .B(_01007_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand2_1 _07923_ (.A(_00982_),
    .B(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__inv_2 _07924_ (.A(_01023_),
    .Y(_01024_));
 sky130_fd_sc_hd__xor2_4 _07925_ (.A(_00828_),
    .B(_00845_),
    .X(_01025_));
 sky130_fd_sc_hd__nor2_1 _07926_ (.A(\sq.out[15] ),
    .B(_01002_),
    .Y(_01026_));
 sky130_fd_sc_hd__nor2_1 _07927_ (.A(_01026_),
    .B(_01004_),
    .Y(_01027_));
 sky130_fd_sc_hd__o21ai_4 _07928_ (.A1(\sq.out[14] ),
    .A2(_01025_),
    .B1(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand3_1 _07929_ (.A(_00951_),
    .B(_01024_),
    .C(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _07930_ (.A(_00937_),
    .B(_00939_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _07931_ (.A(_00947_),
    .B(_00940_),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_1 _07932_ (.A(_01031_),
    .B(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hd__nor2_1 _07933_ (.A(_00923_),
    .B(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__nor2_1 _07934_ (.A(_00899_),
    .B(_00897_),
    .Y(_01035_));
 sky130_fd_sc_hd__nand2_1 _07935_ (.A(_00897_),
    .B(_00899_),
    .Y(_01036_));
 sky130_fd_sc_hd__o21ai_1 _07936_ (.A1(_00881_),
    .A2(_01035_),
    .B1(_01036_),
    .Y(_01037_));
 sky130_fd_sc_hd__nor2_1 _07937_ (.A(_00939_),
    .B(_00937_),
    .Y(_01038_));
 sky130_fd_sc_hd__o21ai_1 _07938_ (.A1(_00921_),
    .A2(_01038_),
    .B1(_01031_),
    .Y(_01039_));
 sky130_fd_sc_hd__a21oi_2 _07939_ (.A1(_01034_),
    .A2(_01037_),
    .B1(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__nor2_1 _07940_ (.A(_01012_),
    .B(_01018_),
    .Y(_01042_));
 sky130_fd_sc_hd__o21ai_1 _07941_ (.A1(_01006_),
    .A2(_01042_),
    .B1(_01020_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand2_1 _07942_ (.A(_01043_),
    .B(_00982_),
    .Y(_01044_));
 sky130_fd_sc_hd__clkinvlp_2 _07943_ (.A(_00977_),
    .Y(_01045_));
 sky130_fd_sc_hd__a21boi_1 _07944_ (.A1(_01045_),
    .A2(_00965_),
    .B1_N(_00966_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2_1 _07945_ (.A(_01044_),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__nand2_1 _07946_ (.A(_00951_),
    .B(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__nand3_2 _07947_ (.A(_01029_),
    .B(_01040_),
    .C(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand2_1 _07948_ (.A(_00800_),
    .B(_00801_),
    .Y(_01050_));
 sky130_fd_sc_hd__inv_2 _07949_ (.A(_01050_),
    .Y(_01051_));
 sky130_fd_sc_hd__or2_1 _07950_ (.A(_01051_),
    .B(_00849_),
    .X(_01053_));
 sky130_fd_sc_hd__nand2_1 _07951_ (.A(_00849_),
    .B(_01051_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _07952_ (.A(_01053_),
    .B(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__nand2_1 _07953_ (.A(_01055_),
    .B(_00845_),
    .Y(_01056_));
 sky130_fd_sc_hd__o21ai_4 _07954_ (.A1(_00797_),
    .A2(_00845_),
    .B1(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__inv_2 _07955_ (.A(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__nand2_1 _07956_ (.A(_01054_),
    .B(_00800_),
    .Y(_01059_));
 sky130_fd_sc_hd__or2_1 _07957_ (.A(_00796_),
    .B(_01059_),
    .X(_01060_));
 sky130_fd_sc_hd__nand2_1 _07958_ (.A(_01059_),
    .B(_00796_),
    .Y(_01061_));
 sky130_fd_sc_hd__nand3_1 _07959_ (.A(_01060_),
    .B(\sq.out[13] ),
    .C(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__nand2_1 _07960_ (.A(_00842_),
    .B(_00794_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand2_1 _07961_ (.A(_01062_),
    .B(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__or2_4 _07962_ (.A(_01058_),
    .B(_01064_),
    .X(_01065_));
 sky130_fd_sc_hd__nand2_1 _07963_ (.A(_01064_),
    .B(_01058_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_01065_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _07965_ (.A(_00928_),
    .B(_00727_),
    .Y(_01068_));
 sky130_fd_sc_hd__nand2_1 _07966_ (.A(_01068_),
    .B(_00756_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand3_1 _07967_ (.A(_00928_),
    .B(_00763_),
    .C(_00727_),
    .Y(_01070_));
 sky130_fd_sc_hd__nand3_2 _07968_ (.A(_01069_),
    .B(_01070_),
    .C(_00845_),
    .Y(_01071_));
 sky130_fd_sc_hd__or2_1 _07969_ (.A(_00741_),
    .B(_00845_),
    .X(_01072_));
 sky130_fd_sc_hd__nand2_1 _07970_ (.A(_01071_),
    .B(_01072_),
    .Y(_01074_));
 sky130_fd_sc_hd__inv_2 _07971_ (.A(_01074_),
    .Y(_01075_));
 sky130_fd_sc_hd__nand3_1 _07972_ (.A(_01075_),
    .B(_00283_),
    .C(_01057_),
    .Y(_01076_));
 sky130_fd_sc_hd__nand3_1 _07973_ (.A(_01071_),
    .B(_00283_),
    .C(_01072_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand2_1 _07974_ (.A(_01077_),
    .B(_01058_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand2_1 _07975_ (.A(_01076_),
    .B(_01078_),
    .Y(_01079_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(_01074_),
    .B(_00283_),
    .Y(_01080_));
 sky130_fd_sc_hd__clkbuf_8 _07977_ (.A(_03650_),
    .X(_01081_));
 sky130_fd_sc_hd__nand3_1 _07978_ (.A(_01071_),
    .B(_01081_),
    .C(_01072_),
    .Y(_01082_));
 sky130_fd_sc_hd__nand2_1 _07979_ (.A(_01080_),
    .B(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__inv_2 _07980_ (.A(_00935_),
    .Y(_01085_));
 sky130_fd_sc_hd__nand2_1 _07981_ (.A(_01083_),
    .B(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__nand3_2 _07982_ (.A(_01080_),
    .B(_00935_),
    .C(_01082_),
    .Y(_01087_));
 sky130_fd_sc_hd__nand3_1 _07983_ (.A(_01079_),
    .B(_01086_),
    .C(_01087_),
    .Y(_01088_));
 sky130_fd_sc_hd__nor2_2 _07984_ (.A(_01088_),
    .B(_01067_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_2 _07985_ (.A(_01049_),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__buf_4 _07986_ (.A(_01090_),
    .X(_01091_));
 sky130_fd_sc_hd__nor2_1 _07987_ (.A(_01057_),
    .B(_01077_),
    .Y(_01092_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(_01077_),
    .B(_01057_),
    .Y(_01093_));
 sky130_fd_sc_hd__o21ai_2 _07989_ (.A1(_01092_),
    .A2(_01087_),
    .B1(_01093_),
    .Y(_01094_));
 sky130_fd_sc_hd__a21boi_4 _07990_ (.A1(_01094_),
    .A2(_01065_),
    .B1_N(_01066_),
    .Y(_01096_));
 sky130_fd_sc_hd__buf_6 _07991_ (.A(_01096_),
    .X(_01097_));
 sky130_fd_sc_hd__nand2_1 _07992_ (.A(_00873_),
    .B(_00877_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand3_1 _07993_ (.A(_01091_),
    .B(_01097_),
    .C(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__nand2_1 _07994_ (.A(_01048_),
    .B(_01040_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_1 _07995_ (.A(_01100_),
    .B(_01089_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2_1 _07996_ (.A(_00898_),
    .B(_00902_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand2_1 _07997_ (.A(_01102_),
    .B(_01036_),
    .Y(_01103_));
 sky130_fd_sc_hd__nor2_1 _07998_ (.A(_00882_),
    .B(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _07999_ (.A(_01034_),
    .B(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__nor2_1 _08000_ (.A(_01023_),
    .B(_01105_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand3_2 _08001_ (.A(_01089_),
    .B(_01107_),
    .C(_01028_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand3_4 _08002_ (.A(_01101_),
    .B(_01096_),
    .C(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__buf_8 _08003_ (.A(_01109_),
    .X(_01110_));
 sky130_fd_sc_hd__nand2_1 _08004_ (.A(_01022_),
    .B(_01028_),
    .Y(_01111_));
 sky130_fd_sc_hd__inv_2 _08005_ (.A(_01043_),
    .Y(_01112_));
 sky130_fd_sc_hd__nand2_1 _08006_ (.A(_01111_),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__inv_2 _08007_ (.A(_00981_),
    .Y(_01114_));
 sky130_fd_sc_hd__nand2_1 _08008_ (.A(_01113_),
    .B(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _08009_ (.A(_01115_),
    .B(_00977_),
    .Y(_01116_));
 sky130_fd_sc_hd__inv_2 _08010_ (.A(_00967_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand2_1 _08011_ (.A(_01116_),
    .B(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand3_1 _08012_ (.A(_01115_),
    .B(_00967_),
    .C(_00977_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _08013_ (.A(_01119_),
    .B(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__inv_2 _08014_ (.A(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand2_2 _08015_ (.A(_01110_),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__nand2_1 _08016_ (.A(_01099_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _08017_ (.A(_01124_),
    .B(_00460_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand3_1 _08018_ (.A(_01099_),
    .B(_01123_),
    .C(_06045_),
    .Y(_01126_));
 sky130_fd_sc_hd__nand2_1 _08019_ (.A(_01125_),
    .B(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand3_2 _08020_ (.A(_01090_),
    .B(_01096_),
    .C(_00968_),
    .Y(_01129_));
 sky130_fd_sc_hd__or2_1 _08021_ (.A(_01114_),
    .B(_01113_),
    .X(_01130_));
 sky130_fd_sc_hd__nand2_1 _08022_ (.A(_01130_),
    .B(_01115_),
    .Y(_01131_));
 sky130_fd_sc_hd__inv_2 _08023_ (.A(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__nand2_1 _08024_ (.A(_01109_),
    .B(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand3_2 _08025_ (.A(_01129_),
    .B(_01133_),
    .C(\sq.out[19] ),
    .Y(_01134_));
 sky130_fd_sc_hd__inv_2 _08026_ (.A(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_1 _08027_ (.A(_01127_),
    .B(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand3_2 _08028_ (.A(_01125_),
    .B(_01126_),
    .C(_01134_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand2_1 _08029_ (.A(_01136_),
    .B(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__inv_2 _08030_ (.A(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand3_1 _08031_ (.A(_01090_),
    .B(_01096_),
    .C(_00868_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand3_1 _08032_ (.A(_00982_),
    .B(_01022_),
    .C(_01028_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand3b_1 _08033_ (.A_N(_01047_),
    .B(_00882_),
    .C(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand3_1 _08034_ (.A(_01141_),
    .B(_01046_),
    .C(_01044_),
    .Y(_01143_));
 sky130_fd_sc_hd__nand2_1 _08035_ (.A(_01143_),
    .B(_00883_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand2_1 _08036_ (.A(_01142_),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__inv_2 _08037_ (.A(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__nand2_1 _08038_ (.A(_01109_),
    .B(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hd__nand2_1 _08039_ (.A(_01140_),
    .B(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__nand2_1 _08040_ (.A(_01148_),
    .B(_00455_),
    .Y(_01150_));
 sky130_fd_sc_hd__nand3_2 _08041_ (.A(_01140_),
    .B(_01147_),
    .C(\sq.out[21] ),
    .Y(_01151_));
 sky130_fd_sc_hd__nand2_1 _08042_ (.A(_01150_),
    .B(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand3_2 _08043_ (.A(_01099_),
    .B(_01123_),
    .C(_00460_),
    .Y(_01153_));
 sky130_fd_sc_hd__inv_2 _08044_ (.A(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand2_1 _08045_ (.A(_01152_),
    .B(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__nand3_1 _08046_ (.A(_01150_),
    .B(_01153_),
    .C(_01151_),
    .Y(_01156_));
 sky130_fd_sc_hd__nand2_1 _08047_ (.A(_01155_),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand2_1 _08048_ (.A(_01139_),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(_01144_),
    .B(_00881_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_01159_),
    .B(_00904_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand3_1 _08051_ (.A(_01144_),
    .B(_01103_),
    .C(_00881_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2_1 _08052_ (.A(_01161_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _08053_ (.A(_01163_),
    .B(net118),
    .Y(_01164_));
 sky130_fd_sc_hd__nand2_1 _08054_ (.A(_00884_),
    .B(_00892_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand3b_1 _08055_ (.A_N(_01165_),
    .B(_01091_),
    .C(_01097_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand3_1 _08056_ (.A(_01164_),
    .B(_01166_),
    .C(_06106_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand3_2 _08057_ (.A(_01110_),
    .B(_01161_),
    .C(_01162_),
    .Y(_01168_));
 sky130_fd_sc_hd__nand3_1 _08058_ (.A(_01091_),
    .B(_01097_),
    .C(_01165_),
    .Y(_01169_));
 sky130_fd_sc_hd__nand3_2 _08059_ (.A(_01168_),
    .B(_00177_),
    .C(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__nand2_1 _08060_ (.A(_01167_),
    .B(_01170_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand2_1 _08061_ (.A(_01172_),
    .B(_01151_),
    .Y(_01173_));
 sky130_fd_sc_hd__inv_2 _08062_ (.A(_01151_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand3_1 _08063_ (.A(_01174_),
    .B(_01167_),
    .C(_01170_),
    .Y(_01175_));
 sky130_fd_sc_hd__nand2_1 _08064_ (.A(_01173_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__inv_2 _08065_ (.A(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2_1 _08066_ (.A(_01143_),
    .B(_01104_),
    .Y(_01178_));
 sky130_fd_sc_hd__inv_2 _08067_ (.A(_01037_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand2_1 _08068_ (.A(_01178_),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _08069_ (.A(_01180_),
    .B(_00924_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand3_1 _08070_ (.A(_01178_),
    .B(_00923_),
    .C(_01179_),
    .Y(_01183_));
 sky130_fd_sc_hd__nand2_1 _08071_ (.A(_01181_),
    .B(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _08072_ (.A(_01184_),
    .B(_01110_),
    .Y(_01185_));
 sky130_fd_sc_hd__inv_4 _08073_ (.A(_01109_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _08074_ (.A(_01186_),
    .B(_00938_),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _08075_ (.A(_01185_),
    .B(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__nand2_1 _08076_ (.A(_01188_),
    .B(_00437_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand3_1 _08077_ (.A(_01185_),
    .B(_01187_),
    .C(_00743_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(_01189_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__inv_2 _08079_ (.A(_01170_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _08080_ (.A(_01191_),
    .B(_01192_),
    .Y(_01194_));
 sky130_fd_sc_hd__nand3_1 _08081_ (.A(_01185_),
    .B(_01187_),
    .C(_00437_),
    .Y(_01195_));
 sky130_fd_sc_hd__buf_12 _08082_ (.A(_01110_),
    .X(\sq.out[12] ));
 sky130_fd_sc_hd__nand3_1 _08083_ (.A(\sq.out[12] ),
    .B(_01181_),
    .C(_01183_),
    .Y(_01196_));
 sky130_fd_sc_hd__nand3b_1 _08084_ (.A_N(_00938_),
    .B(_01091_),
    .C(_01097_),
    .Y(_01197_));
 sky130_fd_sc_hd__nand3_1 _08085_ (.A(_01196_),
    .B(_01197_),
    .C(_00743_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_1 _08086_ (.A(_01195_),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(_01199_),
    .B(_01170_),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _08088_ (.A(_01194_),
    .B(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__nand2_1 _08089_ (.A(_01177_),
    .B(_01201_),
    .Y(_01202_));
 sky130_fd_sc_hd__nor2_2 _08090_ (.A(_01158_),
    .B(_01202_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand3_1 _08091_ (.A(_01091_),
    .B(_01097_),
    .C(_01002_),
    .Y(_01205_));
 sky130_fd_sc_hd__inv_2 _08092_ (.A(_01025_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_1 _08093_ (.A(_01206_),
    .B(_00749_),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _08094_ (.A(_01025_),
    .B(\sq.out[14] ),
    .Y(_01208_));
 sky130_fd_sc_hd__and2_1 _08095_ (.A(_01207_),
    .B(_01208_),
    .X(_01209_));
 sky130_fd_sc_hd__inv_2 _08096_ (.A(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__xor2_1 _08097_ (.A(_01208_),
    .B(_01027_),
    .X(_01211_));
 sky130_fd_sc_hd__xor2_1 _08098_ (.A(_01210_),
    .B(_01211_),
    .X(_01212_));
 sky130_fd_sc_hd__nand2_1 _08099_ (.A(net118),
    .B(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__buf_8 _08100_ (.A(_00249_),
    .X(\sq.out[16] ));
 sky130_fd_sc_hd__nand3_1 _08101_ (.A(_01205_),
    .B(_01213_),
    .C(\sq.out[16] ),
    .Y(_01214_));
 sky130_fd_sc_hd__clkinvlp_2 _08102_ (.A(_01002_),
    .Y(_01215_));
 sky130_fd_sc_hd__nand3_2 _08103_ (.A(_01091_),
    .B(_01097_),
    .C(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__clkinvlp_2 _08104_ (.A(_01212_),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_1 _08105_ (.A(_01110_),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__nand3_1 _08106_ (.A(_01216_),
    .B(_01218_),
    .C(_00091_),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_1 _08107_ (.A(_01214_),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand3_1 _08108_ (.A(_01090_),
    .B(_01096_),
    .C(_01206_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_1 _08109_ (.A(_01109_),
    .B(_01209_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand3_2 _08110_ (.A(_01221_),
    .B(_01222_),
    .C(\sq.out[15] ),
    .Y(_01224_));
 sky130_fd_sc_hd__inv_2 _08111_ (.A(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_1 _08112_ (.A(_01220_),
    .B(_01225_),
    .Y(_01226_));
 sky130_fd_sc_hd__nand3_1 _08113_ (.A(_01224_),
    .B(_01214_),
    .C(_01219_),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_1 _08114_ (.A(_01226_),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__inv_2 _08115_ (.A(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _08116_ (.A(_00991_),
    .B(_00992_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand3_1 _08117_ (.A(_01091_),
    .B(_01097_),
    .C(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__xor2_2 _08118_ (.A(_01007_),
    .B(_01028_),
    .X(_01232_));
 sky130_fd_sc_hd__clkinvlp_2 _08119_ (.A(_01232_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _08120_ (.A(_01109_),
    .B(_01233_),
    .Y(_01235_));
 sky130_fd_sc_hd__nand3_2 _08121_ (.A(_01231_),
    .B(_01235_),
    .C(\sq.out[17] ),
    .Y(_01236_));
 sky130_fd_sc_hd__inv_2 _08122_ (.A(_01230_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand3_1 _08123_ (.A(_01091_),
    .B(_01097_),
    .C(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__nand2_1 _08124_ (.A(\sq.out[12] ),
    .B(_01232_),
    .Y(_01239_));
 sky130_fd_sc_hd__buf_6 _08125_ (.A(_00194_),
    .X(_01240_));
 sky130_fd_sc_hd__nand3_1 _08126_ (.A(_01238_),
    .B(_01239_),
    .C(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__nand2_1 _08127_ (.A(_01236_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__nand3_2 _08128_ (.A(_01216_),
    .B(_01218_),
    .C(\sq.out[16] ),
    .Y(_01243_));
 sky130_fd_sc_hd__clkinvlp_2 _08129_ (.A(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand2_1 _08130_ (.A(_01242_),
    .B(_01244_),
    .Y(_01246_));
 sky130_fd_sc_hd__nand3_1 _08131_ (.A(_01236_),
    .B(_01243_),
    .C(_01241_),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2_1 _08132_ (.A(_01246_),
    .B(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__nand2_1 _08133_ (.A(_01229_),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand3_1 _08134_ (.A(_01091_),
    .B(_01097_),
    .C(_00978_),
    .Y(_01250_));
 sky130_fd_sc_hd__a21boi_1 _08135_ (.A1(_01028_),
    .A2(_01005_),
    .B1_N(_01006_),
    .Y(_01251_));
 sky130_fd_sc_hd__xor2_1 _08136_ (.A(_01021_),
    .B(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__nand2_1 _08137_ (.A(_01109_),
    .B(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand3_1 _08138_ (.A(_01250_),
    .B(_01253_),
    .C(_00214_),
    .Y(_01254_));
 sky130_fd_sc_hd__clkinvlp_2 _08139_ (.A(_00978_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand3_1 _08140_ (.A(_01091_),
    .B(_01097_),
    .C(_01255_),
    .Y(_01257_));
 sky130_fd_sc_hd__inv_2 _08141_ (.A(_01252_),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _08142_ (.A(net118),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand3_1 _08143_ (.A(_01257_),
    .B(_01259_),
    .C(_06002_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_1 _08144_ (.A(_01254_),
    .B(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__inv_2 _08145_ (.A(_01236_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand2_1 _08146_ (.A(_01261_),
    .B(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__nand3_2 _08147_ (.A(_01254_),
    .B(_01236_),
    .C(_01260_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand2_1 _08148_ (.A(_01263_),
    .B(_01264_),
    .Y(_01265_));
 sky130_fd_sc_hd__inv_2 _08149_ (.A(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _08150_ (.A(_01129_),
    .B(_01133_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_1 _08151_ (.A(_01267_),
    .B(\sq.out[19] ),
    .Y(_01268_));
 sky130_fd_sc_hd__nand3_1 _08152_ (.A(_01129_),
    .B(_01133_),
    .C(_05130_),
    .Y(_01269_));
 sky130_fd_sc_hd__nand2_1 _08153_ (.A(_01268_),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__nand2_1 _08154_ (.A(_01250_),
    .B(_01253_),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_2 _08155_ (.A(_00214_),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__inv_2 _08156_ (.A(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand2_1 _08157_ (.A(_01270_),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2_1 _08158_ (.A(_01267_),
    .B(_05130_),
    .Y(_01275_));
 sky130_fd_sc_hd__nand2_1 _08159_ (.A(_01275_),
    .B(_01134_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand2_1 _08160_ (.A(_01276_),
    .B(_01272_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2_1 _08161_ (.A(_01274_),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__nand2_1 _08162_ (.A(_01266_),
    .B(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_1 _08163_ (.A(_01249_),
    .B(_01280_),
    .Y(_01281_));
 sky130_fd_sc_hd__nand2_1 _08164_ (.A(\sq.out[12] ),
    .B(_00842_),
    .Y(_01282_));
 sky130_fd_sc_hd__nand2_1 _08165_ (.A(\sq.out[13] ),
    .B(_00749_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_1 _08166_ (.A(_01282_),
    .B(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(_01221_),
    .B(_01222_),
    .Y(_01285_));
 sky130_fd_sc_hd__buf_6 _08168_ (.A(_00425_),
    .X(_01286_));
 sky130_fd_sc_hd__nand2_1 _08169_ (.A(_01285_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__nand2_1 _08170_ (.A(_01287_),
    .B(_01224_),
    .Y(_01288_));
 sky130_fd_sc_hd__or2_1 _08171_ (.A(_01284_),
    .B(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__buf_6 _08172_ (.A(_01289_),
    .X(_01290_));
 sky130_fd_sc_hd__nand3_2 _08173_ (.A(_01204_),
    .B(_01281_),
    .C(_01290_),
    .Y(_01291_));
 sky130_fd_sc_hd__nand2_1 _08174_ (.A(_01191_),
    .B(_01170_),
    .Y(_01292_));
 sky130_fd_sc_hd__nand2_1 _08175_ (.A(_01199_),
    .B(_01192_),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_1 _08176_ (.A(_01292_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__nor2_1 _08177_ (.A(_01176_),
    .B(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__nor2_1 _08178_ (.A(_01153_),
    .B(_01152_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand2_1 _08179_ (.A(_01152_),
    .B(_01153_),
    .Y(_01297_));
 sky130_fd_sc_hd__o21ai_1 _08180_ (.A1(_01137_),
    .A2(_01296_),
    .B1(_01297_),
    .Y(_01299_));
 sky130_fd_sc_hd__inv_2 _08181_ (.A(_01293_),
    .Y(_01300_));
 sky130_fd_sc_hd__o21ai_1 _08182_ (.A1(_01173_),
    .A2(_01300_),
    .B1(_01292_),
    .Y(_01301_));
 sky130_fd_sc_hd__a21oi_1 _08183_ (.A1(_01295_),
    .A2(_01299_),
    .B1(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__nor2_1 _08184_ (.A(_01243_),
    .B(_01242_),
    .Y(_01303_));
 sky130_fd_sc_hd__nand2_1 _08185_ (.A(_01242_),
    .B(_01243_),
    .Y(_01304_));
 sky130_fd_sc_hd__o21ai_1 _08186_ (.A1(_01227_),
    .A2(_01303_),
    .B1(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_1 _08187_ (.A(_01276_),
    .B(_01273_),
    .Y(_01306_));
 sky130_fd_sc_hd__nand2_1 _08188_ (.A(_01270_),
    .B(_01272_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _08189_ (.A(_01306_),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_2 _08190_ (.A(_01265_),
    .B(_01308_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand2_1 _08191_ (.A(_01305_),
    .B(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__nor2_1 _08192_ (.A(_01273_),
    .B(_01276_),
    .Y(_01312_));
 sky130_fd_sc_hd__o21a_1 _08193_ (.A1(_01264_),
    .A2(_01312_),
    .B1(_01306_),
    .X(_01313_));
 sky130_fd_sc_hd__nand2_1 _08194_ (.A(_01311_),
    .B(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__nand2_1 _08195_ (.A(_01314_),
    .B(_01204_),
    .Y(_01315_));
 sky130_fd_sc_hd__nand3_4 _08196_ (.A(_01291_),
    .B(_01302_),
    .C(_01315_),
    .Y(_01316_));
 sky130_fd_sc_hd__nand2_1 _08197_ (.A(_01086_),
    .B(_01087_),
    .Y(_01317_));
 sky130_fd_sc_hd__inv_4 _08198_ (.A(_01317_),
    .Y(_01318_));
 sky130_fd_sc_hd__or2_1 _08199_ (.A(_01318_),
    .B(_01049_),
    .X(_01319_));
 sky130_fd_sc_hd__nand2_1 _08200_ (.A(_01049_),
    .B(_01318_),
    .Y(_01321_));
 sky130_fd_sc_hd__a21o_1 _08201_ (.A1(_01319_),
    .A2(_01321_),
    .B1(_01186_),
    .X(_01322_));
 sky130_fd_sc_hd__nand2_1 _08202_ (.A(_01186_),
    .B(_01075_),
    .Y(_01323_));
 sky130_fd_sc_hd__nand2_1 _08203_ (.A(_01322_),
    .B(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hd__inv_2 _08204_ (.A(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__nand2_1 _08205_ (.A(_01321_),
    .B(_01087_),
    .Y(_01326_));
 sky130_fd_sc_hd__or2_1 _08206_ (.A(_01079_),
    .B(_01326_),
    .X(_01327_));
 sky130_fd_sc_hd__nand2_1 _08207_ (.A(_01326_),
    .B(_01079_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand3_1 _08208_ (.A(_01327_),
    .B(\sq.out[12] ),
    .C(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__nand2_1 _08209_ (.A(_01186_),
    .B(_01058_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _08210_ (.A(_01329_),
    .B(_01330_),
    .Y(_01332_));
 sky130_fd_sc_hd__or2_1 _08211_ (.A(_01325_),
    .B(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__a31o_1 _08212_ (.A1(_01049_),
    .A2(_01079_),
    .A3(_01318_),
    .B1(_01094_),
    .X(_01334_));
 sky130_fd_sc_hd__nand3_2 _08213_ (.A(_01334_),
    .B(_01064_),
    .C(_01058_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_1 _08214_ (.A(_01332_),
    .B(_01325_),
    .Y(_01336_));
 sky130_fd_sc_hd__nand3_1 _08215_ (.A(_01333_),
    .B(_01335_),
    .C(_01336_),
    .Y(_01337_));
 sky130_fd_sc_hd__inv_2 _08216_ (.A(_01337_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_01181_),
    .B(_00921_),
    .Y(_01339_));
 sky130_fd_sc_hd__or2_1 _08218_ (.A(_00949_),
    .B(_01339_),
    .X(_01340_));
 sky130_fd_sc_hd__nand2_1 _08219_ (.A(_01339_),
    .B(_00949_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand3_2 _08220_ (.A(_01340_),
    .B(net118),
    .C(_01341_),
    .Y(_01343_));
 sky130_fd_sc_hd__buf_6 _08221_ (.A(_00283_),
    .X(_01344_));
 sky130_fd_sc_hd__or2_4 _08222_ (.A(_00934_),
    .B(net118),
    .X(_01345_));
 sky130_fd_sc_hd__nand3_1 _08223_ (.A(_01343_),
    .B(_01344_),
    .C(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__nor2_1 _08224_ (.A(_01324_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__nand2_2 _08225_ (.A(_01346_),
    .B(_01324_),
    .Y(_01348_));
 sky130_fd_sc_hd__inv_2 _08226_ (.A(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__or2_1 _08227_ (.A(_01347_),
    .B(_01349_),
    .X(_01350_));
 sky130_fd_sc_hd__a21o_1 _08228_ (.A1(_01343_),
    .A2(_01345_),
    .B1(_01344_),
    .X(_01351_));
 sky130_fd_sc_hd__nand3b_1 _08229_ (.A_N(_01189_),
    .B(_01351_),
    .C(_01346_),
    .Y(_01352_));
 sky130_fd_sc_hd__a21o_1 _08230_ (.A1(_01343_),
    .A2(_01345_),
    .B1(_01081_),
    .X(_01354_));
 sky130_fd_sc_hd__nand3_1 _08231_ (.A(_01343_),
    .B(_01081_),
    .C(_01345_),
    .Y(_01355_));
 sky130_fd_sc_hd__nand3_2 _08232_ (.A(_01354_),
    .B(_01189_),
    .C(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(_01352_),
    .B(_01356_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_2 _08234_ (.A(_01350_),
    .B(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__nand3_4 _08235_ (.A(_01316_),
    .B(_01338_),
    .C(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__o21ai_2 _08236_ (.A1(_01347_),
    .A2(_01356_),
    .B1(_01348_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _08237_ (.A(_01336_),
    .B(_01335_),
    .Y(_01361_));
 sky130_fd_sc_hd__a21oi_4 _08238_ (.A1(_01360_),
    .A2(_01338_),
    .B1(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__buf_6 _08239_ (.A(_01186_),
    .X(_01363_));
 sky130_fd_sc_hd__nand3_2 _08240_ (.A(net98),
    .B(_01362_),
    .C(_01363_),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_2 _08241_ (.A(_01359_),
    .B(_01362_),
    .Y(_01366_));
 sky130_fd_sc_hd__buf_6 _08242_ (.A(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__buf_6 _08243_ (.A(_01367_),
    .X(_01368_));
 sky130_fd_sc_hd__nand2_1 _08244_ (.A(_00842_),
    .B(\sq.out[14] ),
    .Y(_01369_));
 sky130_fd_sc_hd__nand2_1 _08245_ (.A(_01369_),
    .B(_01283_),
    .Y(_01370_));
 sky130_fd_sc_hd__nand2_1 _08246_ (.A(_01368_),
    .B(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__o21ai_2 _08247_ (.A1(\sq.out[13] ),
    .A2(_01365_),
    .B1(_01371_),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_2 _08248_ (.A(_01372_),
    .B(\sq.out[15] ),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_1 _08249_ (.A(_01288_),
    .B(_01284_),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _08250_ (.A(_01290_),
    .B(_01374_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _08251_ (.A(_01367_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand3_1 _08252_ (.A(_01359_),
    .B(_01362_),
    .C(_01285_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _08253_ (.A(_01377_),
    .B(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__nand2_1 _08254_ (.A(_01379_),
    .B(_00091_),
    .Y(_01380_));
 sky130_fd_sc_hd__nand3_1 _08255_ (.A(_01377_),
    .B(\sq.out[16] ),
    .C(_01378_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_1 _08256_ (.A(_01380_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand2_1 _08257_ (.A(_01373_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__xor2_1 _08258_ (.A(_01228_),
    .B(_01290_),
    .X(_01384_));
 sky130_fd_sc_hd__inv_2 _08259_ (.A(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_1 _08260_ (.A(_01367_),
    .B(_01385_),
    .Y(_01387_));
 sky130_fd_sc_hd__nand2_1 _08261_ (.A(_01216_),
    .B(_01218_),
    .Y(_01388_));
 sky130_fd_sc_hd__nand3_1 _08262_ (.A(_01359_),
    .B(_01362_),
    .C(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__nand2_1 _08263_ (.A(_01387_),
    .B(_01389_),
    .Y(_01390_));
 sky130_fd_sc_hd__nand2_1 _08264_ (.A(_01390_),
    .B(_01240_),
    .Y(_01391_));
 sky130_fd_sc_hd__nand3_1 _08265_ (.A(_01387_),
    .B(\sq.out[17] ),
    .C(_01389_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand2_1 _08266_ (.A(_01391_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _08267_ (.A(_01381_),
    .B(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__nand2_1 _08268_ (.A(_01393_),
    .B(_01381_),
    .Y(_01395_));
 sky130_fd_sc_hd__o21ai_1 _08269_ (.A1(_01383_),
    .A2(_01394_),
    .B1(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand3_1 _08270_ (.A(_01244_),
    .B(_01236_),
    .C(_01241_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand2_1 _08271_ (.A(_01398_),
    .B(_01304_),
    .Y(_01399_));
 sky130_fd_sc_hd__a21boi_1 _08272_ (.A1(_01290_),
    .A2(_01226_),
    .B1_N(_01227_),
    .Y(_01400_));
 sky130_fd_sc_hd__xor2_1 _08273_ (.A(_01399_),
    .B(_01400_),
    .X(_01401_));
 sky130_fd_sc_hd__nand2_1 _08274_ (.A(_01367_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__nand2_1 _08275_ (.A(_01231_),
    .B(_01235_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand3_1 _08276_ (.A(net98),
    .B(_01362_),
    .C(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _08277_ (.A(_01402_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand2_1 _08278_ (.A(_01405_),
    .B(_00214_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand3_2 _08279_ (.A(_01402_),
    .B(_06002_),
    .C(_01404_),
    .Y(_01407_));
 sky130_fd_sc_hd__nand2_1 _08280_ (.A(_01406_),
    .B(_01407_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2_1 _08281_ (.A(_01409_),
    .B(_01392_),
    .Y(_01410_));
 sky130_fd_sc_hd__inv_2 _08282_ (.A(_01392_),
    .Y(_01411_));
 sky130_fd_sc_hd__nand3_1 _08283_ (.A(_01411_),
    .B(_01406_),
    .C(_01407_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _08284_ (.A(_01410_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_1 _08285_ (.A(_01228_),
    .B(_01399_),
    .Y(_01414_));
 sky130_fd_sc_hd__a21o_1 _08286_ (.A1(_01414_),
    .A2(_01290_),
    .B1(_01305_),
    .X(_01415_));
 sky130_fd_sc_hd__or2_1 _08287_ (.A(_01266_),
    .B(_01415_),
    .X(_01416_));
 sky130_fd_sc_hd__nand2_1 _08288_ (.A(_01415_),
    .B(_01266_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_1 _08289_ (.A(_01416_),
    .B(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__inv_2 _08290_ (.A(_01418_),
    .Y(_01420_));
 sky130_fd_sc_hd__nand2_1 _08291_ (.A(_01367_),
    .B(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__nand3_1 _08292_ (.A(_01359_),
    .B(_01362_),
    .C(_01271_),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _08293_ (.A(_01421_),
    .B(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _08294_ (.A(_01423_),
    .B(_05130_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand3_1 _08295_ (.A(_01421_),
    .B(\sq.out[19] ),
    .C(_01422_),
    .Y(_01425_));
 sky130_fd_sc_hd__nand2_1 _08296_ (.A(_01424_),
    .B(_01425_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _08297_ (.A(_01426_),
    .B(_01407_),
    .Y(_01427_));
 sky130_fd_sc_hd__inv_2 _08298_ (.A(_01407_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand3_1 _08299_ (.A(_01428_),
    .B(_01424_),
    .C(_01425_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_1 _08300_ (.A(_01427_),
    .B(_01429_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_1 _08301_ (.A(_01413_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand2_1 _08302_ (.A(_01396_),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__nor2_1 _08303_ (.A(_01407_),
    .B(_01426_),
    .Y(_01434_));
 sky130_fd_sc_hd__o21a_1 _08304_ (.A1(_01410_),
    .A2(_01434_),
    .B1(_01427_),
    .X(_01435_));
 sky130_fd_sc_hd__nand2_1 _08305_ (.A(_01433_),
    .B(_01435_),
    .Y(_01436_));
 sky130_fd_sc_hd__nand2_1 _08306_ (.A(_01417_),
    .B(_01264_),
    .Y(_01437_));
 sky130_fd_sc_hd__xor2_1 _08307_ (.A(_01279_),
    .B(_01437_),
    .X(_01438_));
 sky130_fd_sc_hd__nand2_1 _08308_ (.A(_01438_),
    .B(_01367_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand3_1 _08309_ (.A(net98),
    .B(_01362_),
    .C(_01267_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand3_2 _08310_ (.A(_01439_),
    .B(_00460_),
    .C(_01440_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _08311_ (.A(_01439_),
    .B(_01440_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _08312_ (.A(_01443_),
    .B(_06045_),
    .Y(_01444_));
 sky130_fd_sc_hd__nand3b_1 _08313_ (.A_N(_01425_),
    .B(_01442_),
    .C(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _08314_ (.A(_01444_),
    .B(_01442_),
    .Y(_01446_));
 sky130_fd_sc_hd__nand2_1 _08315_ (.A(_01446_),
    .B(_01425_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _08316_ (.A(_01445_),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__inv_2 _08317_ (.A(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__inv_2 _08318_ (.A(_01442_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand3_1 _08319_ (.A(_01310_),
    .B(_01414_),
    .C(_01290_),
    .Y(_01451_));
 sky130_fd_sc_hd__nand3_1 _08320_ (.A(_01451_),
    .B(_01313_),
    .C(_01311_),
    .Y(_01453_));
 sky130_fd_sc_hd__or2_1 _08321_ (.A(_01139_),
    .B(_01453_),
    .X(_01454_));
 sky130_fd_sc_hd__nand2_1 _08322_ (.A(_01453_),
    .B(_01139_),
    .Y(_01455_));
 sky130_fd_sc_hd__nand2_1 _08323_ (.A(_01454_),
    .B(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__inv_2 _08324_ (.A(_01456_),
    .Y(_01457_));
 sky130_fd_sc_hd__nand2_1 _08325_ (.A(_01367_),
    .B(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__nand3_1 _08326_ (.A(net98),
    .B(_01362_),
    .C(_01124_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand2_1 _08327_ (.A(_01458_),
    .B(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _08328_ (.A(_01460_),
    .B(_00455_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand3_2 _08329_ (.A(_01458_),
    .B(\sq.out[21] ),
    .C(_01459_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand3_1 _08330_ (.A(_01450_),
    .B(_01461_),
    .C(_01462_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _08331_ (.A(_01461_),
    .B(_01462_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand2_1 _08332_ (.A(_01465_),
    .B(_01442_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_1 _08333_ (.A(_01464_),
    .B(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__inv_2 _08334_ (.A(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _08335_ (.A(_01449_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__inv_2 _08336_ (.A(_01158_),
    .Y(_01470_));
 sky130_fd_sc_hd__nand2_1 _08337_ (.A(_01453_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__inv_2 _08338_ (.A(_01299_),
    .Y(_01472_));
 sky130_fd_sc_hd__nand2_1 _08339_ (.A(_01471_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__or2b_1 _08340_ (.A(_01473_),
    .B_N(_01176_),
    .X(_01475_));
 sky130_fd_sc_hd__nand2_1 _08341_ (.A(_01473_),
    .B(_01177_),
    .Y(_01476_));
 sky130_fd_sc_hd__nand3_1 _08342_ (.A(_01367_),
    .B(_01475_),
    .C(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__inv_2 _08343_ (.A(_01366_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_1 _08344_ (.A(_01168_),
    .B(_01169_),
    .Y(_01479_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(_01478_),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2_1 _08346_ (.A(_01477_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand2_1 _08347_ (.A(_01481_),
    .B(_00743_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand3_2 _08348_ (.A(_01477_),
    .B(_01480_),
    .C(_00437_),
    .Y(_01483_));
 sky130_fd_sc_hd__nand2_1 _08349_ (.A(_01482_),
    .B(_01483_),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _08350_ (.A(_01455_),
    .B(_01137_),
    .Y(_01486_));
 sky130_fd_sc_hd__nand2_1 _08351_ (.A(_01486_),
    .B(_01157_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand3b_1 _08352_ (.A_N(_01157_),
    .B(_01455_),
    .C(_01137_),
    .Y(_01488_));
 sky130_fd_sc_hd__nand2_1 _08353_ (.A(_01487_),
    .B(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_01367_),
    .B(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hd__nand3b_1 _08355_ (.A_N(_01148_),
    .B(_01359_),
    .C(_01362_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _08356_ (.A(_01490_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_2 _08357_ (.A(_01492_),
    .B(_00177_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand2_1 _08358_ (.A(_01484_),
    .B(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hd__inv_2 _08359_ (.A(_01493_),
    .Y(_01495_));
 sky130_fd_sc_hd__nand3_1 _08360_ (.A(_01482_),
    .B(_01495_),
    .C(_01483_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand2_2 _08361_ (.A(_01494_),
    .B(_01497_),
    .Y(_01498_));
 sky130_fd_sc_hd__inv_2 _08362_ (.A(_01498_),
    .Y(_01499_));
 sky130_fd_sc_hd__nand3_1 _08363_ (.A(_01490_),
    .B(_01491_),
    .C(_06106_),
    .Y(_01500_));
 sky130_fd_sc_hd__nand3b_1 _08364_ (.A_N(_01462_),
    .B(_01493_),
    .C(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__nand2_1 _08365_ (.A(_01493_),
    .B(_01500_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand2_2 _08366_ (.A(_01502_),
    .B(_01462_),
    .Y(_01503_));
 sky130_fd_sc_hd__nand2_2 _08367_ (.A(_01501_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__inv_2 _08368_ (.A(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__nand2_1 _08369_ (.A(_01499_),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_2 _08370_ (.A(_01469_),
    .B(_01506_),
    .Y(_01508_));
 sky130_fd_sc_hd__nand2_1 _08371_ (.A(_01436_),
    .B(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__nor2_1 _08372_ (.A(_01504_),
    .B(_01498_),
    .Y(_01510_));
 sky130_fd_sc_hd__nor2_1 _08373_ (.A(_01442_),
    .B(_01465_),
    .Y(_01511_));
 sky130_fd_sc_hd__o21ai_2 _08374_ (.A1(_01447_),
    .A2(_01511_),
    .B1(_01466_),
    .Y(_01512_));
 sky130_fd_sc_hd__inv_2 _08375_ (.A(_01497_),
    .Y(_01513_));
 sky130_fd_sc_hd__o21ai_1 _08376_ (.A1(_01503_),
    .A2(_01513_),
    .B1(_01494_),
    .Y(_01514_));
 sky130_fd_sc_hd__a21oi_1 _08377_ (.A1(_01510_),
    .A2(_01512_),
    .B1(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__nand2_1 _08378_ (.A(_01509_),
    .B(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand2_1 _08379_ (.A(_01316_),
    .B(_01358_),
    .Y(_01517_));
 sky130_fd_sc_hd__inv_2 _08380_ (.A(_01360_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _08381_ (.A(_01333_),
    .B(_01336_),
    .Y(_01520_));
 sky130_fd_sc_hd__a21o_1 _08382_ (.A1(_01517_),
    .A2(_01519_),
    .B1(_01520_),
    .X(_01521_));
 sky130_fd_sc_hd__nand3_1 _08383_ (.A(_01521_),
    .B(_01336_),
    .C(_01368_),
    .Y(_01522_));
 sky130_fd_sc_hd__xnor2_2 _08384_ (.A(_01335_),
    .B(_01522_),
    .Y(_01523_));
 sky130_fd_sc_hd__inv_2 _08385_ (.A(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand2_1 _08386_ (.A(_01476_),
    .B(_01173_),
    .Y(_01525_));
 sky130_fd_sc_hd__nand2_1 _08387_ (.A(_01525_),
    .B(_01201_),
    .Y(_01526_));
 sky130_fd_sc_hd__nand3_1 _08388_ (.A(_01476_),
    .B(_01294_),
    .C(_01173_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand2_1 _08389_ (.A(_01526_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__nand2_1 _08390_ (.A(_01528_),
    .B(_01368_),
    .Y(_01530_));
 sky130_fd_sc_hd__buf_6 _08391_ (.A(_01478_),
    .X(_01531_));
 sky130_fd_sc_hd__nand2_1 _08392_ (.A(_01531_),
    .B(_01188_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _08393_ (.A(_01530_),
    .B(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__nand2_1 _08394_ (.A(_01533_),
    .B(_01344_),
    .Y(_01534_));
 sky130_fd_sc_hd__a21o_1 _08395_ (.A1(_01343_),
    .A2(_01345_),
    .B1(_01367_),
    .X(_01535_));
 sky130_fd_sc_hd__inv_2 _08396_ (.A(_01357_),
    .Y(_01536_));
 sky130_fd_sc_hd__nand2_1 _08397_ (.A(_01316_),
    .B(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__or2_1 _08398_ (.A(_01536_),
    .B(_01316_),
    .X(_01538_));
 sky130_fd_sc_hd__nand3_1 _08399_ (.A(_01368_),
    .B(_01537_),
    .C(_01538_),
    .Y(_01539_));
 sky130_fd_sc_hd__nand2_2 _08400_ (.A(_01535_),
    .B(_01539_),
    .Y(_01541_));
 sky130_fd_sc_hd__inv_2 _08401_ (.A(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2_1 _08402_ (.A(_01534_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__nand3_1 _08403_ (.A(_01533_),
    .B(_01541_),
    .C(_01344_),
    .Y(_01544_));
 sky130_fd_sc_hd__nand2_1 _08404_ (.A(_01543_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand3_1 _08405_ (.A(_01530_),
    .B(_01081_),
    .C(_01532_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_1 _08406_ (.A(_01534_),
    .B(_01546_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand2_1 _08407_ (.A(_01547_),
    .B(_01483_),
    .Y(_01548_));
 sky130_fd_sc_hd__nand3b_1 _08408_ (.A_N(_01483_),
    .B(_01534_),
    .C(_01546_),
    .Y(_01549_));
 sky130_fd_sc_hd__nand2_1 _08409_ (.A(_01548_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__nor2_2 _08410_ (.A(_01545_),
    .B(_01550_),
    .Y(_01552_));
 sky130_fd_sc_hd__clkinvlp_2 _08411_ (.A(_01350_),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_1 _08412_ (.A(_01537_),
    .B(_01356_),
    .Y(_01554_));
 sky130_fd_sc_hd__or2_1 _08413_ (.A(_01553_),
    .B(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__nand2_1 _08414_ (.A(_01554_),
    .B(_01553_),
    .Y(_01556_));
 sky130_fd_sc_hd__nand3_1 _08415_ (.A(_01555_),
    .B(_01368_),
    .C(_01556_),
    .Y(_01557_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(_01531_),
    .B(_01325_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_1 _08417_ (.A(_01557_),
    .B(_01558_),
    .Y(_01559_));
 sky130_fd_sc_hd__or2_1 _08418_ (.A(_01541_),
    .B(_01559_),
    .X(_01560_));
 sky130_fd_sc_hd__nand2_1 _08419_ (.A(_01559_),
    .B(_01541_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand3_1 _08420_ (.A(_01517_),
    .B(_01520_),
    .C(_01519_),
    .Y(_01563_));
 sky130_fd_sc_hd__nand2_1 _08421_ (.A(_01521_),
    .B(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__nand2_1 _08422_ (.A(_01531_),
    .B(_01332_),
    .Y(_01565_));
 sky130_fd_sc_hd__o21ai_1 _08423_ (.A1(_01531_),
    .A2(_01564_),
    .B1(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__inv_4 _08424_ (.A(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__nand3_1 _08425_ (.A(_01560_),
    .B(_01561_),
    .C(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__inv_2 _08426_ (.A(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__nand2_2 _08427_ (.A(_01552_),
    .B(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__nor2_4 _08428_ (.A(_01524_),
    .B(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__o21ai_1 _08429_ (.A1(_01545_),
    .A2(_01548_),
    .B1(_01543_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_1 _08430_ (.A(_01572_),
    .B(_01569_),
    .Y(_01574_));
 sky130_fd_sc_hd__and2_1 _08431_ (.A(_01567_),
    .B(_01561_),
    .X(_01575_));
 sky130_fd_sc_hd__nand3_1 _08432_ (.A(_01574_),
    .B(_01523_),
    .C(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__a21oi_4 _08433_ (.A1(_01516_),
    .A2(_01571_),
    .B1(_01576_),
    .Y(_01577_));
 sky130_fd_sc_hd__clkinvlp_2 _08434_ (.A(_01432_),
    .Y(_01578_));
 sky130_fd_sc_hd__nor3_1 _08435_ (.A(\sq.out[14] ),
    .B(_00843_),
    .C(_01365_),
    .Y(_01579_));
 sky130_fd_sc_hd__nand2_1 _08436_ (.A(_01363_),
    .B(\sq.out[13] ),
    .Y(_01580_));
 sky130_fd_sc_hd__nand2_2 _08437_ (.A(_01580_),
    .B(_01282_),
    .Y(_01581_));
 sky130_fd_sc_hd__a21oi_1 _08438_ (.A1(_01368_),
    .A2(_00843_),
    .B1(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__nand2_1 _08439_ (.A(_01368_),
    .B(_01581_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _08440_ (.A(_01583_),
    .B(_01365_),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _08441_ (.A(_01585_),
    .B(\sq.out[14] ),
    .Y(_01586_));
 sky130_fd_sc_hd__buf_6 _08442_ (.A(_00749_),
    .X(_01587_));
 sky130_fd_sc_hd__nand3_1 _08443_ (.A(_01583_),
    .B(_01587_),
    .C(_01365_),
    .Y(_01588_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_01586_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__or2_1 _08445_ (.A(_00843_),
    .B(_01365_),
    .X(_01590_));
 sky130_fd_sc_hd__nand2_1 _08446_ (.A(_01589_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__o21ai_2 _08447_ (.A1(_01579_),
    .A2(_01582_),
    .B1(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__nand3_1 _08448_ (.A(_01531_),
    .B(_00843_),
    .C(_01363_),
    .Y(_01593_));
 sky130_fd_sc_hd__nand3_1 _08449_ (.A(_01593_),
    .B(_01286_),
    .C(_01371_),
    .Y(_01594_));
 sky130_fd_sc_hd__nand2_1 _08450_ (.A(_01373_),
    .B(_01594_),
    .Y(_01596_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(_01596_),
    .B(_01586_),
    .Y(_01597_));
 sky130_fd_sc_hd__nand3b_1 _08452_ (.A_N(_01586_),
    .B(_01373_),
    .C(_01594_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand3_2 _08453_ (.A(_01592_),
    .B(_01597_),
    .C(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand2_2 _08454_ (.A(_01599_),
    .B(_01597_),
    .Y(_01600_));
 sky130_fd_sc_hd__or2b_1 _08455_ (.A(_01394_),
    .B_N(_01395_),
    .X(_01601_));
 sky130_fd_sc_hd__inv_2 _08456_ (.A(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__or2_1 _08457_ (.A(_01382_),
    .B(_01373_),
    .X(_01603_));
 sky130_fd_sc_hd__and2_1 _08458_ (.A(_01603_),
    .B(_01383_),
    .X(_01604_));
 sky130_fd_sc_hd__nand3_2 _08459_ (.A(_01600_),
    .B(_01602_),
    .C(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_4 _08460_ (.A(_01578_),
    .B(_01605_),
    .Y(_01607_));
 sky130_fd_sc_hd__nand3_4 _08461_ (.A(_01607_),
    .B(_01571_),
    .C(_01508_),
    .Y(_01608_));
 sky130_fd_sc_hd__nand2_4 _08462_ (.A(_01608_),
    .B(_01577_),
    .Y(_01609_));
 sky130_fd_sc_hd__buf_6 _08463_ (.A(_01609_),
    .X(_01610_));
 sky130_fd_sc_hd__inv_2 _08464_ (.A(_01581_),
    .Y(_01611_));
 sky130_fd_sc_hd__nand2_1 _08465_ (.A(_01610_),
    .B(_01611_),
    .Y(_01612_));
 sky130_fd_sc_hd__nand3_1 _08466_ (.A(_01577_),
    .B(_01365_),
    .C(_01608_),
    .Y(_01613_));
 sky130_fd_sc_hd__nand2_1 _08467_ (.A(_01612_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__nand2_1 _08468_ (.A(_01614_),
    .B(_01587_),
    .Y(_01615_));
 sky130_fd_sc_hd__nand3_1 _08469_ (.A(_01612_),
    .B(\sq.out[14] ),
    .C(_01613_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _08470_ (.A(_01615_),
    .B(_01616_),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _08471_ (.A(_01531_),
    .B(\sq.out[12] ),
    .Y(_01619_));
 sky130_fd_sc_hd__nand2_1 _08472_ (.A(_01368_),
    .B(_01363_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_1 _08473_ (.A(_01619_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__inv_2 _08474_ (.A(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _08475_ (.A(_01610_),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__nand3_2 _08476_ (.A(_01577_),
    .B(_01368_),
    .C(_01608_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand3_2 _08477_ (.A(_01623_),
    .B(\sq.out[13] ),
    .C(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__nand2_1 _08478_ (.A(_01618_),
    .B(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__clkinvlp_2 _08479_ (.A(_01625_),
    .Y(_01627_));
 sky130_fd_sc_hd__nand3_1 _08480_ (.A(_01627_),
    .B(_01615_),
    .C(_01616_),
    .Y(_01629_));
 sky130_fd_sc_hd__nand2_1 _08481_ (.A(_01623_),
    .B(_01624_),
    .Y(_01630_));
 sky130_fd_sc_hd__nand2_1 _08482_ (.A(_01630_),
    .B(_00843_),
    .Y(_01631_));
 sky130_fd_sc_hd__buf_6 _08483_ (.A(_01610_),
    .X(_01632_));
 sky130_fd_sc_hd__nand2_1 _08484_ (.A(_01632_),
    .B(_01531_),
    .Y(_01633_));
 sky130_fd_sc_hd__and2_1 _08485_ (.A(_01633_),
    .B(_01620_),
    .X(_01634_));
 sky130_fd_sc_hd__nand3_2 _08486_ (.A(_01631_),
    .B(_01634_),
    .C(_01625_),
    .Y(_01635_));
 sky130_fd_sc_hd__nand3_1 _08487_ (.A(_01626_),
    .B(_01629_),
    .C(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(_01636_),
    .B(_01626_),
    .Y(_01637_));
 sky130_fd_sc_hd__or2b_1 _08489_ (.A(_01579_),
    .B_N(_01591_),
    .X(_01638_));
 sky130_fd_sc_hd__or2_1 _08490_ (.A(_01582_),
    .B(_01638_),
    .X(_01640_));
 sky130_fd_sc_hd__nand2_1 _08491_ (.A(_01638_),
    .B(_01582_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand3_1 _08492_ (.A(_01610_),
    .B(_01640_),
    .C(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__inv_2 _08493_ (.A(_01609_),
    .Y(_01643_));
 sky130_fd_sc_hd__buf_6 _08494_ (.A(_01643_),
    .X(_01644_));
 sky130_fd_sc_hd__inv_2 _08495_ (.A(_01585_),
    .Y(_01645_));
 sky130_fd_sc_hd__nand2_1 _08496_ (.A(_01644_),
    .B(_01645_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _08497_ (.A(_01642_),
    .B(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _08498_ (.A(_01647_),
    .B(_01286_),
    .Y(_01648_));
 sky130_fd_sc_hd__nand3_2 _08499_ (.A(_01642_),
    .B(_01646_),
    .C(\sq.out[15] ),
    .Y(_01649_));
 sky130_fd_sc_hd__nand2_1 _08500_ (.A(_01648_),
    .B(_01649_),
    .Y(_01651_));
 sky130_fd_sc_hd__nand2_1 _08501_ (.A(_01651_),
    .B(_01616_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand3b_1 _08502_ (.A_N(_01616_),
    .B(_01648_),
    .C(_01649_),
    .Y(_01653_));
 sky130_fd_sc_hd__nand2_1 _08503_ (.A(_01652_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__inv_2 _08504_ (.A(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_1 _08505_ (.A(_01637_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _08506_ (.A(_01656_),
    .B(_01652_),
    .Y(_01657_));
 sky130_fd_sc_hd__a21o_1 _08507_ (.A1(_01597_),
    .A2(_01598_),
    .B1(_01592_),
    .X(_01658_));
 sky130_fd_sc_hd__nand3_1 _08508_ (.A(_01609_),
    .B(_01599_),
    .C(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand3b_1 _08509_ (.A_N(_01372_),
    .B(_01577_),
    .C(_01608_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _08510_ (.A(_01659_),
    .B(_01660_),
    .Y(_01662_));
 sky130_fd_sc_hd__inv_2 _08511_ (.A(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand2_1 _08512_ (.A(_01663_),
    .B(\sq.out[16] ),
    .Y(_01664_));
 sky130_fd_sc_hd__nand2_1 _08513_ (.A(_01600_),
    .B(_01604_),
    .Y(_01665_));
 sky130_fd_sc_hd__or2_1 _08514_ (.A(_01604_),
    .B(_01600_),
    .X(_01666_));
 sky130_fd_sc_hd__nand3_1 _08515_ (.A(_01609_),
    .B(_01665_),
    .C(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _08516_ (.A(_01643_),
    .B(_01379_),
    .Y(_01668_));
 sky130_fd_sc_hd__nand2_1 _08517_ (.A(_01667_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__inv_2 _08518_ (.A(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _08519_ (.A(_01670_),
    .B(\sq.out[17] ),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _08520_ (.A(_01669_),
    .B(_01240_),
    .Y(_01673_));
 sky130_fd_sc_hd__nand2_1 _08521_ (.A(_01671_),
    .B(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__nor2_1 _08522_ (.A(_01664_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_1 _08523_ (.A(_01674_),
    .B(_01664_),
    .Y(_01676_));
 sky130_fd_sc_hd__or2b_1 _08524_ (.A(_01675_),
    .B_N(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__inv_2 _08525_ (.A(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(_01662_),
    .B(_00091_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _08527_ (.A(_01664_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__or2_1 _08528_ (.A(_01649_),
    .B(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(_01680_),
    .B(_01649_),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2_1 _08530_ (.A(_01681_),
    .B(_01682_),
    .Y(_01684_));
 sky130_fd_sc_hd__inv_2 _08531_ (.A(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__nand3_1 _08532_ (.A(_01657_),
    .B(_01678_),
    .C(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__o21a_1 _08533_ (.A1(_01682_),
    .A2(_01675_),
    .B1(_01676_),
    .X(_01687_));
 sky130_fd_sc_hd__nand2_1 _08534_ (.A(_01686_),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__nand2_1 _08535_ (.A(_01665_),
    .B(_01383_),
    .Y(_01689_));
 sky130_fd_sc_hd__or2_1 _08536_ (.A(_01602_),
    .B(_01689_),
    .X(_01690_));
 sky130_fd_sc_hd__nand2_1 _08537_ (.A(_01689_),
    .B(_01602_),
    .Y(_01691_));
 sky130_fd_sc_hd__a21o_1 _08538_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01644_),
    .X(_01692_));
 sky130_fd_sc_hd__or2_1 _08539_ (.A(_01390_),
    .B(_01610_),
    .X(_01693_));
 sky130_fd_sc_hd__nand2_1 _08540_ (.A(_01692_),
    .B(_01693_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _08541_ (.A(_01695_),
    .B(_06002_),
    .Y(_01696_));
 sky130_fd_sc_hd__nand2b_1 _08542_ (.A_N(_01396_),
    .B(_01605_),
    .Y(_01697_));
 sky130_fd_sc_hd__nand2b_1 _08543_ (.A_N(_01413_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__or2b_1 _08544_ (.A(_01697_),
    .B_N(_01413_),
    .X(_01699_));
 sky130_fd_sc_hd__nand3_1 _08545_ (.A(_01610_),
    .B(_01698_),
    .C(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__nand2_1 _08546_ (.A(_01643_),
    .B(_01405_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_1 _08547_ (.A(_01700_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__inv_2 _08548_ (.A(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_1 _08549_ (.A(_01703_),
    .B(\sq.out[19] ),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _08550_ (.A(_01702_),
    .B(_05130_),
    .Y(_01706_));
 sky130_fd_sc_hd__nand2_1 _08551_ (.A(_01704_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__or2_1 _08552_ (.A(_01696_),
    .B(_01707_),
    .X(_01708_));
 sky130_fd_sc_hd__nand2_1 _08553_ (.A(_01707_),
    .B(_01696_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_1 _08554_ (.A(_01708_),
    .B(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__inv_2 _08555_ (.A(_01695_),
    .Y(_01711_));
 sky130_fd_sc_hd__buf_6 _08556_ (.A(_00214_),
    .X(_01712_));
 sky130_fd_sc_hd__nand2_1 _08557_ (.A(_01711_),
    .B(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(_01713_),
    .B(_01696_),
    .Y(_01714_));
 sky130_fd_sc_hd__or2_1 _08559_ (.A(_01671_),
    .B(_01714_),
    .X(_01715_));
 sky130_fd_sc_hd__nand2_1 _08560_ (.A(_01714_),
    .B(_01671_),
    .Y(_01717_));
 sky130_fd_sc_hd__nand2_1 _08561_ (.A(_01715_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__nor2_1 _08562_ (.A(_01710_),
    .B(_01718_),
    .Y(_01719_));
 sky130_fd_sc_hd__nand2_1 _08563_ (.A(_01688_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__o21a_1 _08564_ (.A1(_01717_),
    .A2(_01710_),
    .B1(_01709_),
    .X(_01721_));
 sky130_fd_sc_hd__nand2_2 _08565_ (.A(_01720_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__nand2_1 _08566_ (.A(_01698_),
    .B(_01410_),
    .Y(_01723_));
 sky130_fd_sc_hd__xor2_1 _08567_ (.A(_01431_),
    .B(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__nand2_1 _08568_ (.A(_01724_),
    .B(_01632_),
    .Y(_01725_));
 sky130_fd_sc_hd__or2_1 _08569_ (.A(_01423_),
    .B(_01610_),
    .X(_01726_));
 sky130_fd_sc_hd__nand2_1 _08570_ (.A(_01725_),
    .B(_01726_),
    .Y(_01728_));
 sky130_fd_sc_hd__inv_2 _08571_ (.A(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__buf_6 _08572_ (.A(_06045_),
    .X(_01730_));
 sky130_fd_sc_hd__nand2_1 _08573_ (.A(_01729_),
    .B(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__nand2_1 _08574_ (.A(_01728_),
    .B(_00460_),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_1 _08575_ (.A(_01731_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand2_1 _08576_ (.A(_01733_),
    .B(_01704_),
    .Y(_01734_));
 sky130_fd_sc_hd__nand3b_1 _08577_ (.A_N(_01704_),
    .B(_01731_),
    .C(_01732_),
    .Y(_01735_));
 sky130_fd_sc_hd__nand2_1 _08578_ (.A(_01734_),
    .B(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__inv_2 _08579_ (.A(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__or2_1 _08580_ (.A(_01436_),
    .B(_01607_),
    .X(_01739_));
 sky130_fd_sc_hd__or2_1 _08581_ (.A(_01449_),
    .B(_01739_),
    .X(_01740_));
 sky130_fd_sc_hd__nand2_1 _08582_ (.A(_01739_),
    .B(_01449_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand3_1 _08583_ (.A(_01740_),
    .B(_01610_),
    .C(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand2_1 _08584_ (.A(_01644_),
    .B(_01443_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_2 _08585_ (.A(_01742_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__inv_2 _08586_ (.A(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__nand2_1 _08587_ (.A(_01745_),
    .B(\sq.out[21] ),
    .Y(_01746_));
 sky130_fd_sc_hd__nand2_1 _08588_ (.A(_01744_),
    .B(_00455_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand2_1 _08589_ (.A(_01746_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _08590_ (.A(_01732_),
    .B(_01748_),
    .Y(_01750_));
 sky130_fd_sc_hd__nand2_1 _08591_ (.A(_01748_),
    .B(_01732_),
    .Y(_01751_));
 sky130_fd_sc_hd__and2b_1 _08592_ (.A_N(_01750_),
    .B(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__nand2_1 _08593_ (.A(_01737_),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__nand2_1 _08594_ (.A(_01741_),
    .B(_01447_),
    .Y(_01754_));
 sky130_fd_sc_hd__xor2_1 _08595_ (.A(_01467_),
    .B(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__nand2_1 _08596_ (.A(_01755_),
    .B(_01632_),
    .Y(_01756_));
 sky130_fd_sc_hd__or2_1 _08597_ (.A(_01460_),
    .B(_01610_),
    .X(_01757_));
 sky130_fd_sc_hd__nand2_2 _08598_ (.A(_01756_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__or2b_1 _08599_ (.A(_01758_),
    .B_N(_06106_),
    .X(_01759_));
 sky130_fd_sc_hd__buf_8 _08600_ (.A(_00177_),
    .X(\sq.out[22] ));
 sky130_fd_sc_hd__nand2_2 _08601_ (.A(_01758_),
    .B(\sq.out[22] ),
    .Y(_01761_));
 sky130_fd_sc_hd__nand2_1 _08602_ (.A(_01759_),
    .B(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2_1 _08603_ (.A(_01762_),
    .B(_01746_),
    .Y(_01763_));
 sky130_fd_sc_hd__nand3b_1 _08604_ (.A_N(_01746_),
    .B(_01759_),
    .C(_01761_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_1 _08605_ (.A(_01763_),
    .B(_01764_),
    .Y(_01765_));
 sky130_fd_sc_hd__inv_2 _08606_ (.A(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__nand2b_1 _08607_ (.A_N(_01469_),
    .B(_01739_),
    .Y(_01767_));
 sky130_fd_sc_hd__inv_2 _08608_ (.A(_01512_),
    .Y(_01768_));
 sky130_fd_sc_hd__nand2_1 _08609_ (.A(_01767_),
    .B(_01768_),
    .Y(_01769_));
 sky130_fd_sc_hd__nand2_1 _08610_ (.A(_01769_),
    .B(_01505_),
    .Y(_01771_));
 sky130_fd_sc_hd__nand3_1 _08611_ (.A(_01767_),
    .B(_01504_),
    .C(_01768_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand3_1 _08612_ (.A(_01771_),
    .B(_01632_),
    .C(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__or2_1 _08613_ (.A(_01492_),
    .B(_01610_),
    .X(_01774_));
 sky130_fd_sc_hd__nand2_2 _08614_ (.A(_01773_),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__inv_2 _08615_ (.A(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__clkbuf_8 _08616_ (.A(_00437_),
    .X(\sq.out[23] ));
 sky130_fd_sc_hd__nand2_1 _08617_ (.A(_01776_),
    .B(\sq.out[23] ),
    .Y(_01777_));
 sky130_fd_sc_hd__nand2_1 _08618_ (.A(_01775_),
    .B(_00743_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand2_1 _08619_ (.A(_01777_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__nor2_1 _08620_ (.A(_01761_),
    .B(_01779_),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _08621_ (.A(_01779_),
    .B(_01761_),
    .Y(_01782_));
 sky130_fd_sc_hd__and2b_1 _08622_ (.A_N(_01781_),
    .B(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__nand2_1 _08623_ (.A(_01766_),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _08624_ (.A(_01753_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__nand2_2 _08625_ (.A(_01722_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__xnor2_1 _08626_ (.A(_01761_),
    .B(_01779_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _08627_ (.A(_01765_),
    .B(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__o21ai_1 _08628_ (.A1(_01750_),
    .A2(_01734_),
    .B1(_01751_),
    .Y(_01789_));
 sky130_fd_sc_hd__o21ai_1 _08629_ (.A1(_01781_),
    .A2(_01763_),
    .B1(_01782_),
    .Y(_01790_));
 sky130_fd_sc_hd__a21oi_2 _08630_ (.A1(_01788_),
    .A2(_01789_),
    .B1(_01790_),
    .Y(_01792_));
 sky130_fd_sc_hd__nand2_4 _08631_ (.A(_01786_),
    .B(_01792_),
    .Y(_01793_));
 sky130_fd_sc_hd__a21o_1 _08632_ (.A1(_01607_),
    .A2(_01508_),
    .B1(_01516_),
    .X(_01794_));
 sky130_fd_sc_hd__xor2_1 _08633_ (.A(_01550_),
    .B(_01794_),
    .X(_01795_));
 sky130_fd_sc_hd__or2_1 _08634_ (.A(_01533_),
    .B(_01632_),
    .X(_01796_));
 sky130_fd_sc_hd__o21ai_2 _08635_ (.A1(_01644_),
    .A2(_01795_),
    .B1(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__a21bo_1 _08636_ (.A1(_01794_),
    .A2(_01549_),
    .B1_N(_01548_),
    .X(_01798_));
 sky130_fd_sc_hd__inv_2 _08637_ (.A(_01545_),
    .Y(_01799_));
 sky130_fd_sc_hd__and2_1 _08638_ (.A(_01798_),
    .B(_01799_),
    .X(_01800_));
 sky130_fd_sc_hd__o21ai_1 _08639_ (.A1(_01799_),
    .A2(_01798_),
    .B1(_01632_),
    .Y(_01801_));
 sky130_fd_sc_hd__o22ai_2 _08640_ (.A1(_01542_),
    .A2(_01632_),
    .B1(_01800_),
    .B2(_01801_),
    .Y(_01803_));
 sky130_fd_sc_hd__or2_1 _08641_ (.A(_01797_),
    .B(_01803_),
    .X(_01804_));
 sky130_fd_sc_hd__nand2_1 _08642_ (.A(_01803_),
    .B(_01797_),
    .Y(_01805_));
 sky130_fd_sc_hd__nand2_1 _08643_ (.A(_01804_),
    .B(_01805_),
    .Y(_01806_));
 sky130_fd_sc_hd__inv_2 _08644_ (.A(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__and2_1 _08645_ (.A(_01560_),
    .B(_01561_),
    .X(_01808_));
 sky130_fd_sc_hd__a21o_1 _08646_ (.A1(_01794_),
    .A2(_01552_),
    .B1(_01572_),
    .X(_01809_));
 sky130_fd_sc_hd__or2_1 _08647_ (.A(_01808_),
    .B(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__clkbuf_8 _08648_ (.A(_01632_),
    .X(\sq.out[10] ));
 sky130_fd_sc_hd__nand2_1 _08649_ (.A(_01809_),
    .B(_01808_),
    .Y(_01811_));
 sky130_fd_sc_hd__nand3_1 _08650_ (.A(_01810_),
    .B(\sq.out[10] ),
    .C(_01811_),
    .Y(_01813_));
 sky130_fd_sc_hd__nand2_1 _08651_ (.A(_01644_),
    .B(_01559_),
    .Y(_01814_));
 sky130_fd_sc_hd__nand2_2 _08652_ (.A(_01813_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__inv_2 _08653_ (.A(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand2_1 _08654_ (.A(_01807_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__nand2_1 _08655_ (.A(_01771_),
    .B(_01503_),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_1 _08656_ (.A(_01818_),
    .B(_01499_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand3_1 _08657_ (.A(_01771_),
    .B(_01498_),
    .C(_01503_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2_1 _08658_ (.A(_01819_),
    .B(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_01821_),
    .B(\sq.out[10] ),
    .Y(_01822_));
 sky130_fd_sc_hd__or2_1 _08660_ (.A(_01481_),
    .B(_01632_),
    .X(_01824_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(_01822_),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__a21o_1 _08662_ (.A1(_01825_),
    .A2(_01344_),
    .B1(_01797_),
    .X(_01826_));
 sky130_fd_sc_hd__nand3_1 _08663_ (.A(_01825_),
    .B(_01797_),
    .C(_01344_),
    .Y(_01827_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hd__nand2_1 _08665_ (.A(_01825_),
    .B(_01344_),
    .Y(_01829_));
 sky130_fd_sc_hd__nand3_1 _08666_ (.A(_01822_),
    .B(_01081_),
    .C(_01824_),
    .Y(_01830_));
 sky130_fd_sc_hd__nand2_1 _08667_ (.A(_01829_),
    .B(_01830_),
    .Y(_01831_));
 sky130_fd_sc_hd__nand2_1 _08668_ (.A(_01831_),
    .B(_01777_),
    .Y(_01832_));
 sky130_fd_sc_hd__or2_1 _08669_ (.A(_01777_),
    .B(_01831_),
    .X(_01833_));
 sky130_fd_sc_hd__nand3b_1 _08670_ (.A_N(_01828_),
    .B(_01832_),
    .C(_01833_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor2_2 _08671_ (.A(_01817_),
    .B(_01835_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_2 _08672_ (.A(_01793_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__inv_2 _08673_ (.A(_01827_),
    .Y(_01838_));
 sky130_fd_sc_hd__o21ai_1 _08674_ (.A1(_01838_),
    .A2(_01832_),
    .B1(_01826_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand3_1 _08675_ (.A(_01839_),
    .B(_01807_),
    .C(_01816_),
    .Y(_01840_));
 sky130_fd_sc_hd__and2_1 _08676_ (.A(_01805_),
    .B(_01816_),
    .X(_01841_));
 sky130_fd_sc_hd__nand2_1 _08677_ (.A(_01574_),
    .B(_01575_),
    .Y(_01842_));
 sky130_fd_sc_hd__a311o_4 _08678_ (.A1(_01794_),
    .A2(_01569_),
    .A3(_01552_),
    .B1(_01842_),
    .C1(_01644_),
    .X(_01843_));
 sky130_fd_sc_hd__or2_1 _08679_ (.A(_01524_),
    .B(_01843_),
    .X(_01844_));
 sky130_fd_sc_hd__buf_6 _08680_ (.A(_01844_),
    .X(_01846_));
 sky130_fd_sc_hd__nand3_1 _08681_ (.A(_01811_),
    .B(_01561_),
    .C(_01632_),
    .Y(_01847_));
 sky130_fd_sc_hd__xor2_2 _08682_ (.A(_01567_),
    .B(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__inv_2 _08683_ (.A(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_01843_),
    .B(_01524_),
    .Y(_01850_));
 sky130_fd_sc_hd__and3_1 _08685_ (.A(_01846_),
    .B(_01849_),
    .C(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__nand3_2 _08686_ (.A(_01840_),
    .B(_01841_),
    .C(_01851_),
    .Y(_01852_));
 sky130_fd_sc_hd__clkinvlp_2 _08687_ (.A(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand3_4 _08688_ (.A(_01837_),
    .B(_01853_),
    .C(_01846_),
    .Y(_01854_));
 sky130_fd_sc_hd__buf_8 _08689_ (.A(_01854_),
    .X(_01855_));
 sky130_fd_sc_hd__buf_6 _08690_ (.A(_01855_),
    .X(_01857_));
 sky130_fd_sc_hd__buf_6 _08691_ (.A(_01857_),
    .X(\sq.out[9] ));
 sky130_fd_sc_hd__a21oi_4 _08692_ (.A1(_01793_),
    .A2(_01836_),
    .B1(_01852_),
    .Y(_01858_));
 sky130_fd_sc_hd__nand2_1 _08693_ (.A(\sq.out[9] ),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__and2b_1 _08694_ (.A_N(_01859_),
    .B(_01846_),
    .X(_01860_));
 sky130_fd_sc_hd__buf_6 _08695_ (.A(_01860_),
    .X(_01861_));
 sky130_fd_sc_hd__nor2_2 _08696_ (.A(_01524_),
    .B(_01843_),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_2 _08697_ (.A(\sq.out[10] ),
    .B(_01855_),
    .Y(_01863_));
 sky130_fd_sc_hd__clkbuf_8 _08698_ (.A(_01368_),
    .X(\sq.out[11] ));
 sky130_fd_sc_hd__nand3_1 _08699_ (.A(_01863_),
    .B(_01363_),
    .C(\sq.out[11] ),
    .Y(_01864_));
 sky130_fd_sc_hd__inv_2 _08700_ (.A(_01864_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand2_2 _08701_ (.A(_01633_),
    .B(_01624_),
    .Y(_01867_));
 sky130_fd_sc_hd__a21oi_1 _08702_ (.A1(_01857_),
    .A2(_01531_),
    .B1(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__nand3_1 _08703_ (.A(_01858_),
    .B(_01644_),
    .C(_01846_),
    .Y(_01869_));
 sky130_fd_sc_hd__nand2_1 _08704_ (.A(_01855_),
    .B(_01867_),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _08705_ (.A(_01869_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__nand2_1 _08706_ (.A(_01871_),
    .B(\sq.out[12] ),
    .Y(_01872_));
 sky130_fd_sc_hd__nand3_1 _08707_ (.A(_01869_),
    .B(_01870_),
    .C(_01363_),
    .Y(_01873_));
 sky130_fd_sc_hd__nand2_1 _08708_ (.A(_01872_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2_1 _08709_ (.A(_01863_),
    .B(\sq.out[11] ),
    .Y(_01875_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_01874_),
    .B(_01875_),
    .Y(_01877_));
 sky130_fd_sc_hd__o21ai_2 _08711_ (.A1(_01866_),
    .A2(_01868_),
    .B1(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _08712_ (.A(_01863_),
    .B(_01531_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(_01855_),
    .B(_01621_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(_01879_),
    .B(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_2 _08715_ (.A(_01881_),
    .B(\sq.out[13] ),
    .Y(_01882_));
 sky130_fd_sc_hd__nand3_1 _08716_ (.A(_01879_),
    .B(_00843_),
    .C(_01880_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand2_1 _08717_ (.A(_01882_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(_01884_),
    .B(_01872_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand3b_1 _08719_ (.A_N(_01872_),
    .B(_01882_),
    .C(_01883_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand3_1 _08720_ (.A(_01878_),
    .B(_01885_),
    .C(_01886_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_1 _08721_ (.A(_01888_),
    .B(_01885_),
    .Y(_01889_));
 sky130_fd_sc_hd__clkinv_4 _08722_ (.A(_01854_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _08723_ (.A(_01890_),
    .B(_01630_),
    .Y(_01891_));
 sky130_fd_sc_hd__a21o_1 _08724_ (.A1(_01631_),
    .A2(_01625_),
    .B1(_01634_),
    .X(_01892_));
 sky130_fd_sc_hd__nand2_1 _08725_ (.A(_01892_),
    .B(_01635_),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _08726_ (.A(_01854_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand2_1 _08727_ (.A(_01891_),
    .B(_01894_),
    .Y(_01895_));
 sky130_fd_sc_hd__or2_4 _08728_ (.A(_01587_),
    .B(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__inv_2 _08729_ (.A(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__a21o_1 _08730_ (.A1(_01626_),
    .A2(_01629_),
    .B1(_01635_),
    .X(_01899_));
 sky130_fd_sc_hd__nand3_1 _08731_ (.A(_01854_),
    .B(_01636_),
    .C(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__nand2_1 _08732_ (.A(_01890_),
    .B(_01614_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _08733_ (.A(_01900_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__or2_4 _08734_ (.A(_01286_),
    .B(_01902_),
    .X(_01903_));
 sky130_fd_sc_hd__nand2_1 _08735_ (.A(_01902_),
    .B(_01286_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand3_1 _08736_ (.A(_01897_),
    .B(_01903_),
    .C(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_1 _08737_ (.A(_01903_),
    .B(_01904_),
    .Y(_01906_));
 sky130_fd_sc_hd__nand2_1 _08738_ (.A(_01906_),
    .B(_01896_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_2 _08739_ (.A(_01905_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__inv_2 _08740_ (.A(_01908_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand2_1 _08741_ (.A(_01895_),
    .B(_01587_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_2 _08742_ (.A(_01896_),
    .B(_01911_),
    .Y(_01912_));
 sky130_fd_sc_hd__xor2_2 _08743_ (.A(_01882_),
    .B(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__nand3_1 _08744_ (.A(_01889_),
    .B(_01910_),
    .C(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__and2_1 _08745_ (.A(_01906_),
    .B(_01896_),
    .X(_01915_));
 sky130_fd_sc_hd__nand2_1 _08746_ (.A(_01912_),
    .B(_01882_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _08747_ (.A(_01916_),
    .B(_01908_),
    .Y(_01917_));
 sky130_fd_sc_hd__nor2_1 _08748_ (.A(_01915_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__nand2_1 _08749_ (.A(_01914_),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__or2_1 _08750_ (.A(_01655_),
    .B(_01637_),
    .X(_01921_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(_01921_),
    .B(_01656_),
    .Y(_01922_));
 sky130_fd_sc_hd__nand2_1 _08752_ (.A(_01890_),
    .B(_01647_),
    .Y(_01923_));
 sky130_fd_sc_hd__o21ai_2 _08753_ (.A1(_01922_),
    .A2(_01890_),
    .B1(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__or2_1 _08754_ (.A(_00091_),
    .B(_01924_),
    .X(_01925_));
 sky130_fd_sc_hd__nand2_1 _08755_ (.A(_01657_),
    .B(_01685_),
    .Y(_01926_));
 sky130_fd_sc_hd__or2_1 _08756_ (.A(_01685_),
    .B(_01657_),
    .X(_01927_));
 sky130_fd_sc_hd__nand3_1 _08757_ (.A(_01855_),
    .B(_01926_),
    .C(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__o21ai_2 _08758_ (.A1(_01663_),
    .A2(_01855_),
    .B1(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__or2_1 _08759_ (.A(_01240_),
    .B(_01929_),
    .X(_01930_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_01929_),
    .B(_01240_),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_1 _08761_ (.A(_01930_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__or2_1 _08762_ (.A(_01925_),
    .B(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__nand2_1 _08763_ (.A(_01933_),
    .B(_01925_),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_1 _08764_ (.A(_01934_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__inv_2 _08765_ (.A(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(_01924_),
    .B(_00091_),
    .Y(_01938_));
 sky130_fd_sc_hd__nand2_1 _08767_ (.A(_01925_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__or2_1 _08768_ (.A(_01903_),
    .B(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__nand2_1 _08769_ (.A(_01939_),
    .B(_01903_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand2_1 _08770_ (.A(_01940_),
    .B(_01941_),
    .Y(_01943_));
 sky130_fd_sc_hd__inv_2 _08771_ (.A(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__nand3_1 _08772_ (.A(_01919_),
    .B(_01937_),
    .C(_01944_),
    .Y(_01945_));
 sky130_fd_sc_hd__o21a_1 _08773_ (.A1(_01941_),
    .A2(_01936_),
    .B1(_01935_),
    .X(_01946_));
 sky130_fd_sc_hd__nand2_1 _08774_ (.A(_01945_),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__a21o_1 _08775_ (.A1(_01686_),
    .A2(_01687_),
    .B1(_01718_),
    .X(_01948_));
 sky130_fd_sc_hd__or2b_1 _08776_ (.A(_01688_),
    .B_N(_01718_),
    .X(_01949_));
 sky130_fd_sc_hd__nand3_1 _08777_ (.A(_01857_),
    .B(_01948_),
    .C(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(_01890_),
    .B(_01711_),
    .Y(_01951_));
 sky130_fd_sc_hd__nand2_1 _08779_ (.A(_01950_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__inv_2 _08780_ (.A(_01952_),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_1 _08781_ (.A(_01954_),
    .B(\sq.out[19] ),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _08782_ (.A(_01952_),
    .B(_05130_),
    .Y(_01956_));
 sky130_fd_sc_hd__nand2_1 _08783_ (.A(_01955_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _08784_ (.A(_01926_),
    .B(_01682_),
    .Y(_01958_));
 sky130_fd_sc_hd__or2_1 _08785_ (.A(_01678_),
    .B(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__nand2_1 _08786_ (.A(_01958_),
    .B(_01678_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2_1 _08787_ (.A(_01670_),
    .B(_01855_),
    .Y(_01961_));
 sky130_fd_sc_hd__a31o_1 _08788_ (.A1(_01857_),
    .A2(_01959_),
    .A3(_01960_),
    .B1(_01961_),
    .X(_01962_));
 sky130_fd_sc_hd__or2_1 _08789_ (.A(_01712_),
    .B(_01962_),
    .X(_01963_));
 sky130_fd_sc_hd__or2_1 _08790_ (.A(_01957_),
    .B(_01963_),
    .X(_01965_));
 sky130_fd_sc_hd__nand2_1 _08791_ (.A(_01963_),
    .B(_01957_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _08792_ (.A(_01965_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__nand2_1 _08793_ (.A(_01962_),
    .B(_01712_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _08794_ (.A(_01963_),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__or2_1 _08795_ (.A(_01930_),
    .B(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__nand2_1 _08796_ (.A(_01969_),
    .B(_01930_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_01970_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__nor2_1 _08798_ (.A(_01967_),
    .B(_01972_),
    .Y(_01973_));
 sky130_fd_sc_hd__nand2_1 _08799_ (.A(_01947_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__o21a_1 _08800_ (.A1(_01971_),
    .A2(_01967_),
    .B1(_01966_),
    .X(_01976_));
 sky130_fd_sc_hd__nand2_2 _08801_ (.A(_01974_),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__nand2_1 _08802_ (.A(_01722_),
    .B(_01737_),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _08803_ (.A(_01978_),
    .B(_01734_),
    .Y(_01979_));
 sky130_fd_sc_hd__or2_1 _08804_ (.A(_01752_),
    .B(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_01979_),
    .B(_01752_),
    .Y(_01981_));
 sky130_fd_sc_hd__a21o_1 _08806_ (.A1(_01980_),
    .A2(_01981_),
    .B1(_01890_),
    .X(_01982_));
 sky130_fd_sc_hd__nand2_1 _08807_ (.A(_01890_),
    .B(_01745_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _08808_ (.A(_01982_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand2_1 _08809_ (.A(_01984_),
    .B(\sq.out[22] ),
    .Y(_01985_));
 sky130_fd_sc_hd__a31o_1 _08810_ (.A1(_01722_),
    .A2(_01752_),
    .A3(_01737_),
    .B1(_01789_),
    .X(_01987_));
 sky130_fd_sc_hd__or2_1 _08811_ (.A(_01766_),
    .B(_01987_),
    .X(_01988_));
 sky130_fd_sc_hd__nand2_1 _08812_ (.A(_01987_),
    .B(_01766_),
    .Y(_01989_));
 sky130_fd_sc_hd__nand3_1 _08813_ (.A(_01988_),
    .B(_01855_),
    .C(_01989_),
    .Y(_01990_));
 sky130_fd_sc_hd__o21ai_2 _08814_ (.A1(_01758_),
    .A2(_01855_),
    .B1(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__or2_1 _08815_ (.A(_00743_),
    .B(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__buf_6 _08816_ (.A(_00743_),
    .X(_01993_));
 sky130_fd_sc_hd__nand2_1 _08817_ (.A(_01991_),
    .B(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__nand2_1 _08818_ (.A(_01992_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__or2_1 _08819_ (.A(_01985_),
    .B(_01995_),
    .X(_01996_));
 sky130_fd_sc_hd__nand2_1 _08820_ (.A(_01995_),
    .B(_01985_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_1 _08821_ (.A(_01996_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__clkinvlp_2 _08822_ (.A(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__or2_1 _08823_ (.A(_01737_),
    .B(_01722_),
    .X(_02001_));
 sky130_fd_sc_hd__nand3_1 _08824_ (.A(_01855_),
    .B(_01978_),
    .C(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hd__nand2_1 _08825_ (.A(_01890_),
    .B(_01729_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _08826_ (.A(_02002_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__inv_2 _08827_ (.A(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_1 _08828_ (.A(_02005_),
    .B(\sq.out[21] ),
    .Y(_02006_));
 sky130_fd_sc_hd__inv_2 _08829_ (.A(_01984_),
    .Y(_02007_));
 sky130_fd_sc_hd__buf_6 _08830_ (.A(_06106_),
    .X(_02009_));
 sky130_fd_sc_hd__nand2_1 _08831_ (.A(_02007_),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _08832_ (.A(_02010_),
    .B(_01985_),
    .Y(_02011_));
 sky130_fd_sc_hd__or2_1 _08833_ (.A(_02006_),
    .B(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__nand2_1 _08834_ (.A(_02011_),
    .B(_02006_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(_02012_),
    .B(_02013_),
    .Y(_02014_));
 sky130_fd_sc_hd__clkinvlp_2 _08836_ (.A(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__buf_6 _08837_ (.A(_01890_),
    .X(_02016_));
 sky130_fd_sc_hd__nand2_1 _08838_ (.A(_02016_),
    .B(_01703_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand2_1 _08839_ (.A(_01948_),
    .B(_01717_),
    .Y(_02018_));
 sky130_fd_sc_hd__xor2_1 _08840_ (.A(_01710_),
    .B(_02018_),
    .X(_02020_));
 sky130_fd_sc_hd__nand2_1 _08841_ (.A(_01857_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(_02017_),
    .B(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__inv_2 _08843_ (.A(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__nand2_1 _08844_ (.A(_02023_),
    .B(_01730_),
    .Y(_02024_));
 sky130_fd_sc_hd__clkbuf_8 _08845_ (.A(_00460_),
    .X(\sq.out[20] ));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(_02022_),
    .B(\sq.out[20] ),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _08847_ (.A(_02024_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__or2_1 _08848_ (.A(_01955_),
    .B(_02026_),
    .X(_02027_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(_02026_),
    .B(_01955_),
    .Y(_02028_));
 sky130_fd_sc_hd__nand2_1 _08850_ (.A(_02027_),
    .B(_02028_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _08851_ (.A(_02004_),
    .B(_00455_),
    .Y(_02031_));
 sky130_fd_sc_hd__nand2_1 _08852_ (.A(_02006_),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__or2_1 _08853_ (.A(_02025_),
    .B(_02032_),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_02032_),
    .B(_02025_),
    .Y(_02034_));
 sky130_fd_sc_hd__nand2_1 _08855_ (.A(_02033_),
    .B(_02034_),
    .Y(_02035_));
 sky130_fd_sc_hd__nor2_1 _08856_ (.A(_02030_),
    .B(_02035_),
    .Y(_02036_));
 sky130_fd_sc_hd__and3_1 _08857_ (.A(_02000_),
    .B(_02015_),
    .C(_02036_),
    .X(_02037_));
 sky130_fd_sc_hd__nand2_2 _08858_ (.A(_01977_),
    .B(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__o21a_1 _08859_ (.A1(_02028_),
    .A2(_02035_),
    .B1(_02034_),
    .X(_02039_));
 sky130_fd_sc_hd__o21a_1 _08860_ (.A1(_02013_),
    .A2(_01999_),
    .B1(_01998_),
    .X(_02041_));
 sky130_fd_sc_hd__o31a_1 _08861_ (.A1(_01999_),
    .A2(_02014_),
    .A3(_02039_),
    .B1(_02041_),
    .X(_02042_));
 sky130_fd_sc_hd__nand2_4 _08862_ (.A(_02038_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21oi_1 _08863_ (.A1(_01786_),
    .A2(_01792_),
    .B1(_01835_),
    .Y(_02044_));
 sky130_fd_sc_hd__or2_1 _08864_ (.A(_01839_),
    .B(_02044_),
    .X(_02045_));
 sky130_fd_sc_hd__or2_1 _08865_ (.A(_01807_),
    .B(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_02045_),
    .B(_01807_),
    .Y(_02047_));
 sky130_fd_sc_hd__nand3_1 _08867_ (.A(_02046_),
    .B(_01857_),
    .C(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(_02016_),
    .B(_01803_),
    .Y(_02049_));
 sky130_fd_sc_hd__nand2_4 _08869_ (.A(_02048_),
    .B(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_01833_),
    .B(_01832_),
    .Y(_02052_));
 sky130_fd_sc_hd__xor2_2 _08871_ (.A(_02052_),
    .B(_01793_),
    .X(_02053_));
 sky130_fd_sc_hd__or2_1 _08872_ (.A(_01825_),
    .B(_01857_),
    .X(_02054_));
 sky130_fd_sc_hd__o21ai_4 _08873_ (.A1(_02016_),
    .A2(_02053_),
    .B1(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__a21bo_1 _08874_ (.A1(_01793_),
    .A2(_01833_),
    .B1_N(_01832_),
    .X(_02056_));
 sky130_fd_sc_hd__xor2_1 _08875_ (.A(_01828_),
    .B(_02056_),
    .X(_02057_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(_02016_),
    .B(_01797_),
    .Y(_02058_));
 sky130_fd_sc_hd__o21ai_2 _08877_ (.A1(_02016_),
    .A2(_02057_),
    .B1(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__or2_1 _08878_ (.A(_02055_),
    .B(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__nand2_1 _08879_ (.A(_02059_),
    .B(_02055_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _08880_ (.A(_02060_),
    .B(_02061_),
    .Y(_02063_));
 sky130_fd_sc_hd__or2_1 _08881_ (.A(_02050_),
    .B(_02063_),
    .X(_02064_));
 sky130_fd_sc_hd__nand2_1 _08882_ (.A(_01989_),
    .B(_01763_),
    .Y(_02065_));
 sky130_fd_sc_hd__xor2_1 _08883_ (.A(_01787_),
    .B(_02065_),
    .X(_02066_));
 sky130_fd_sc_hd__nand2_1 _08884_ (.A(_02066_),
    .B(_01857_),
    .Y(_02067_));
 sky130_fd_sc_hd__o21ai_4 _08885_ (.A1(_01775_),
    .A2(_01857_),
    .B1(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(_02068_),
    .B(_01344_),
    .Y(_02069_));
 sky130_fd_sc_hd__nand2b_1 _08887_ (.A_N(_02069_),
    .B(_02055_),
    .Y(_02070_));
 sky130_fd_sc_hd__buf_6 _08888_ (.A(_01344_),
    .X(_02071_));
 sky130_fd_sc_hd__a21o_1 _08889_ (.A1(_02068_),
    .A2(_02071_),
    .B1(_02055_),
    .X(_02072_));
 sky130_fd_sc_hd__nand2_1 _08890_ (.A(_02070_),
    .B(_02072_),
    .Y(_02074_));
 sky130_fd_sc_hd__or2_1 _08891_ (.A(_01344_),
    .B(_02068_),
    .X(_02075_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(_02075_),
    .B(_02069_),
    .Y(_02076_));
 sky130_fd_sc_hd__or2_1 _08893_ (.A(_01992_),
    .B(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__nand2_1 _08894_ (.A(_02076_),
    .B(_01992_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand2_1 _08895_ (.A(_02077_),
    .B(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__nor2_1 _08896_ (.A(_02074_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__and2b_1 _08897_ (.A_N(_02064_),
    .B(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__nand2_2 _08898_ (.A(_02043_),
    .B(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__or2_1 _08899_ (.A(_01524_),
    .B(_01843_),
    .X(_02083_));
 sky130_fd_sc_hd__buf_6 _08900_ (.A(_02083_),
    .X(_02085_));
 sky130_fd_sc_hd__o21a_1 _08901_ (.A1(_02074_),
    .A2(_02078_),
    .B1(_02072_),
    .X(_02086_));
 sky130_fd_sc_hd__inv_2 _08902_ (.A(_02050_),
    .Y(_02087_));
 sky130_fd_sc_hd__and2_1 _08903_ (.A(_02061_),
    .B(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__o21a_1 _08904_ (.A1(_02064_),
    .A2(_02086_),
    .B1(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__clkinvlp_2 _08905_ (.A(_01837_),
    .Y(_02090_));
 sky130_fd_sc_hd__and2_1 _08906_ (.A(_01840_),
    .B(_01841_),
    .X(_02091_));
 sky130_fd_sc_hd__or3b_1 _08907_ (.A(_02090_),
    .B(_02016_),
    .C_N(_02091_),
    .X(_02092_));
 sky130_fd_sc_hd__or2_1 _08908_ (.A(_01848_),
    .B(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__nand2_1 _08909_ (.A(_02092_),
    .B(_01848_),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_2 _08910_ (.A(_02093_),
    .B(_02094_),
    .Y(_02096_));
 sky130_fd_sc_hd__or2_1 _08911_ (.A(_01524_),
    .B(_01843_),
    .X(_02097_));
 sky130_fd_sc_hd__a32oi_1 _08912_ (.A1(_01837_),
    .A2(_02091_),
    .A3(_01849_),
    .B1(_01846_),
    .B2(_01850_),
    .Y(_02098_));
 sky130_fd_sc_hd__inv_1 _08913_ (.A(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand3_1 _08914_ (.A(_02047_),
    .B(_01805_),
    .C(_01857_),
    .Y(_02100_));
 sky130_fd_sc_hd__xor2_2 _08915_ (.A(_01815_),
    .B(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__and4b_1 _08916_ (.A_N(_02096_),
    .B(_02097_),
    .C(_02099_),
    .D(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__nand2_1 _08917_ (.A(_02089_),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__inv_2 _08918_ (.A(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__nand3_4 _08919_ (.A(_02082_),
    .B(_02085_),
    .C(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__buf_6 _08920_ (.A(_02105_),
    .X(_02107_));
 sky130_fd_sc_hd__buf_8 _08921_ (.A(_02107_),
    .X(_02108_));
 sky130_fd_sc_hd__a21oi_4 _08922_ (.A1(_02043_),
    .A2(_02081_),
    .B1(_02103_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_4 _08923_ (.A(_02108_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__or2_4 _08924_ (.A(_01862_),
    .B(_02110_),
    .X(_02111_));
 sky130_fd_sc_hd__inv_2 _08925_ (.A(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__nor2_1 _08926_ (.A(_01861_),
    .B(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__or2b_1 _08927_ (.A(_01859_),
    .B_N(_01846_),
    .X(_02114_));
 sky130_fd_sc_hd__inv_2 _08928_ (.A(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__or2_1 _08929_ (.A(_01524_),
    .B(_01843_),
    .X(_02116_));
 sky130_fd_sc_hd__a211o_1 _08930_ (.A1(_02109_),
    .A2(_02116_),
    .B1(_01846_),
    .C1(_01858_),
    .X(_02118_));
 sky130_fd_sc_hd__inv_2 _08931_ (.A(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand3_1 _08932_ (.A(_02105_),
    .B(_02082_),
    .C(_02089_),
    .Y(_02120_));
 sky130_fd_sc_hd__inv_2 _08933_ (.A(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_1 _08934_ (.A(_02121_),
    .B(_02101_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _08935_ (.A(_02096_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _08936_ (.A(_02123_),
    .B(_02099_),
    .Y(_02124_));
 sky130_fd_sc_hd__xor2_1 _08937_ (.A(_02097_),
    .B(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__nand3_1 _08938_ (.A(_02109_),
    .B(_02085_),
    .C(_01902_),
    .Y(_02126_));
 sky130_fd_sc_hd__a21bo_1 _08939_ (.A1(_01889_),
    .A2(_01913_),
    .B1_N(_01916_),
    .X(_02127_));
 sky130_fd_sc_hd__xor2_1 _08940_ (.A(_01908_),
    .B(_02127_),
    .X(_02129_));
 sky130_fd_sc_hd__clkinvlp_2 _08941_ (.A(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_1 _08942_ (.A(_02108_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(_02126_),
    .B(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__nand2_1 _08944_ (.A(_02132_),
    .B(_00091_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand3_1 _08945_ (.A(_02126_),
    .B(\sq.out[16] ),
    .C(_02131_),
    .Y(_02134_));
 sky130_fd_sc_hd__nand2_1 _08946_ (.A(_02133_),
    .B(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__inv_6 _08947_ (.A(_02105_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_1 _08948_ (.A(_02136_),
    .B(_01895_),
    .Y(_02137_));
 sky130_fd_sc_hd__xor2_1 _08949_ (.A(_01913_),
    .B(_01889_),
    .X(_02138_));
 sky130_fd_sc_hd__nand2_1 _08950_ (.A(_02107_),
    .B(_02138_),
    .Y(_02140_));
 sky130_fd_sc_hd__nand3_1 _08951_ (.A(_02137_),
    .B(\sq.out[15] ),
    .C(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(_02135_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__nand3_1 _08953_ (.A(_02109_),
    .B(_02085_),
    .C(_01924_),
    .Y(_02143_));
 sky130_fd_sc_hd__xor2_1 _08954_ (.A(_01943_),
    .B(_01919_),
    .X(_02144_));
 sky130_fd_sc_hd__inv_2 _08955_ (.A(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand2_1 _08956_ (.A(_02107_),
    .B(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(_02143_),
    .B(_02146_),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_1 _08958_ (.A(_02147_),
    .B(_01240_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand3_2 _08959_ (.A(_02143_),
    .B(\sq.out[17] ),
    .C(_02146_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand2_1 _08960_ (.A(_02148_),
    .B(_02149_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_1 _08961_ (.A(_02134_),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_1 _08962_ (.A(_02151_),
    .B(_02134_),
    .Y(_02153_));
 sky130_fd_sc_hd__o21ai_1 _08963_ (.A1(_02142_),
    .A2(_02152_),
    .B1(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__nand3_1 _08964_ (.A(_02109_),
    .B(_02085_),
    .C(_01962_),
    .Y(_02155_));
 sky130_fd_sc_hd__xor2_1 _08965_ (.A(_01972_),
    .B(_01947_),
    .X(_02156_));
 sky130_fd_sc_hd__inv_2 _08966_ (.A(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__nand2_1 _08967_ (.A(_02108_),
    .B(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__nand2_1 _08968_ (.A(_02155_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_02159_),
    .B(_05130_),
    .Y(_02160_));
 sky130_fd_sc_hd__nand3_1 _08970_ (.A(_02155_),
    .B(\sq.out[19] ),
    .C(_02158_),
    .Y(_02162_));
 sky130_fd_sc_hd__nand2_1 _08971_ (.A(_02160_),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__nand3_1 _08972_ (.A(_02109_),
    .B(_02085_),
    .C(_01929_),
    .Y(_02164_));
 sky130_fd_sc_hd__buf_6 _08973_ (.A(_06002_),
    .X(\sq.out[18] ));
 sky130_fd_sc_hd__a21bo_1 _08974_ (.A1(_01919_),
    .A2(_01944_),
    .B1_N(_01941_),
    .X(_02165_));
 sky130_fd_sc_hd__xor2_1 _08975_ (.A(_01937_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__nand2_1 _08976_ (.A(net105),
    .B(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__nand3_2 _08977_ (.A(_02164_),
    .B(\sq.out[18] ),
    .C(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _08978_ (.A(_02163_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__inv_2 _08979_ (.A(_02168_),
    .Y(_02170_));
 sky130_fd_sc_hd__nand3_1 _08980_ (.A(_02170_),
    .B(_02160_),
    .C(_02162_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _08981_ (.A(_02169_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_1 _08982_ (.A(_02164_),
    .B(_02167_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand2_1 _08983_ (.A(_02174_),
    .B(_01712_),
    .Y(_02175_));
 sky130_fd_sc_hd__nand2_1 _08984_ (.A(_02175_),
    .B(_02168_),
    .Y(_02176_));
 sky130_fd_sc_hd__nand2_1 _08985_ (.A(_02176_),
    .B(_02149_),
    .Y(_02177_));
 sky130_fd_sc_hd__inv_2 _08986_ (.A(_02149_),
    .Y(_02178_));
 sky130_fd_sc_hd__nand3_1 _08987_ (.A(_02178_),
    .B(_02175_),
    .C(_02168_),
    .Y(_02179_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(_02177_),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _08989_ (.A(_02173_),
    .B(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _08990_ (.A(_02154_),
    .B(_02181_),
    .Y(_02183_));
 sky130_fd_sc_hd__and2_1 _08991_ (.A(_02176_),
    .B(_02149_),
    .X(_02184_));
 sky130_fd_sc_hd__a21boi_1 _08992_ (.A1(_02184_),
    .A2(_02172_),
    .B1_N(_02169_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand2_1 _08993_ (.A(_02183_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _08994_ (.A(_02136_),
    .B(_02005_),
    .Y(_02187_));
 sky130_fd_sc_hd__inv_2 _08995_ (.A(_02030_),
    .Y(_02188_));
 sky130_fd_sc_hd__nand2_1 _08996_ (.A(_01977_),
    .B(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__nand2_1 _08997_ (.A(_02189_),
    .B(_02028_),
    .Y(_02190_));
 sky130_fd_sc_hd__xor2_1 _08998_ (.A(_02035_),
    .B(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__nand2_1 _08999_ (.A(_02191_),
    .B(_02105_),
    .Y(_02192_));
 sky130_fd_sc_hd__nand2_1 _09000_ (.A(_02187_),
    .B(_02192_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_1 _09001_ (.A(_02194_),
    .B(\sq.out[22] ),
    .Y(_02195_));
 sky130_fd_sc_hd__inv_2 _09002_ (.A(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _09003_ (.A(_01977_),
    .B(_02036_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _09004_ (.A(_02197_),
    .B(_02039_),
    .Y(_02198_));
 sky130_fd_sc_hd__nand2_1 _09005_ (.A(_02198_),
    .B(_02015_),
    .Y(_02199_));
 sky130_fd_sc_hd__or2_1 _09006_ (.A(_02015_),
    .B(_02198_),
    .X(_02200_));
 sky130_fd_sc_hd__nand3_2 _09007_ (.A(net105),
    .B(_02199_),
    .C(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__nand2_1 _09008_ (.A(_02136_),
    .B(_02007_),
    .Y(_02202_));
 sky130_fd_sc_hd__nand3_2 _09009_ (.A(_02201_),
    .B(_02202_),
    .C(\sq.out[23] ),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2_1 _09010_ (.A(_02201_),
    .B(_02202_),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(_02205_),
    .B(_01993_),
    .Y(_02206_));
 sky130_fd_sc_hd__nand3_1 _09012_ (.A(_02196_),
    .B(_02203_),
    .C(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__nand2_1 _09013_ (.A(_02206_),
    .B(_02203_),
    .Y(_02208_));
 sky130_fd_sc_hd__nand2_1 _09014_ (.A(_02208_),
    .B(_02195_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_02207_),
    .B(_02209_),
    .Y(_02210_));
 sky130_fd_sc_hd__inv_2 _09016_ (.A(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__nand3_1 _09017_ (.A(_02187_),
    .B(_02192_),
    .C(_02009_),
    .Y(_02212_));
 sky130_fd_sc_hd__nand2_1 _09018_ (.A(_02195_),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__nand2_1 _09019_ (.A(_02136_),
    .B(_02023_),
    .Y(_02214_));
 sky130_fd_sc_hd__or2_1 _09020_ (.A(_02188_),
    .B(_01977_),
    .X(_02216_));
 sky130_fd_sc_hd__nand2_1 _09021_ (.A(_02216_),
    .B(_02189_),
    .Y(_02217_));
 sky130_fd_sc_hd__inv_2 _09022_ (.A(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nand2_1 _09023_ (.A(net105),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__nand3_2 _09024_ (.A(_02214_),
    .B(\sq.out[21] ),
    .C(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand2_1 _09025_ (.A(_02213_),
    .B(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__inv_2 _09026_ (.A(_02220_),
    .Y(_02222_));
 sky130_fd_sc_hd__nand3_1 _09027_ (.A(_02222_),
    .B(_02195_),
    .C(_02212_),
    .Y(_02223_));
 sky130_fd_sc_hd__nand2_1 _09028_ (.A(_02221_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__inv_2 _09029_ (.A(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__nand2_1 _09030_ (.A(_02211_),
    .B(_02225_),
    .Y(_02227_));
 sky130_fd_sc_hd__nand2_1 _09031_ (.A(_02136_),
    .B(_01954_),
    .Y(_02228_));
 sky130_fd_sc_hd__a21bo_1 _09032_ (.A1(_01947_),
    .A2(_01970_),
    .B1_N(_01971_),
    .X(_02229_));
 sky130_fd_sc_hd__xor2_1 _09033_ (.A(_01967_),
    .B(_02229_),
    .X(_02230_));
 sky130_fd_sc_hd__nand2_1 _09034_ (.A(_02107_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__nand2_1 _09035_ (.A(_02228_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__nand2_2 _09036_ (.A(_02232_),
    .B(\sq.out[20] ),
    .Y(_02233_));
 sky130_fd_sc_hd__inv_2 _09037_ (.A(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2_1 _09038_ (.A(_02214_),
    .B(_02219_),
    .Y(_02235_));
 sky130_fd_sc_hd__nand2_1 _09039_ (.A(_02235_),
    .B(_00455_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand3_1 _09040_ (.A(_02234_),
    .B(_02220_),
    .C(_02236_),
    .Y(_02238_));
 sky130_fd_sc_hd__nand2_1 _09041_ (.A(_02236_),
    .B(_02220_),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_1 _09042_ (.A(_02239_),
    .B(_02233_),
    .Y(_02240_));
 sky130_fd_sc_hd__nand2_1 _09043_ (.A(_02238_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__inv_2 _09044_ (.A(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand3_1 _09045_ (.A(_02228_),
    .B(_01730_),
    .C(_02231_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand3b_1 _09046_ (.A_N(_02162_),
    .B(_02233_),
    .C(_02243_),
    .Y(_02244_));
 sky130_fd_sc_hd__nand2_1 _09047_ (.A(_02233_),
    .B(_02243_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand2_1 _09048_ (.A(_02245_),
    .B(_02162_),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_1 _09049_ (.A(_02244_),
    .B(_02246_),
    .Y(_02247_));
 sky130_fd_sc_hd__inv_2 _09050_ (.A(_02247_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_1 _09051_ (.A(_02242_),
    .B(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _09052_ (.A(_02227_),
    .B(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__nand2_1 _09053_ (.A(_02186_),
    .B(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor2_1 _09054_ (.A(_02233_),
    .B(_02239_),
    .Y(_02253_));
 sky130_fd_sc_hd__o21ai_1 _09055_ (.A1(_02246_),
    .A2(_02253_),
    .B1(_02240_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor2_1 _09056_ (.A(_02224_),
    .B(_02210_),
    .Y(_02255_));
 sky130_fd_sc_hd__inv_2 _09057_ (.A(_02207_),
    .Y(_02256_));
 sky130_fd_sc_hd__o21ai_1 _09058_ (.A1(_02221_),
    .A2(_02256_),
    .B1(_02209_),
    .Y(_02257_));
 sky130_fd_sc_hd__a21oi_1 _09059_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__nand2_1 _09060_ (.A(_02252_),
    .B(_02258_),
    .Y(_02260_));
 sky130_fd_sc_hd__nand2_1 _09061_ (.A(_02043_),
    .B(_02080_),
    .Y(_02261_));
 sky130_fd_sc_hd__a21o_1 _09062_ (.A1(_02261_),
    .A2(_02086_),
    .B1(_02063_),
    .X(_02262_));
 sky130_fd_sc_hd__and3_1 _09063_ (.A(_02262_),
    .B(_02061_),
    .C(_02108_),
    .X(_02263_));
 sky130_fd_sc_hd__xor2_2 _09064_ (.A(_02050_),
    .B(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__nand2_1 _09065_ (.A(_02122_),
    .B(_02096_),
    .Y(_02265_));
 sky130_fd_sc_hd__and2b_1 _09066_ (.A_N(_02123_),
    .B(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__or2_1 _09067_ (.A(_02101_),
    .B(_02121_),
    .X(_02267_));
 sky130_fd_sc_hd__nand2_1 _09068_ (.A(_02267_),
    .B(_02122_),
    .Y(_02268_));
 sky130_fd_sc_hd__inv_2 _09069_ (.A(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _09070_ (.A(_02266_),
    .B(_02269_),
    .Y(_02271_));
 sky130_fd_sc_hd__nor2_1 _09071_ (.A(_02264_),
    .B(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__or2_1 _09072_ (.A(_02099_),
    .B(_02123_),
    .X(_02273_));
 sky130_fd_sc_hd__nand2_1 _09073_ (.A(_02273_),
    .B(_02124_),
    .Y(_02274_));
 sky130_fd_sc_hd__inv_2 _09074_ (.A(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_1 _09075_ (.A(_02272_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__xor2_1 _09076_ (.A(_02079_),
    .B(_02043_),
    .X(_02277_));
 sky130_fd_sc_hd__nand2b_1 _09077_ (.A_N(_02277_),
    .B(net105),
    .Y(_02278_));
 sky130_fd_sc_hd__o21ai_4 _09078_ (.A1(_02068_),
    .A2(_02108_),
    .B1(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__nand2_1 _09079_ (.A(_02199_),
    .B(_02013_),
    .Y(_02280_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(_02280_),
    .B(_02000_),
    .Y(_02282_));
 sky130_fd_sc_hd__nand3_1 _09081_ (.A(_02199_),
    .B(_01999_),
    .C(_02013_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _09082_ (.A(_02282_),
    .B(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hd__buf_8 _09083_ (.A(_02108_),
    .X(\sq.out[8] ));
 sky130_fd_sc_hd__nand2_1 _09084_ (.A(_02284_),
    .B(\sq.out[8] ),
    .Y(_02285_));
 sky130_fd_sc_hd__or2_1 _09085_ (.A(_01991_),
    .B(_02108_),
    .X(_02286_));
 sky130_fd_sc_hd__nand2_1 _09086_ (.A(_02285_),
    .B(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand3_1 _09087_ (.A(_02279_),
    .B(_02071_),
    .C(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__inv_2 _09088_ (.A(_02279_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _09089_ (.A(_02287_),
    .B(_02071_),
    .Y(_02290_));
 sky130_fd_sc_hd__nand2_1 _09090_ (.A(_02289_),
    .B(_02290_),
    .Y(_02292_));
 sky130_fd_sc_hd__nand2_1 _09091_ (.A(_02288_),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__nand3_1 _09092_ (.A(_02285_),
    .B(_02286_),
    .C(_01081_),
    .Y(_02294_));
 sky130_fd_sc_hd__inv_2 _09093_ (.A(_02203_),
    .Y(_02295_));
 sky130_fd_sc_hd__a21o_1 _09094_ (.A1(_02290_),
    .A2(_02294_),
    .B1(_02295_),
    .X(_02296_));
 sky130_fd_sc_hd__nand3_1 _09095_ (.A(_02290_),
    .B(_02295_),
    .C(_02294_),
    .Y(_02297_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_02296_),
    .B(_02297_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_2 _09097_ (.A(_02298_),
    .B(_02293_),
    .Y(_02299_));
 sky130_fd_sc_hd__inv_2 _09098_ (.A(_02074_),
    .Y(_02300_));
 sky130_fd_sc_hd__a21bo_1 _09099_ (.A1(_02043_),
    .A2(_02077_),
    .B1_N(_02078_),
    .X(_02301_));
 sky130_fd_sc_hd__or2_1 _09100_ (.A(_02300_),
    .B(_02301_),
    .X(_02303_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(_02301_),
    .B(_02300_),
    .Y(_02304_));
 sky130_fd_sc_hd__nand3_1 _09102_ (.A(_02303_),
    .B(\sq.out[8] ),
    .C(_02304_),
    .Y(_02305_));
 sky130_fd_sc_hd__nand2_1 _09103_ (.A(_02136_),
    .B(_02055_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand2_1 _09104_ (.A(_02305_),
    .B(_02306_),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_1 _09105_ (.A(_02307_),
    .B(_02279_),
    .Y(_02308_));
 sky130_fd_sc_hd__nand3_1 _09106_ (.A(_02289_),
    .B(_02305_),
    .C(_02306_),
    .Y(_02309_));
 sky130_fd_sc_hd__nand3_1 _09107_ (.A(_02261_),
    .B(_02063_),
    .C(_02086_),
    .Y(_02310_));
 sky130_fd_sc_hd__nand3_1 _09108_ (.A(_02262_),
    .B(\sq.out[8] ),
    .C(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__nand2_1 _09109_ (.A(_02136_),
    .B(_02059_),
    .Y(_02312_));
 sky130_fd_sc_hd__nand2_1 _09110_ (.A(_02311_),
    .B(_02312_),
    .Y(_02314_));
 sky130_fd_sc_hd__inv_2 _09111_ (.A(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__nand3_1 _09112_ (.A(_02308_),
    .B(_02309_),
    .C(_02315_),
    .Y(_02316_));
 sky130_fd_sc_hd__inv_2 _09113_ (.A(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__nand2_2 _09114_ (.A(_02299_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_4 _09115_ (.A(_02276_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__o21ai_1 _09116_ (.A1(_02293_),
    .A2(_02296_),
    .B1(_02292_),
    .Y(_02320_));
 sky130_fd_sc_hd__nand2_1 _09117_ (.A(_02320_),
    .B(_02317_),
    .Y(_02321_));
 sky130_fd_sc_hd__inv_2 _09118_ (.A(_02276_),
    .Y(_02322_));
 sky130_fd_sc_hd__and2_1 _09119_ (.A(_02308_),
    .B(_02315_),
    .X(_02323_));
 sky130_fd_sc_hd__nand3_2 _09120_ (.A(_02321_),
    .B(_02322_),
    .C(_02323_),
    .Y(_02325_));
 sky130_fd_sc_hd__a21oi_4 _09121_ (.A1(_02260_),
    .A2(_02319_),
    .B1(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand3_1 _09122_ (.A(_02109_),
    .B(_02085_),
    .C(_01869_),
    .Y(_02327_));
 sky130_fd_sc_hd__clkinvlp_2 _09123_ (.A(_01867_),
    .Y(_02328_));
 sky130_fd_sc_hd__nand2_1 _09124_ (.A(_02108_),
    .B(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _09125_ (.A(_02327_),
    .B(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__nand2_1 _09126_ (.A(_02330_),
    .B(_01363_),
    .Y(_02331_));
 sky130_fd_sc_hd__nand3_2 _09127_ (.A(_02327_),
    .B(\sq.out[12] ),
    .C(_02329_),
    .Y(_02332_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(_02331_),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__nand3_2 _09129_ (.A(_02109_),
    .B(\sq.out[9] ),
    .C(_02085_),
    .Y(_02334_));
 sky130_fd_sc_hd__nand2_1 _09130_ (.A(_02016_),
    .B(\sq.out[10] ),
    .Y(_02336_));
 sky130_fd_sc_hd__nand2_1 _09131_ (.A(\sq.out[9] ),
    .B(_01644_),
    .Y(_02337_));
 sky130_fd_sc_hd__and2_1 _09132_ (.A(_02336_),
    .B(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__nand2_1 _09133_ (.A(_02108_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__nand3_2 _09134_ (.A(_02334_),
    .B(\sq.out[11] ),
    .C(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__nand2_1 _09135_ (.A(_02333_),
    .B(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__inv_2 _09136_ (.A(_02340_),
    .Y(_02342_));
 sky130_fd_sc_hd__nand3_1 _09137_ (.A(_02342_),
    .B(_02331_),
    .C(_02332_),
    .Y(_02343_));
 sky130_fd_sc_hd__nand2_1 _09138_ (.A(_02334_),
    .B(_02339_),
    .Y(_02344_));
 sky130_fd_sc_hd__buf_6 _09139_ (.A(_01531_),
    .X(_02345_));
 sky130_fd_sc_hd__nand2_1 _09140_ (.A(_02344_),
    .B(_02345_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _09141_ (.A(_02108_),
    .B(_02016_),
    .Y(_02348_));
 sky130_fd_sc_hd__and2_1 _09142_ (.A(_02348_),
    .B(_02337_),
    .X(_02349_));
 sky130_fd_sc_hd__nand3_1 _09143_ (.A(_02347_),
    .B(_02340_),
    .C(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand3_1 _09144_ (.A(_02341_),
    .B(_02343_),
    .C(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__nand2_1 _09145_ (.A(_02351_),
    .B(_02341_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _09146_ (.A(_01877_),
    .B(_01864_),
    .Y(_02353_));
 sky130_fd_sc_hd__or2_1 _09147_ (.A(_01868_),
    .B(_02353_),
    .X(_02354_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(_02353_),
    .B(_01868_),
    .Y(_02355_));
 sky130_fd_sc_hd__nand3_1 _09149_ (.A(net105),
    .B(_02354_),
    .C(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__clkinvlp_2 _09150_ (.A(_01871_),
    .Y(_02358_));
 sky130_fd_sc_hd__nand2_1 _09151_ (.A(_02136_),
    .B(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__nand3_2 _09152_ (.A(_02356_),
    .B(_02359_),
    .C(\sq.out[13] ),
    .Y(_02360_));
 sky130_fd_sc_hd__nand2_1 _09153_ (.A(_02356_),
    .B(_02359_),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_1 _09154_ (.A(_02361_),
    .B(_00843_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand3b_1 _09155_ (.A_N(_02332_),
    .B(_02360_),
    .C(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand2_1 _09156_ (.A(_02362_),
    .B(_02360_),
    .Y(_02364_));
 sky130_fd_sc_hd__nand2_1 _09157_ (.A(_02364_),
    .B(_02332_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(_02363_),
    .B(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__inv_2 _09159_ (.A(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__nand2_1 _09160_ (.A(_02352_),
    .B(_02367_),
    .Y(_02369_));
 sky130_fd_sc_hd__nand2_2 _09161_ (.A(_02369_),
    .B(_02365_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand2_1 _09162_ (.A(_02137_),
    .B(_02140_),
    .Y(_02371_));
 sky130_fd_sc_hd__nand2_1 _09163_ (.A(_02371_),
    .B(_01286_),
    .Y(_02372_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(_02372_),
    .B(_02141_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_1 _09165_ (.A(_01885_),
    .B(_01886_),
    .Y(_02374_));
 sky130_fd_sc_hd__xnor2_1 _09166_ (.A(_01878_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand2_1 _09167_ (.A(_02105_),
    .B(_02375_),
    .Y(_02376_));
 sky130_fd_sc_hd__o21ai_2 _09168_ (.A1(_01881_),
    .A2(_02107_),
    .B1(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__or2_1 _09169_ (.A(_01587_),
    .B(_02377_),
    .X(_02378_));
 sky130_fd_sc_hd__nor2_1 _09170_ (.A(_02373_),
    .B(_02378_),
    .Y(_02380_));
 sky130_fd_sc_hd__and2_1 _09171_ (.A(_02378_),
    .B(_02373_),
    .X(_02381_));
 sky130_fd_sc_hd__or2_1 _09172_ (.A(_02380_),
    .B(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__inv_2 _09173_ (.A(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _09174_ (.A(_02377_),
    .B(_01587_),
    .Y(_02384_));
 sky130_fd_sc_hd__inv_2 _09175_ (.A(_02360_),
    .Y(_02385_));
 sky130_fd_sc_hd__a21o_1 _09176_ (.A1(_02378_),
    .A2(_02384_),
    .B1(_02385_),
    .X(_02386_));
 sky130_fd_sc_hd__nand3_1 _09177_ (.A(_02378_),
    .B(_02385_),
    .C(_02384_),
    .Y(_02387_));
 sky130_fd_sc_hd__nand2_1 _09178_ (.A(_02386_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__inv_2 _09179_ (.A(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__nand3_1 _09180_ (.A(_02370_),
    .B(_02383_),
    .C(_02389_),
    .Y(_02391_));
 sky130_fd_sc_hd__o21ba_1 _09181_ (.A1(_02380_),
    .A2(_02386_),
    .B1_N(_02381_),
    .X(_02392_));
 sky130_fd_sc_hd__nand2_2 _09182_ (.A(_02391_),
    .B(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__or2_1 _09183_ (.A(_02141_),
    .B(_02135_),
    .X(_02394_));
 sky130_fd_sc_hd__nand2_1 _09184_ (.A(_02394_),
    .B(_02142_),
    .Y(_02395_));
 sky130_fd_sc_hd__nand2b_1 _09185_ (.A_N(_02152_),
    .B(_02153_),
    .Y(_02396_));
 sky130_fd_sc_hd__nor2_1 _09186_ (.A(_02395_),
    .B(_02396_),
    .Y(_02397_));
 sky130_fd_sc_hd__nand2_1 _09187_ (.A(_02397_),
    .B(_02181_),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2b_4 _09188_ (.A(_02398_),
    .B_N(_02251_),
    .Y(_02399_));
 sky130_fd_sc_hd__nand3_4 _09189_ (.A(_02393_),
    .B(_02319_),
    .C(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _09190_ (.A(_01861_),
    .B(_02111_),
    .Y(_02402_));
 sky130_fd_sc_hd__inv_2 _09191_ (.A(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__inv_2 _09192_ (.A(_02110_),
    .Y(_02404_));
 sky130_fd_sc_hd__nand2_1 _09193_ (.A(_02404_),
    .B(_02085_),
    .Y(_02405_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_02403_),
    .B(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__or2_1 _09195_ (.A(_01861_),
    .B(_02112_),
    .X(_02407_));
 sky130_fd_sc_hd__o22a_1 _09196_ (.A1(_01846_),
    .A2(_01858_),
    .B1(_02116_),
    .B2(_02109_),
    .X(_02408_));
 sky130_fd_sc_hd__nor3b_1 _09197_ (.A(_02407_),
    .B(_02125_),
    .C_N(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(_02409_),
    .B(_02403_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor2_4 _09199_ (.A(_02406_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__nand3_4 _09200_ (.A(_02326_),
    .B(_02400_),
    .C(_02411_),
    .Y(_02413_));
 sky130_fd_sc_hd__buf_6 _09201_ (.A(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__nand2_1 _09202_ (.A(_02326_),
    .B(_02400_),
    .Y(_02415_));
 sky130_fd_sc_hd__inv_2 _09203_ (.A(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__nand2_2 _09204_ (.A(_02414_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__nor2_2 _09205_ (.A(_02125_),
    .B(_02417_),
    .Y(_02418_));
 sky130_fd_sc_hd__xnor2_1 _09206_ (.A(_02116_),
    .B(_02110_),
    .Y(_02419_));
 sky130_fd_sc_hd__nand2_1 _09207_ (.A(_02418_),
    .B(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__or2_4 _09208_ (.A(_02119_),
    .B(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__nor2_1 _09209_ (.A(_02115_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__nor2_1 _09210_ (.A(_02113_),
    .B(_02422_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_1 _09211_ (.A(_02422_),
    .B(_02113_),
    .Y(_02425_));
 sky130_fd_sc_hd__inv_2 _09212_ (.A(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__nor2_1 _09213_ (.A(_02424_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__inv_2 _09214_ (.A(_02427_),
    .Y(_02428_));
 sky130_fd_sc_hd__and2_1 _09215_ (.A(_02421_),
    .B(_02115_),
    .X(_02429_));
 sky130_fd_sc_hd__nor2_1 _09216_ (.A(_02422_),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__inv_2 _09217_ (.A(_02430_),
    .Y(_02431_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(_02420_),
    .B(_02119_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_1 _09219_ (.A(_02421_),
    .B(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__or2_1 _09220_ (.A(_02419_),
    .B(_02418_),
    .X(_02435_));
 sky130_fd_sc_hd__and2_1 _09221_ (.A(_02435_),
    .B(_02420_),
    .X(_02436_));
 sky130_fd_sc_hd__inv_2 _09222_ (.A(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__a21o_1 _09223_ (.A1(_02393_),
    .A2(_02399_),
    .B1(_02260_),
    .X(_02438_));
 sky130_fd_sc_hd__nand2_1 _09224_ (.A(_02321_),
    .B(_02323_),
    .Y(_02439_));
 sky130_fd_sc_hd__inv_6 _09225_ (.A(_02413_),
    .Y(_02440_));
 sky130_fd_sc_hd__buf_6 _09226_ (.A(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__a311o_1 _09227_ (.A1(_02438_),
    .A2(_02317_),
    .A3(_02299_),
    .B1(_02439_),
    .C1(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__nor2_1 _09228_ (.A(_02264_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _09229_ (.A(_02443_),
    .B(_02269_),
    .Y(_02444_));
 sky130_fd_sc_hd__inv_2 _09230_ (.A(_02444_),
    .Y(_02446_));
 sky130_fd_sc_hd__nand2_1 _09231_ (.A(_02446_),
    .B(_02266_),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _09232_ (.A(_02447_),
    .B(_02275_),
    .Y(_02448_));
 sky130_fd_sc_hd__nand3_1 _09233_ (.A(_02446_),
    .B(_02274_),
    .C(_02266_),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_1 _09234_ (.A(_02448_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__clkinvlp_2 _09235_ (.A(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__inv_2 _09236_ (.A(_02395_),
    .Y(_02452_));
 sky130_fd_sc_hd__nand2_1 _09237_ (.A(_02393_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__nand2_1 _09238_ (.A(_02453_),
    .B(_02142_),
    .Y(_02454_));
 sky130_fd_sc_hd__xor2_1 _09239_ (.A(_02396_),
    .B(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__nand2_1 _09240_ (.A(_02455_),
    .B(net114),
    .Y(_02457_));
 sky130_fd_sc_hd__or2_1 _09241_ (.A(_02147_),
    .B(_02414_),
    .X(_02458_));
 sky130_fd_sc_hd__nand2_1 _09242_ (.A(_02457_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__or2_1 _09243_ (.A(\sq.out[18] ),
    .B(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__nand2_1 _09244_ (.A(_02459_),
    .B(\sq.out[18] ),
    .Y(_02461_));
 sky130_fd_sc_hd__or2_1 _09245_ (.A(_02452_),
    .B(_02393_),
    .X(_02462_));
 sky130_fd_sc_hd__nand2_1 _09246_ (.A(_02462_),
    .B(_02453_),
    .Y(_02463_));
 sky130_fd_sc_hd__nand2_1 _09247_ (.A(_02440_),
    .B(_02132_),
    .Y(_02464_));
 sky130_fd_sc_hd__o21ai_2 _09248_ (.A1(_02463_),
    .A2(_02440_),
    .B1(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__or2_1 _09249_ (.A(_01240_),
    .B(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__inv_2 _09250_ (.A(_02466_),
    .Y(_02468_));
 sky130_fd_sc_hd__a21o_1 _09251_ (.A1(_02460_),
    .A2(_02461_),
    .B1(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__nand3_1 _09252_ (.A(_02468_),
    .B(_02460_),
    .C(_02461_),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_1 _09253_ (.A(_02469_),
    .B(_02470_),
    .Y(_02471_));
 sky130_fd_sc_hd__inv_2 _09254_ (.A(_02180_),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(_02393_),
    .B(_02397_),
    .Y(_02473_));
 sky130_fd_sc_hd__inv_2 _09256_ (.A(_02154_),
    .Y(_02474_));
 sky130_fd_sc_hd__nand2_1 _09257_ (.A(_02473_),
    .B(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__or2_1 _09258_ (.A(_02472_),
    .B(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_02475_),
    .B(_02472_),
    .Y(_02477_));
 sky130_fd_sc_hd__nand3_1 _09260_ (.A(_02476_),
    .B(_02414_),
    .C(_02477_),
    .Y(_02479_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(_02440_),
    .B(_02174_),
    .Y(_02480_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(_02479_),
    .B(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__or2_1 _09263_ (.A(_05130_),
    .B(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__nand2_1 _09264_ (.A(_02481_),
    .B(_05130_),
    .Y(_02483_));
 sky130_fd_sc_hd__nand2_1 _09265_ (.A(_02482_),
    .B(_02483_),
    .Y(_02484_));
 sky130_fd_sc_hd__nor2_1 _09266_ (.A(_02461_),
    .B(_02484_),
    .Y(_02485_));
 sky130_fd_sc_hd__nand2_1 _09267_ (.A(_02484_),
    .B(_02461_),
    .Y(_02486_));
 sky130_fd_sc_hd__nand2b_1 _09268_ (.A_N(_02485_),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__nor2_1 _09269_ (.A(_02471_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__inv_2 _09270_ (.A(_02488_),
    .Y(_02490_));
 sky130_fd_sc_hd__nor2_2 _09271_ (.A(\sq.out[8] ),
    .B(_02414_),
    .Y(_02491_));
 sky130_fd_sc_hd__nand3_1 _09272_ (.A(_02491_),
    .B(_01644_),
    .C(\sq.out[9] ),
    .Y(_02492_));
 sky130_fd_sc_hd__clkinvlp_2 _09273_ (.A(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hd__buf_6 _09274_ (.A(_02414_),
    .X(_02494_));
 sky130_fd_sc_hd__buf_6 _09275_ (.A(_02494_),
    .X(\sq.out[7] ));
 sky130_fd_sc_hd__buf_6 _09276_ (.A(_02016_),
    .X(_02495_));
 sky130_fd_sc_hd__nand2_1 _09277_ (.A(_02334_),
    .B(_02348_),
    .Y(_02496_));
 sky130_fd_sc_hd__a21oi_1 _09278_ (.A1(\sq.out[7] ),
    .A2(_02495_),
    .B1(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__buf_6 _09279_ (.A(_02136_),
    .X(_02498_));
 sky130_fd_sc_hd__nand3_2 _09280_ (.A(_02416_),
    .B(_02498_),
    .C(_02411_),
    .Y(_02500_));
 sky130_fd_sc_hd__nand2_1 _09281_ (.A(_02494_),
    .B(_02496_),
    .Y(_02501_));
 sky130_fd_sc_hd__nand2_1 _09282_ (.A(_02500_),
    .B(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__nand2_1 _09283_ (.A(_02502_),
    .B(\sq.out[10] ),
    .Y(_02503_));
 sky130_fd_sc_hd__buf_6 _09284_ (.A(_01644_),
    .X(_02504_));
 sky130_fd_sc_hd__nand3_1 _09285_ (.A(_02500_),
    .B(_02504_),
    .C(_02501_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_1 _09286_ (.A(_02503_),
    .B(_02505_),
    .Y(_02506_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_02491_),
    .B(\sq.out[9] ),
    .Y(_02507_));
 sky130_fd_sc_hd__nand2_1 _09288_ (.A(_02506_),
    .B(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__o21ai_2 _09289_ (.A1(_02493_),
    .A2(_02497_),
    .B1(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(_02491_),
    .B(_02016_),
    .Y(_02511_));
 sky130_fd_sc_hd__or2b_1 _09291_ (.A(_02338_),
    .B_N(_02413_),
    .X(_02512_));
 sky130_fd_sc_hd__nand2_1 _09292_ (.A(_02511_),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__nand2_1 _09293_ (.A(_02513_),
    .B(\sq.out[11] ),
    .Y(_02514_));
 sky130_fd_sc_hd__nand3_1 _09294_ (.A(_02511_),
    .B(_02512_),
    .C(_02345_),
    .Y(_02515_));
 sky130_fd_sc_hd__nand2_1 _09295_ (.A(_02514_),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__nand2_1 _09296_ (.A(_02516_),
    .B(_02503_),
    .Y(_02517_));
 sky130_fd_sc_hd__nand3b_1 _09297_ (.A_N(_02503_),
    .B(_02514_),
    .C(_02515_),
    .Y(_02518_));
 sky130_fd_sc_hd__nand3_1 _09298_ (.A(_02509_),
    .B(_02517_),
    .C(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__nand2_1 _09299_ (.A(_02519_),
    .B(_02517_),
    .Y(_02520_));
 sky130_fd_sc_hd__a21o_1 _09300_ (.A1(_02347_),
    .A2(_02340_),
    .B1(_02349_),
    .X(_02522_));
 sky130_fd_sc_hd__a21o_1 _09301_ (.A1(_02350_),
    .A2(_02522_),
    .B1(_02440_),
    .X(_02523_));
 sky130_fd_sc_hd__nand2_1 _09302_ (.A(_02441_),
    .B(_02344_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand3_1 _09303_ (.A(_02523_),
    .B(_02524_),
    .C(\sq.out[12] ),
    .Y(_02525_));
 sky130_fd_sc_hd__a21o_1 _09304_ (.A1(_02341_),
    .A2(_02343_),
    .B1(_02350_),
    .X(_02526_));
 sky130_fd_sc_hd__nand3_1 _09305_ (.A(_02413_),
    .B(_02351_),
    .C(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2_1 _09306_ (.A(_02440_),
    .B(_02330_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand2_1 _09307_ (.A(_02527_),
    .B(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__inv_2 _09308_ (.A(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__nand2_1 _09309_ (.A(_02530_),
    .B(\sq.out[13] ),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _09310_ (.A(_02529_),
    .B(_00843_),
    .Y(_02533_));
 sky130_fd_sc_hd__nand2_1 _09311_ (.A(_02531_),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__or2_1 _09312_ (.A(_02525_),
    .B(_02534_),
    .X(_02535_));
 sky130_fd_sc_hd__nand2_1 _09313_ (.A(_02534_),
    .B(_02525_),
    .Y(_02536_));
 sky130_fd_sc_hd__nand2_1 _09314_ (.A(_02535_),
    .B(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__inv_2 _09315_ (.A(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__nand2_1 _09316_ (.A(_02523_),
    .B(_02524_),
    .Y(_02539_));
 sky130_fd_sc_hd__nand2_1 _09317_ (.A(_02539_),
    .B(_01363_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand2_1 _09318_ (.A(_02540_),
    .B(_02525_),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _09319_ (.A(_02514_),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_1 _09320_ (.A(_02541_),
    .B(_02514_),
    .Y(_02544_));
 sky130_fd_sc_hd__inv_2 _09321_ (.A(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _09322_ (.A(_02542_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand3_1 _09323_ (.A(_02520_),
    .B(_02538_),
    .C(_02546_),
    .Y(_02547_));
 sky130_fd_sc_hd__a21boi_1 _09324_ (.A1(_02545_),
    .A2(_02535_),
    .B1_N(_02536_),
    .Y(_02548_));
 sky130_fd_sc_hd__nand2_1 _09325_ (.A(_02547_),
    .B(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__or2_1 _09326_ (.A(_02367_),
    .B(_02352_),
    .X(_02550_));
 sky130_fd_sc_hd__nand2_1 _09327_ (.A(_02550_),
    .B(_02369_),
    .Y(_02551_));
 sky130_fd_sc_hd__nand2_1 _09328_ (.A(_02440_),
    .B(_02361_),
    .Y(_02552_));
 sky130_fd_sc_hd__o21ai_2 _09329_ (.A1(_02551_),
    .A2(_02440_),
    .B1(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__or2_1 _09330_ (.A(_01587_),
    .B(_02553_),
    .X(_02555_));
 sky130_fd_sc_hd__xor2_1 _09331_ (.A(_02388_),
    .B(_02370_),
    .X(_02556_));
 sky130_fd_sc_hd__nand2_1 _09332_ (.A(_02440_),
    .B(_02377_),
    .Y(_02557_));
 sky130_fd_sc_hd__o21ai_2 _09333_ (.A1(_02556_),
    .A2(_02440_),
    .B1(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__or2_1 _09334_ (.A(_01286_),
    .B(_02558_),
    .X(_02559_));
 sky130_fd_sc_hd__nand2_1 _09335_ (.A(_02558_),
    .B(_01286_),
    .Y(_02560_));
 sky130_fd_sc_hd__nand2_1 _09336_ (.A(_02559_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__or2_1 _09337_ (.A(_02555_),
    .B(_02561_),
    .X(_02562_));
 sky130_fd_sc_hd__nand2_1 _09338_ (.A(_02561_),
    .B(_02555_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand2_1 _09339_ (.A(_02562_),
    .B(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__inv_2 _09340_ (.A(_02564_),
    .Y(_02566_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_02553_),
    .B(_01587_),
    .Y(_02567_));
 sky130_fd_sc_hd__nand2_1 _09342_ (.A(_02555_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__or2_1 _09343_ (.A(_02531_),
    .B(_02568_),
    .X(_02569_));
 sky130_fd_sc_hd__nand2_1 _09344_ (.A(_02568_),
    .B(_02531_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _09345_ (.A(_02569_),
    .B(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__inv_2 _09346_ (.A(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__nand3_2 _09347_ (.A(_02549_),
    .B(_02566_),
    .C(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__o21a_1 _09348_ (.A1(_02570_),
    .A2(_02564_),
    .B1(_02563_),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_2 _09349_ (.A(_02573_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__a21bo_1 _09350_ (.A1(_02370_),
    .A2(_02387_),
    .B1_N(_02386_),
    .X(_02577_));
 sky130_fd_sc_hd__xor2_1 _09351_ (.A(_02382_),
    .B(_02577_),
    .X(_02578_));
 sky130_fd_sc_hd__nand2_1 _09352_ (.A(_02494_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__o21ai_1 _09353_ (.A1(_02371_),
    .A2(_02494_),
    .B1(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__nand2_1 _09354_ (.A(_02580_),
    .B(\sq.out[16] ),
    .Y(_02581_));
 sky130_fd_sc_hd__nand2_1 _09355_ (.A(_02465_),
    .B(_01240_),
    .Y(_02582_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(_02466_),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hd__nor2_1 _09357_ (.A(_02581_),
    .B(_02583_),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_1 _09358_ (.A(_02583_),
    .B(_02581_),
    .Y(_02585_));
 sky130_fd_sc_hd__or2b_1 _09359_ (.A(_02584_),
    .B_N(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__clkinvlp_2 _09360_ (.A(_02586_),
    .Y(_02588_));
 sky130_fd_sc_hd__or2_1 _09361_ (.A(\sq.out[16] ),
    .B(_02580_),
    .X(_02589_));
 sky130_fd_sc_hd__nand2_1 _09362_ (.A(_02589_),
    .B(_02581_),
    .Y(_02590_));
 sky130_fd_sc_hd__or2_1 _09363_ (.A(_02559_),
    .B(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__nand2_1 _09364_ (.A(_02590_),
    .B(_02559_),
    .Y(_02592_));
 sky130_fd_sc_hd__nand2_1 _09365_ (.A(_02591_),
    .B(_02592_),
    .Y(_02593_));
 sky130_fd_sc_hd__inv_2 _09366_ (.A(_02593_),
    .Y(_02594_));
 sky130_fd_sc_hd__nand3_4 _09367_ (.A(_02575_),
    .B(_02588_),
    .C(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__nor2_4 _09368_ (.A(_02490_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__or2_1 _09369_ (.A(_02269_),
    .B(_02443_),
    .X(_02597_));
 sky130_fd_sc_hd__nand3_1 _09370_ (.A(_02597_),
    .B(_02266_),
    .C(_02444_),
    .Y(_02599_));
 sky130_fd_sc_hd__a21o_1 _09371_ (.A1(_02438_),
    .A2(_02299_),
    .B1(_02320_),
    .X(_02600_));
 sky130_fd_sc_hd__and2_1 _09372_ (.A(_02308_),
    .B(_02309_),
    .X(_02601_));
 sky130_fd_sc_hd__a21oi_1 _09373_ (.A1(_02600_),
    .A2(_02601_),
    .B1(_02441_),
    .Y(_02602_));
 sky130_fd_sc_hd__nand2_1 _09374_ (.A(_02602_),
    .B(_02308_),
    .Y(_02603_));
 sky130_fd_sc_hd__xor2_1 _09375_ (.A(_02315_),
    .B(_02603_),
    .X(_02604_));
 sky130_fd_sc_hd__and2_1 _09376_ (.A(_02442_),
    .B(_02264_),
    .X(_02605_));
 sky130_fd_sc_hd__or2_1 _09377_ (.A(_02443_),
    .B(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__or2_1 _09378_ (.A(_02604_),
    .B(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__nor2_1 _09379_ (.A(_02599_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hd__a31o_1 _09380_ (.A1(_02393_),
    .A2(_02181_),
    .A3(_02397_),
    .B1(_02186_),
    .X(_02610_));
 sky130_fd_sc_hd__inv_2 _09381_ (.A(_02250_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(_02610_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__inv_2 _09383_ (.A(_02254_),
    .Y(_02613_));
 sky130_fd_sc_hd__nand2_1 _09384_ (.A(_02612_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(_02614_),
    .B(_02225_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _09386_ (.A(_02615_),
    .B(_02221_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _09387_ (.A(_02616_),
    .B(_02211_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand3_1 _09388_ (.A(_02615_),
    .B(_02210_),
    .C(_02221_),
    .Y(_02618_));
 sky130_fd_sc_hd__nand2_1 _09389_ (.A(_02617_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__nand2_1 _09390_ (.A(_02619_),
    .B(\sq.out[7] ),
    .Y(_02621_));
 sky130_fd_sc_hd__or2_1 _09391_ (.A(_02205_),
    .B(_02494_),
    .X(_02622_));
 sky130_fd_sc_hd__nand2_1 _09392_ (.A(_02621_),
    .B(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_1 _09393_ (.A(_02623_),
    .B(_02071_),
    .Y(_02624_));
 sky130_fd_sc_hd__xor2_1 _09394_ (.A(_02298_),
    .B(_02438_),
    .X(_02625_));
 sky130_fd_sc_hd__or2_1 _09395_ (.A(_02287_),
    .B(net114),
    .X(_02626_));
 sky130_fd_sc_hd__o21a_1 _09396_ (.A1(_02441_),
    .A2(_02625_),
    .B1(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__nand2_1 _09397_ (.A(_02624_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__inv_2 _09398_ (.A(_02627_),
    .Y(_02629_));
 sky130_fd_sc_hd__nand3_1 _09399_ (.A(_02623_),
    .B(_02071_),
    .C(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2_1 _09400_ (.A(_02628_),
    .B(_02630_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand3_1 _09401_ (.A(_02621_),
    .B(_01081_),
    .C(_02622_),
    .Y(_02633_));
 sky130_fd_sc_hd__nand2_1 _09402_ (.A(_02624_),
    .B(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__nand3_1 _09403_ (.A(_02612_),
    .B(_02224_),
    .C(_02613_),
    .Y(_02635_));
 sky130_fd_sc_hd__nand3_1 _09404_ (.A(_02615_),
    .B(net114),
    .C(_02635_),
    .Y(_02636_));
 sky130_fd_sc_hd__or2_1 _09405_ (.A(_02194_),
    .B(net114),
    .X(_02637_));
 sky130_fd_sc_hd__nand2_1 _09406_ (.A(_02636_),
    .B(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__inv_2 _09407_ (.A(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hd__nand2_1 _09408_ (.A(_02639_),
    .B(\sq.out[23] ),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _09409_ (.A(_02634_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__nand3b_1 _09410_ (.A_N(_02640_),
    .B(_02624_),
    .C(_02633_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _09411_ (.A(_02641_),
    .B(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__nor2_1 _09412_ (.A(_02632_),
    .B(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__o21ai_1 _09413_ (.A1(_02601_),
    .A2(_02600_),
    .B1(_02602_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand2_1 _09414_ (.A(_02441_),
    .B(_02307_),
    .Y(_02647_));
 sky130_fd_sc_hd__nand2_1 _09415_ (.A(_02646_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__a21bo_1 _09416_ (.A1(_02438_),
    .A2(_02297_),
    .B1_N(_02296_),
    .X(_02649_));
 sky130_fd_sc_hd__or2b_1 _09417_ (.A(_02649_),
    .B_N(_02293_),
    .X(_02650_));
 sky130_fd_sc_hd__nand2_1 _09418_ (.A(_02650_),
    .B(\sq.out[7] ),
    .Y(_02651_));
 sky130_fd_sc_hd__a31o_1 _09419_ (.A1(_02292_),
    .A2(_02288_),
    .A3(_02649_),
    .B1(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__nand2_1 _09420_ (.A(_02441_),
    .B(_02279_),
    .Y(_02654_));
 sky130_fd_sc_hd__nand2_1 _09421_ (.A(_02652_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__nand2_1 _09422_ (.A(_02655_),
    .B(_02629_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand3_1 _09423_ (.A(_02652_),
    .B(_02627_),
    .C(_02654_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(_02656_),
    .B(_02657_),
    .Y(_02658_));
 sky130_fd_sc_hd__nor2_1 _09425_ (.A(_02648_),
    .B(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__nand3_1 _09426_ (.A(_02608_),
    .B(_02645_),
    .C(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__inv_2 _09427_ (.A(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__nand2_1 _09428_ (.A(_02610_),
    .B(_02249_),
    .Y(_02662_));
 sky130_fd_sc_hd__nand2_1 _09429_ (.A(_02662_),
    .B(_02246_),
    .Y(_02663_));
 sky130_fd_sc_hd__nand2_1 _09430_ (.A(_02663_),
    .B(_02242_),
    .Y(_02665_));
 sky130_fd_sc_hd__nand3_1 _09431_ (.A(_02662_),
    .B(_02241_),
    .C(_02246_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(_02665_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand2_1 _09433_ (.A(_02667_),
    .B(_02494_),
    .Y(_02668_));
 sky130_fd_sc_hd__or2_1 _09434_ (.A(_02235_),
    .B(_02494_),
    .X(_02669_));
 sky130_fd_sc_hd__nand2_1 _09435_ (.A(_02668_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand2_1 _09436_ (.A(_02670_),
    .B(\sq.out[22] ),
    .Y(_02671_));
 sky130_fd_sc_hd__nand3_1 _09437_ (.A(_02668_),
    .B(_02009_),
    .C(_02669_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand2_1 _09438_ (.A(_02671_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__or2_1 _09439_ (.A(_02249_),
    .B(_02610_),
    .X(_02674_));
 sky130_fd_sc_hd__nand3_1 _09440_ (.A(_02674_),
    .B(_02494_),
    .C(_02662_),
    .Y(_02676_));
 sky130_fd_sc_hd__or2_1 _09441_ (.A(_02232_),
    .B(net114),
    .X(_02677_));
 sky130_fd_sc_hd__nand3_1 _09442_ (.A(_02676_),
    .B(\sq.out[21] ),
    .C(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__nand2_1 _09443_ (.A(_02673_),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand3b_1 _09444_ (.A_N(_02678_),
    .B(_02671_),
    .C(_02672_),
    .Y(_02680_));
 sky130_fd_sc_hd__nand2_1 _09445_ (.A(_02679_),
    .B(_02680_),
    .Y(_02681_));
 sky130_fd_sc_hd__nand2_1 _09446_ (.A(_02638_),
    .B(_01993_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand3b_1 _09447_ (.A_N(_02671_),
    .B(_02640_),
    .C(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _09448_ (.A(_02640_),
    .B(_02682_),
    .Y(_02684_));
 sky130_fd_sc_hd__nand2_1 _09449_ (.A(_02684_),
    .B(_02671_),
    .Y(_02685_));
 sky130_fd_sc_hd__nand2_1 _09450_ (.A(_02683_),
    .B(_02685_),
    .Y(_02687_));
 sky130_fd_sc_hd__nor2_1 _09451_ (.A(_02681_),
    .B(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_02477_),
    .B(_02177_),
    .Y(_02689_));
 sky130_fd_sc_hd__xor2_1 _09453_ (.A(_02173_),
    .B(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__nand2_1 _09454_ (.A(_02690_),
    .B(_02494_),
    .Y(_02691_));
 sky130_fd_sc_hd__o21ai_2 _09455_ (.A1(_02159_),
    .A2(_02494_),
    .B1(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _09456_ (.A(_02692_),
    .B(\sq.out[20] ),
    .Y(_02693_));
 sky130_fd_sc_hd__nand2_1 _09457_ (.A(_02676_),
    .B(_02677_),
    .Y(_02694_));
 sky130_fd_sc_hd__nand2_1 _09458_ (.A(_02694_),
    .B(_00455_),
    .Y(_02695_));
 sky130_fd_sc_hd__nand2_1 _09459_ (.A(_02695_),
    .B(_02678_),
    .Y(_02696_));
 sky130_fd_sc_hd__nor2_1 _09460_ (.A(_02693_),
    .B(_02696_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_1 _09461_ (.A(_02696_),
    .B(_02693_),
    .Y(_02699_));
 sky130_fd_sc_hd__or2b_1 _09462_ (.A(_02698_),
    .B_N(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__or2_1 _09463_ (.A(\sq.out[20] ),
    .B(_02692_),
    .X(_02701_));
 sky130_fd_sc_hd__nand2_1 _09464_ (.A(_02701_),
    .B(_02693_),
    .Y(_02702_));
 sky130_fd_sc_hd__nand2_1 _09465_ (.A(_02702_),
    .B(_02482_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand3b_1 _09466_ (.A_N(_02482_),
    .B(_02701_),
    .C(_02693_),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2_1 _09467_ (.A(_02703_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__nor2_1 _09468_ (.A(_02705_),
    .B(_02700_),
    .Y(_02706_));
 sky130_fd_sc_hd__nand2_1 _09469_ (.A(_02706_),
    .B(_02688_),
    .Y(_02707_));
 sky130_fd_sc_hd__clkinvlp_2 _09470_ (.A(_02707_),
    .Y(_02709_));
 sky130_fd_sc_hd__nand3_4 _09471_ (.A(_02596_),
    .B(_02661_),
    .C(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__o21ai_1 _09472_ (.A1(_02632_),
    .A2(_02641_),
    .B1(_02628_),
    .Y(_02711_));
 sky130_fd_sc_hd__nand2_1 _09473_ (.A(_02711_),
    .B(_02659_),
    .Y(_02712_));
 sky130_fd_sc_hd__and3_1 _09474_ (.A(_02656_),
    .B(_02646_),
    .C(_02647_),
    .X(_02713_));
 sky130_fd_sc_hd__nand3_1 _09475_ (.A(_02712_),
    .B(_02608_),
    .C(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__o21ai_1 _09476_ (.A1(_02698_),
    .A2(_02703_),
    .B1(_02699_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(_02688_),
    .B(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hd__nor2_1 _09478_ (.A(_02671_),
    .B(_02684_),
    .Y(_02717_));
 sky130_fd_sc_hd__o21a_1 _09479_ (.A1(_02679_),
    .A2(_02717_),
    .B1(_02685_),
    .X(_02718_));
 sky130_fd_sc_hd__nand2_1 _09480_ (.A(_02716_),
    .B(_02718_),
    .Y(_02720_));
 sky130_fd_sc_hd__o21ai_1 _09481_ (.A1(_02592_),
    .A2(_02584_),
    .B1(_02585_),
    .Y(_02721_));
 sky130_fd_sc_hd__o21ai_1 _09482_ (.A1(_02485_),
    .A2(_02469_),
    .B1(_02486_),
    .Y(_02722_));
 sky130_fd_sc_hd__a21oi_2 _09483_ (.A1(_02488_),
    .A2(_02721_),
    .B1(_02722_),
    .Y(_02723_));
 sky130_fd_sc_hd__nor2_1 _09484_ (.A(_02723_),
    .B(_02707_),
    .Y(_02724_));
 sky130_fd_sc_hd__nor2_1 _09485_ (.A(_02720_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__nor2_1 _09486_ (.A(_02660_),
    .B(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__nor2_2 _09487_ (.A(_02726_),
    .B(_02714_),
    .Y(_02727_));
 sky130_fd_sc_hd__a21o_1 _09488_ (.A1(_02421_),
    .A2(_02111_),
    .B1(_01861_),
    .X(_02728_));
 sky130_fd_sc_hd__or3_1 _09489_ (.A(_01861_),
    .B(_01862_),
    .C(_02110_),
    .X(_02729_));
 sky130_fd_sc_hd__nand2_1 _09490_ (.A(_02728_),
    .B(_02729_),
    .Y(_02731_));
 sky130_fd_sc_hd__or3_1 _09491_ (.A(_01861_),
    .B(_02112_),
    .C(_02422_),
    .X(_02732_));
 sky130_fd_sc_hd__nand2_1 _09492_ (.A(_02417_),
    .B(_02125_),
    .Y(_02733_));
 sky130_fd_sc_hd__and2b_1 _09493_ (.A_N(_02418_),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__nand2_1 _09494_ (.A(_02436_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__nor3_1 _09495_ (.A(_02433_),
    .B(_02735_),
    .C(_02431_),
    .Y(_02736_));
 sky130_fd_sc_hd__nand3_1 _09496_ (.A(_02450_),
    .B(_02427_),
    .C(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__nor2_1 _09497_ (.A(_02732_),
    .B(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__a21o_1 _09498_ (.A1(_02421_),
    .A2(_02111_),
    .B1(_01861_),
    .X(_02739_));
 sky130_fd_sc_hd__nand2_1 _09499_ (.A(_02404_),
    .B(_02085_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand3_1 _09500_ (.A(_02738_),
    .B(_02739_),
    .C(_02740_),
    .Y(_02742_));
 sky130_fd_sc_hd__nor2_2 _09501_ (.A(_02731_),
    .B(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__nand3_4 _09502_ (.A(_02710_),
    .B(_02727_),
    .C(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand3_4 _09503_ (.A(_02744_),
    .B(_02710_),
    .C(_02727_),
    .Y(_02745_));
 sky130_fd_sc_hd__nor2_2 _09504_ (.A(_02451_),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__nand2_1 _09505_ (.A(_02746_),
    .B(_02734_),
    .Y(_02747_));
 sky130_fd_sc_hd__or2_1 _09506_ (.A(_02437_),
    .B(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__or2_1 _09507_ (.A(_02433_),
    .B(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__or2_1 _09508_ (.A(_02431_),
    .B(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__or2_1 _09509_ (.A(_02428_),
    .B(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__nand2_1 _09510_ (.A(_02750_),
    .B(_02428_),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _09511_ (.A(_02751_),
    .B(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _09512_ (.A(_02748_),
    .B(_02433_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _09513_ (.A(_02749_),
    .B(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__nand2_1 _09514_ (.A(_02749_),
    .B(_02431_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_1 _09515_ (.A(_02750_),
    .B(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__or2_1 _09516_ (.A(_02756_),
    .B(_02758_),
    .X(_02759_));
 sky130_fd_sc_hd__nor2_1 _09517_ (.A(_02732_),
    .B(_02751_),
    .Y(_02760_));
 sky130_fd_sc_hd__and2_1 _09518_ (.A(_02751_),
    .B(_02732_),
    .X(_02761_));
 sky130_fd_sc_hd__or2_1 _09519_ (.A(_02760_),
    .B(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__or3_4 _09520_ (.A(_02754_),
    .B(_02759_),
    .C(_02762_),
    .X(_02764_));
 sky130_fd_sc_hd__inv_2 _09521_ (.A(_02744_),
    .Y(_02765_));
 sky130_fd_sc_hd__nand3_1 _09522_ (.A(_02765_),
    .B(_02498_),
    .C(_02441_),
    .Y(_02766_));
 sky130_fd_sc_hd__buf_6 _09523_ (.A(_02744_),
    .X(_02767_));
 sky130_fd_sc_hd__nand2_1 _09524_ (.A(_02767_),
    .B(_02496_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand2_1 _09525_ (.A(_02766_),
    .B(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2_1 _09526_ (.A(_02769_),
    .B(\sq.out[10] ),
    .Y(_02770_));
 sky130_fd_sc_hd__nand3_1 _09527_ (.A(_02766_),
    .B(_02504_),
    .C(_02768_),
    .Y(_02771_));
 sky130_fd_sc_hd__nand2_1 _09528_ (.A(_02770_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__buf_6 _09529_ (.A(_02765_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_1 _09530_ (.A(_02773_),
    .B(_02441_),
    .Y(_02775_));
 sky130_fd_sc_hd__nand2_1 _09531_ (.A(_02441_),
    .B(\sq.out[8] ),
    .Y(_02776_));
 sky130_fd_sc_hd__nand2_1 _09532_ (.A(\sq.out[7] ),
    .B(_02498_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _09533_ (.A(_02776_),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand2_1 _09534_ (.A(_02767_),
    .B(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_02775_),
    .B(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2_2 _09536_ (.A(_02780_),
    .B(\sq.out[9] ),
    .Y(_02781_));
 sky130_fd_sc_hd__nand2_2 _09537_ (.A(_02772_),
    .B(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__a21oi_1 _09538_ (.A1(_02775_),
    .A2(_02779_),
    .B1(_02495_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand3_1 _09539_ (.A(_02770_),
    .B(_02783_),
    .C(_02771_),
    .Y(_02784_));
 sky130_fd_sc_hd__o21ai_1 _09540_ (.A1(\sq.out[7] ),
    .A2(_02773_),
    .B1(_02777_),
    .Y(_02786_));
 sky130_fd_sc_hd__nand3_1 _09541_ (.A(_02775_),
    .B(_02495_),
    .C(_02779_),
    .Y(_02787_));
 sky130_fd_sc_hd__nand3b_2 _09542_ (.A_N(_02786_),
    .B(_02781_),
    .C(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand3_2 _09543_ (.A(_02782_),
    .B(_02784_),
    .C(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__inv_2 _09544_ (.A(_02789_),
    .Y(_02790_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_02508_),
    .B(_02492_),
    .Y(_02791_));
 sky130_fd_sc_hd__or2_1 _09546_ (.A(_02497_),
    .B(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__nand2_1 _09547_ (.A(_02791_),
    .B(_02497_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand3_1 _09548_ (.A(_02767_),
    .B(_02792_),
    .C(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__inv_2 _09549_ (.A(_02502_),
    .Y(_02795_));
 sky130_fd_sc_hd__nand2_1 _09550_ (.A(_02773_),
    .B(_02795_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_1 _09551_ (.A(_02794_),
    .B(_02797_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_1 _09552_ (.A(_02798_),
    .B(_02345_),
    .Y(_02799_));
 sky130_fd_sc_hd__nand3_1 _09553_ (.A(_02794_),
    .B(_02797_),
    .C(\sq.out[11] ),
    .Y(_02800_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(_02799_),
    .B(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__nor2_1 _09555_ (.A(_02770_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(_02801_),
    .B(_02770_),
    .Y(_02803_));
 sky130_fd_sc_hd__nor2b_2 _09557_ (.A(_02802_),
    .B_N(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__nand2_1 _09558_ (.A(_02790_),
    .B(_02804_),
    .Y(_02805_));
 sky130_fd_sc_hd__o21a_1 _09559_ (.A1(_02802_),
    .A2(_02782_),
    .B1(_02803_),
    .X(_02806_));
 sky130_fd_sc_hd__nand2_1 _09560_ (.A(_02805_),
    .B(_02806_),
    .Y(_02808_));
 sky130_fd_sc_hd__or2_1 _09561_ (.A(_02546_),
    .B(_02520_),
    .X(_02809_));
 sky130_fd_sc_hd__nand2_1 _09562_ (.A(_02520_),
    .B(_02546_),
    .Y(_02810_));
 sky130_fd_sc_hd__nand2_1 _09563_ (.A(_02809_),
    .B(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand2_1 _09564_ (.A(_02773_),
    .B(_02539_),
    .Y(_02812_));
 sky130_fd_sc_hd__o21ai_2 _09565_ (.A1(_02811_),
    .A2(_02773_),
    .B1(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__or2_1 _09566_ (.A(_00843_),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__nand2_1 _09567_ (.A(_02813_),
    .B(_00844_),
    .Y(_02815_));
 sky130_fd_sc_hd__nand2_1 _09568_ (.A(_02517_),
    .B(_02518_),
    .Y(_02816_));
 sky130_fd_sc_hd__xnor2_1 _09569_ (.A(_02509_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__nand2_1 _09570_ (.A(_02744_),
    .B(_02817_),
    .Y(_02819_));
 sky130_fd_sc_hd__o21ai_1 _09571_ (.A1(_02513_),
    .A2(_02744_),
    .B1(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__or2_1 _09572_ (.A(_01363_),
    .B(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__a21bo_1 _09573_ (.A1(_02814_),
    .A2(_02815_),
    .B1_N(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__nand3b_1 _09574_ (.A_N(_02821_),
    .B(_02814_),
    .C(_02815_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _09575_ (.A(_02822_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__inv_2 _09576_ (.A(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__buf_6 _09577_ (.A(_01363_),
    .X(_02826_));
 sky130_fd_sc_hd__nand2_1 _09578_ (.A(_02820_),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__nand2_1 _09579_ (.A(_02821_),
    .B(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__and2_1 _09580_ (.A(_02828_),
    .B(_02800_),
    .X(_02830_));
 sky130_fd_sc_hd__inv_2 _09581_ (.A(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__or2_1 _09582_ (.A(_02800_),
    .B(_02828_),
    .X(_02832_));
 sky130_fd_sc_hd__nand2_1 _09583_ (.A(_02831_),
    .B(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__inv_2 _09584_ (.A(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__nand3_1 _09585_ (.A(_02808_),
    .B(_02825_),
    .C(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__a21boi_1 _09586_ (.A1(_02823_),
    .A2(_02830_),
    .B1_N(_02822_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand2_1 _09587_ (.A(_02835_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__xor2_1 _09588_ (.A(_02571_),
    .B(_02549_),
    .X(_02838_));
 sky130_fd_sc_hd__nand2_1 _09589_ (.A(_02773_),
    .B(_02553_),
    .Y(_02839_));
 sky130_fd_sc_hd__o21ai_2 _09590_ (.A1(_02838_),
    .A2(_02773_),
    .B1(_02839_),
    .Y(_02841_));
 sky130_fd_sc_hd__or2_1 _09591_ (.A(_01286_),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__buf_6 _09592_ (.A(_01286_),
    .X(_02843_));
 sky130_fd_sc_hd__nand2_1 _09593_ (.A(_02841_),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__nand2_1 _09594_ (.A(_02842_),
    .B(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _09595_ (.A(_02810_),
    .B(_02544_),
    .Y(_02846_));
 sky130_fd_sc_hd__nand2_1 _09596_ (.A(_02846_),
    .B(_02538_),
    .Y(_02847_));
 sky130_fd_sc_hd__or2_1 _09597_ (.A(_02538_),
    .B(_02846_),
    .X(_02848_));
 sky130_fd_sc_hd__nor2_1 _09598_ (.A(_02530_),
    .B(_02767_),
    .Y(_02849_));
 sky130_fd_sc_hd__a31o_1 _09599_ (.A1(_02767_),
    .A2(_02847_),
    .A3(_02848_),
    .B1(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__or2_1 _09600_ (.A(_01587_),
    .B(_02850_),
    .X(_02852_));
 sky130_fd_sc_hd__or2_1 _09601_ (.A(_02845_),
    .B(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__nand2_1 _09602_ (.A(_02852_),
    .B(_02845_),
    .Y(_02854_));
 sky130_fd_sc_hd__nand2_1 _09603_ (.A(_02853_),
    .B(_02854_),
    .Y(_02855_));
 sky130_fd_sc_hd__buf_6 _09604_ (.A(_01587_),
    .X(_02856_));
 sky130_fd_sc_hd__nand2_1 _09605_ (.A(_02850_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__nand2_1 _09606_ (.A(_02852_),
    .B(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hd__or2_1 _09607_ (.A(_02814_),
    .B(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__nand2_1 _09608_ (.A(_02858_),
    .B(_02814_),
    .Y(_02860_));
 sky130_fd_sc_hd__nand2_1 _09609_ (.A(_02859_),
    .B(_02860_),
    .Y(_02861_));
 sky130_fd_sc_hd__nor2_1 _09610_ (.A(_02855_),
    .B(_02861_),
    .Y(_02863_));
 sky130_fd_sc_hd__nand2_1 _09611_ (.A(_02837_),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__o21a_1 _09612_ (.A1(_02860_),
    .A2(_02855_),
    .B1(_02854_),
    .X(_02865_));
 sky130_fd_sc_hd__nand2_1 _09613_ (.A(_02864_),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__a21bo_1 _09614_ (.A1(_02549_),
    .A2(_02569_),
    .B1_N(_02570_),
    .X(_02867_));
 sky130_fd_sc_hd__xor2_1 _09615_ (.A(_02566_),
    .B(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__mux2_1 _09616_ (.A0(_02558_),
    .A1(_02868_),
    .S(_02744_),
    .X(_02869_));
 sky130_fd_sc_hd__or2_1 _09617_ (.A(_00092_),
    .B(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__nand2_1 _09618_ (.A(_02575_),
    .B(_02594_),
    .Y(_02871_));
 sky130_fd_sc_hd__or2_1 _09619_ (.A(_02594_),
    .B(_02575_),
    .X(_02872_));
 sky130_fd_sc_hd__nor2_1 _09620_ (.A(_02580_),
    .B(_02767_),
    .Y(_02874_));
 sky130_fd_sc_hd__a31o_1 _09621_ (.A1(_02871_),
    .A2(_02767_),
    .A3(_02872_),
    .B1(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__or2_1 _09622_ (.A(_01240_),
    .B(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__buf_6 _09623_ (.A(_01240_),
    .X(_02877_));
 sky130_fd_sc_hd__nand2_1 _09624_ (.A(_02875_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _09625_ (.A(_02876_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__or2_1 _09626_ (.A(_02870_),
    .B(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(_02879_),
    .B(_02870_),
    .Y(_02881_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(_02880_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__inv_2 _09629_ (.A(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2_1 _09630_ (.A(_02869_),
    .B(_00092_),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_1 _09631_ (.A(_02870_),
    .B(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__or2_1 _09632_ (.A(_02842_),
    .B(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__nand2_1 _09633_ (.A(_02886_),
    .B(_02842_),
    .Y(_02888_));
 sky130_fd_sc_hd__nand2_1 _09634_ (.A(_02887_),
    .B(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__inv_2 _09635_ (.A(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__nand3_1 _09636_ (.A(_02866_),
    .B(_02883_),
    .C(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__o21a_1 _09637_ (.A1(_02888_),
    .A2(_02882_),
    .B1(_02881_),
    .X(_02892_));
 sky130_fd_sc_hd__nand2_1 _09638_ (.A(_02891_),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__nand2_1 _09639_ (.A(_02871_),
    .B(_02592_),
    .Y(_02894_));
 sky130_fd_sc_hd__or2_1 _09640_ (.A(_02588_),
    .B(_02894_),
    .X(_02896_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(_02894_),
    .B(_02588_),
    .Y(_02897_));
 sky130_fd_sc_hd__buf_6 _09642_ (.A(_02773_),
    .X(_02898_));
 sky130_fd_sc_hd__a21o_1 _09643_ (.A1(_02896_),
    .A2(_02897_),
    .B1(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__buf_6 _09644_ (.A(_02767_),
    .X(_02900_));
 sky130_fd_sc_hd__or2_1 _09645_ (.A(_02465_),
    .B(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__nand2_1 _09646_ (.A(_02899_),
    .B(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__inv_2 _09647_ (.A(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__nand2_1 _09648_ (.A(_02903_),
    .B(_01712_),
    .Y(_02904_));
 sky130_fd_sc_hd__nand2_1 _09649_ (.A(_02902_),
    .B(\sq.out[18] ),
    .Y(_02905_));
 sky130_fd_sc_hd__nand2_1 _09650_ (.A(_02904_),
    .B(_02905_),
    .Y(_02907_));
 sky130_fd_sc_hd__or2_1 _09651_ (.A(_02907_),
    .B(_02876_),
    .X(_02908_));
 sky130_fd_sc_hd__nand2_1 _09652_ (.A(_02876_),
    .B(_02907_),
    .Y(_02909_));
 sky130_fd_sc_hd__nand2_1 _09653_ (.A(_02908_),
    .B(_02909_),
    .Y(_02910_));
 sky130_fd_sc_hd__nand2b_1 _09654_ (.A_N(_02721_),
    .B(_02595_),
    .Y(_02911_));
 sky130_fd_sc_hd__or2b_1 _09655_ (.A(_02471_),
    .B_N(_02911_),
    .X(_02912_));
 sky130_fd_sc_hd__or2b_1 _09656_ (.A(_02911_),
    .B_N(_02471_),
    .X(_02913_));
 sky130_fd_sc_hd__nor2_1 _09657_ (.A(_02459_),
    .B(_02900_),
    .Y(_02914_));
 sky130_fd_sc_hd__a31o_1 _09658_ (.A1(_02900_),
    .A2(_02912_),
    .A3(_02913_),
    .B1(_02914_),
    .X(_02915_));
 sky130_fd_sc_hd__or2_1 _09659_ (.A(_05130_),
    .B(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__nand2_1 _09660_ (.A(_02915_),
    .B(_05140_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand2_1 _09661_ (.A(_02916_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__or2_1 _09662_ (.A(_02905_),
    .B(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__nand2_1 _09663_ (.A(_02919_),
    .B(_02905_),
    .Y(_02921_));
 sky130_fd_sc_hd__nand2_1 _09664_ (.A(_02920_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__nor2_1 _09665_ (.A(_02910_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__nand2_1 _09666_ (.A(_02893_),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__o21a_1 _09667_ (.A1(_02909_),
    .A2(_02922_),
    .B1(_02921_),
    .X(_02925_));
 sky130_fd_sc_hd__nand2_2 _09668_ (.A(_02924_),
    .B(_02925_),
    .Y(_02926_));
 sky130_fd_sc_hd__buf_6 _09669_ (.A(_00455_),
    .X(_02927_));
 sky130_fd_sc_hd__o21ai_2 _09670_ (.A1(_02490_),
    .A2(_02595_),
    .B1(_02723_),
    .Y(_02929_));
 sky130_fd_sc_hd__xor2_1 _09671_ (.A(_02705_),
    .B(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__or2_1 _09672_ (.A(_02692_),
    .B(_02767_),
    .X(_02931_));
 sky130_fd_sc_hd__o21ai_2 _09673_ (.A1(_02898_),
    .A2(_02930_),
    .B1(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__or2_1 _09674_ (.A(_02927_),
    .B(_02932_),
    .X(_02933_));
 sky130_fd_sc_hd__a21bo_1 _09675_ (.A1(_02929_),
    .A2(_02704_),
    .B1_N(_02703_),
    .X(_02934_));
 sky130_fd_sc_hd__xor2_1 _09676_ (.A(_02700_),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__nand2_1 _09677_ (.A(_02935_),
    .B(_02767_),
    .Y(_02936_));
 sky130_fd_sc_hd__or2_1 _09678_ (.A(_02694_),
    .B(_02744_),
    .X(_02937_));
 sky130_fd_sc_hd__nand2_1 _09679_ (.A(_02936_),
    .B(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__inv_2 _09680_ (.A(_02938_),
    .Y(_02940_));
 sky130_fd_sc_hd__nor2_1 _09681_ (.A(_02009_),
    .B(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__inv_2 _09682_ (.A(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2_1 _09683_ (.A(_02940_),
    .B(_02009_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand2_1 _09684_ (.A(_02942_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__or2_1 _09685_ (.A(_02933_),
    .B(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__nand2_1 _09686_ (.A(_02944_),
    .B(_02933_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand2_1 _09687_ (.A(_02945_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__inv_2 _09688_ (.A(_02947_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand2_1 _09689_ (.A(_02912_),
    .B(_02469_),
    .Y(_02949_));
 sky130_fd_sc_hd__xor2_1 _09690_ (.A(_02487_),
    .B(_02949_),
    .X(_02951_));
 sky130_fd_sc_hd__nand2_1 _09691_ (.A(_02951_),
    .B(_02900_),
    .Y(_02952_));
 sky130_fd_sc_hd__o21ai_2 _09692_ (.A1(_02481_),
    .A2(_02900_),
    .B1(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__nand2_1 _09693_ (.A(_02953_),
    .B(\sq.out[20] ),
    .Y(_02954_));
 sky130_fd_sc_hd__nand2_1 _09694_ (.A(_02932_),
    .B(_02927_),
    .Y(_02955_));
 sky130_fd_sc_hd__nand2_1 _09695_ (.A(_02933_),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hd__or2_1 _09696_ (.A(_02954_),
    .B(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__nand2_1 _09697_ (.A(_02956_),
    .B(_02954_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand2_1 _09698_ (.A(_02957_),
    .B(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__inv_2 _09699_ (.A(_02953_),
    .Y(_02960_));
 sky130_fd_sc_hd__nand2_1 _09700_ (.A(_02960_),
    .B(_01730_),
    .Y(_02962_));
 sky130_fd_sc_hd__nand2_1 _09701_ (.A(_02962_),
    .B(_02954_),
    .Y(_02963_));
 sky130_fd_sc_hd__or2_1 _09702_ (.A(_02916_),
    .B(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__nand2_1 _09703_ (.A(_02963_),
    .B(_02916_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_02964_),
    .B(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__nor2_1 _09705_ (.A(_02959_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__inv_2 _09706_ (.A(_02681_),
    .Y(_02968_));
 sky130_fd_sc_hd__a21o_1 _09707_ (.A1(_02929_),
    .A2(_02706_),
    .B1(_02715_),
    .X(_02969_));
 sky130_fd_sc_hd__or2_1 _09708_ (.A(_02968_),
    .B(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__nand2_1 _09709_ (.A(_02969_),
    .B(_02968_),
    .Y(_02971_));
 sky130_fd_sc_hd__nand3_1 _09710_ (.A(_02970_),
    .B(_02900_),
    .C(_02971_),
    .Y(_02973_));
 sky130_fd_sc_hd__or2_1 _09711_ (.A(_02670_),
    .B(_02900_),
    .X(_02974_));
 sky130_fd_sc_hd__nand2_2 _09712_ (.A(_02973_),
    .B(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__inv_2 _09713_ (.A(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__nand2_1 _09714_ (.A(_02976_),
    .B(\sq.out[23] ),
    .Y(_02977_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(_02975_),
    .B(_01993_),
    .Y(_02978_));
 sky130_fd_sc_hd__nand2_1 _09716_ (.A(_02977_),
    .B(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__nor2_1 _09717_ (.A(_02979_),
    .B(_02942_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand2_1 _09718_ (.A(_02942_),
    .B(_02979_),
    .Y(_02981_));
 sky130_fd_sc_hd__nor2b_1 _09719_ (.A(_02980_),
    .B_N(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__and3_1 _09720_ (.A(_02948_),
    .B(_02967_),
    .C(_02982_),
    .X(_02984_));
 sky130_fd_sc_hd__nand2_1 _09721_ (.A(_02926_),
    .B(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__o21a_1 _09722_ (.A1(_02965_),
    .A2(_02959_),
    .B1(_02958_),
    .X(_02986_));
 sky130_fd_sc_hd__nand2_1 _09723_ (.A(_02948_),
    .B(_02982_),
    .Y(_02987_));
 sky130_fd_sc_hd__o221a_1 _09724_ (.A1(_02980_),
    .A2(_02946_),
    .B1(_02986_),
    .B2(_02987_),
    .C1(_02981_),
    .X(_02988_));
 sky130_fd_sc_hd__nand2_2 _09725_ (.A(_02985_),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand2_1 _09726_ (.A(_02971_),
    .B(_02679_),
    .Y(_02990_));
 sky130_fd_sc_hd__xor2_1 _09727_ (.A(_02687_),
    .B(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _09728_ (.A0(_02991_),
    .A1(_02639_),
    .S(_02773_),
    .X(_02992_));
 sky130_fd_sc_hd__nand2_1 _09729_ (.A(_02992_),
    .B(_02071_),
    .Y(_02993_));
 sky130_fd_sc_hd__a21bo_1 _09730_ (.A1(_02596_),
    .A2(_02709_),
    .B1_N(_02725_),
    .X(_02995_));
 sky130_fd_sc_hd__xor2_1 _09731_ (.A(_02644_),
    .B(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__or2_1 _09732_ (.A(_02623_),
    .B(_02900_),
    .X(_02997_));
 sky130_fd_sc_hd__o21ai_2 _09733_ (.A1(_02898_),
    .A2(_02996_),
    .B1(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand2b_1 _09734_ (.A_N(_02993_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21o_1 _09735_ (.A1(_02992_),
    .A2(_02071_),
    .B1(_02998_),
    .X(_03000_));
 sky130_fd_sc_hd__nand2_1 _09736_ (.A(_02999_),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__or2_1 _09737_ (.A(_02071_),
    .B(_02992_),
    .X(_03002_));
 sky130_fd_sc_hd__nand2_1 _09738_ (.A(_03002_),
    .B(_02993_),
    .Y(_03003_));
 sky130_fd_sc_hd__or2_1 _09739_ (.A(_02977_),
    .B(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__nand2_1 _09740_ (.A(_03003_),
    .B(_02977_),
    .Y(_03006_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_03004_),
    .B(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__nor2_1 _09742_ (.A(_03001_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__inv_2 _09743_ (.A(_02658_),
    .Y(_03009_));
 sky130_fd_sc_hd__a21o_1 _09744_ (.A1(_02995_),
    .A2(_02645_),
    .B1(_02711_),
    .X(_03010_));
 sky130_fd_sc_hd__or2_1 _09745_ (.A(_03009_),
    .B(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__buf_6 _09746_ (.A(_02900_),
    .X(\sq.out[6] ));
 sky130_fd_sc_hd__nand2_1 _09747_ (.A(_03010_),
    .B(_03009_),
    .Y(_03012_));
 sky130_fd_sc_hd__nand3_1 _09748_ (.A(_03011_),
    .B(\sq.out[6] ),
    .C(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hd__nand2_1 _09749_ (.A(_02898_),
    .B(_02655_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_1 _09750_ (.A(_03013_),
    .B(_03014_),
    .Y(_03016_));
 sky130_fd_sc_hd__inv_2 _09751_ (.A(_02632_),
    .Y(_03017_));
 sky130_fd_sc_hd__a21bo_1 _09752_ (.A1(_02995_),
    .A2(_02643_),
    .B1_N(_02641_),
    .X(_03018_));
 sky130_fd_sc_hd__or2_1 _09753_ (.A(_03017_),
    .B(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__nand2_1 _09754_ (.A(_03018_),
    .B(_03017_),
    .Y(_03020_));
 sky130_fd_sc_hd__nor2_1 _09755_ (.A(_02627_),
    .B(_02900_),
    .Y(_03021_));
 sky130_fd_sc_hd__a31o_1 _09756_ (.A1(_03019_),
    .A2(\sq.out[6] ),
    .A3(_03020_),
    .B1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__or2_1 _09757_ (.A(_02998_),
    .B(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__nand2_1 _09758_ (.A(_03022_),
    .B(_02998_),
    .Y(_03024_));
 sky130_fd_sc_hd__nand2_1 _09759_ (.A(_03023_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nor2_1 _09760_ (.A(_03016_),
    .B(_03025_),
    .Y(_03027_));
 sky130_fd_sc_hd__and2_1 _09761_ (.A(_03008_),
    .B(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__nand2_2 _09762_ (.A(_02989_),
    .B(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__o21ai_1 _09763_ (.A1(_03001_),
    .A2(_03006_),
    .B1(_03000_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand2_1 _09764_ (.A(_03030_),
    .B(_03027_),
    .Y(_03031_));
 sky130_fd_sc_hd__and3_1 _09765_ (.A(_03024_),
    .B(_03013_),
    .C(_03014_),
    .X(_03032_));
 sky130_fd_sc_hd__nand2_1 _09766_ (.A(_03031_),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__nand2_1 _09767_ (.A(_02712_),
    .B(_02713_),
    .Y(_03034_));
 sky130_fd_sc_hd__a311o_1 _09768_ (.A1(_02995_),
    .A2(_02659_),
    .A3(_02645_),
    .B1(_03034_),
    .C1(_02773_),
    .X(_03035_));
 sky130_fd_sc_hd__or2_1 _09769_ (.A(_02604_),
    .B(_03035_),
    .X(_03036_));
 sky130_fd_sc_hd__nand2_1 _09770_ (.A(_03035_),
    .B(_02604_),
    .Y(_03038_));
 sky130_fd_sc_hd__nand2_1 _09771_ (.A(_03036_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__nand2_1 _09772_ (.A(_02597_),
    .B(_02444_),
    .Y(_03040_));
 sky130_fd_sc_hd__or2_1 _09773_ (.A(_02607_),
    .B(_03035_),
    .X(_03041_));
 sky130_fd_sc_hd__or2_1 _09774_ (.A(_03040_),
    .B(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__nand2_1 _09775_ (.A(_03041_),
    .B(_03040_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand2_1 _09776_ (.A(_03042_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__a21boi_1 _09777_ (.A1(_02606_),
    .A2(_03036_),
    .B1_N(_03041_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2b_1 _09778_ (.A_N(_03044_),
    .B(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hd__and3_1 _09779_ (.A(_03012_),
    .B(_02656_),
    .C(\sq.out[6] ),
    .X(_03047_));
 sky130_fd_sc_hd__xnor2_1 _09780_ (.A(_02648_),
    .B(_03047_),
    .Y(_03049_));
 sky130_fd_sc_hd__nor3b_1 _09781_ (.A(_03039_),
    .B(_03046_),
    .C_N(_03049_),
    .Y(_03050_));
 sky130_fd_sc_hd__nand2b_1 _09782_ (.A_N(_03033_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__clkinvlp_2 _09783_ (.A(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__nand2_1 _09784_ (.A(_02747_),
    .B(_02437_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2_1 _09785_ (.A(_02748_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__or2_1 _09786_ (.A(_02734_),
    .B(_02746_),
    .X(_03055_));
 sky130_fd_sc_hd__and2_1 _09787_ (.A(_03055_),
    .B(_02747_),
    .X(_03056_));
 sky130_fd_sc_hd__nand2_1 _09788_ (.A(_02745_),
    .B(_02451_),
    .Y(_03057_));
 sky130_fd_sc_hd__and2b_1 _09789_ (.A_N(_02746_),
    .B(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__nand2_1 _09790_ (.A(_03056_),
    .B(_03058_),
    .Y(_03060_));
 sky130_fd_sc_hd__or2_1 _09791_ (.A(_02266_),
    .B(_02446_),
    .X(_03061_));
 sky130_fd_sc_hd__nand2_1 _09792_ (.A(_03061_),
    .B(_02447_),
    .Y(_03062_));
 sky130_fd_sc_hd__xnor2_2 _09793_ (.A(_03062_),
    .B(_03042_),
    .Y(_03063_));
 sky130_fd_sc_hd__nor3_1 _09794_ (.A(_03054_),
    .B(_03060_),
    .C(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__nand3_4 _09795_ (.A(_03029_),
    .B(_03052_),
    .C(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__nor2_4 _09796_ (.A(_03065_),
    .B(_02764_),
    .Y(_03066_));
 sky130_fd_sc_hd__and3b_1 _09797_ (.A_N(_02745_),
    .B(_02739_),
    .C(_02738_),
    .X(_03067_));
 sky130_fd_sc_hd__o21ba_1 _09798_ (.A1(_02739_),
    .A2(_02760_),
    .B1_N(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__or2_1 _09799_ (.A(_02728_),
    .B(_03067_),
    .X(_03069_));
 sky130_fd_sc_hd__nand2_1 _09800_ (.A(_03067_),
    .B(_02728_),
    .Y(_03071_));
 sky130_fd_sc_hd__and2_1 _09801_ (.A(_03069_),
    .B(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__and2_1 _09802_ (.A(_03068_),
    .B(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__or3_1 _09803_ (.A(_01861_),
    .B(_01862_),
    .C(_02110_),
    .X(_03074_));
 sky130_fd_sc_hd__or2b_1 _09804_ (.A(_03071_),
    .B_N(_03074_),
    .X(_03075_));
 sky130_fd_sc_hd__a21o_1 _09805_ (.A1(_03067_),
    .A2(_02728_),
    .B1(_03074_),
    .X(_03076_));
 sky130_fd_sc_hd__nand2_1 _09806_ (.A(_03075_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__or3_1 _09807_ (.A(_01861_),
    .B(_01862_),
    .C(_02110_),
    .X(_03078_));
 sky130_fd_sc_hd__xor2_1 _09808_ (.A(_03078_),
    .B(_03075_),
    .X(_03079_));
 sky130_fd_sc_hd__or2_1 _09809_ (.A(_03077_),
    .B(_03079_),
    .X(_03080_));
 sky130_fd_sc_hd__inv_2 _09810_ (.A(_03080_),
    .Y(_03082_));
 sky130_fd_sc_hd__nand2_1 _09811_ (.A(_03073_),
    .B(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hd__clkinvlp_2 _09812_ (.A(_03083_),
    .Y(_03084_));
 sky130_fd_sc_hd__a31oi_2 _09813_ (.A1(_03067_),
    .A2(_02728_),
    .A3(_02729_),
    .B1(_02740_),
    .Y(_03085_));
 sky130_fd_sc_hd__or2_1 _09814_ (.A(_02410_),
    .B(_02417_),
    .X(_03086_));
 sky130_fd_sc_hd__o311ai_4 _09815_ (.A1(_01861_),
    .A2(_01862_),
    .A3(_02110_),
    .B1(_03086_),
    .C1(_03071_),
    .Y(_03087_));
 sky130_fd_sc_hd__or2_1 _09816_ (.A(_03085_),
    .B(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__inv_2 _09817_ (.A(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__nand3_4 _09818_ (.A(_03066_),
    .B(_03084_),
    .C(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__nand2_1 _09819_ (.A(_02808_),
    .B(_02834_),
    .Y(_03091_));
 sky130_fd_sc_hd__or2_1 _09820_ (.A(_02834_),
    .B(_02808_),
    .X(_03093_));
 sky130_fd_sc_hd__nand3_1 _09821_ (.A(net85),
    .B(_03091_),
    .C(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__inv_4 _09822_ (.A(_03090_),
    .Y(_03095_));
 sky130_fd_sc_hd__nand2_1 _09823_ (.A(_03095_),
    .B(_02820_),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _09824_ (.A(_03094_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__or2_1 _09825_ (.A(_00844_),
    .B(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__buf_6 _09826_ (.A(_03095_),
    .X(_03099_));
 sky130_fd_sc_hd__nand2_1 _09827_ (.A(_03091_),
    .B(_02831_),
    .Y(_03100_));
 sky130_fd_sc_hd__or2_1 _09828_ (.A(_02825_),
    .B(_03100_),
    .X(_03101_));
 sky130_fd_sc_hd__nand2_1 _09829_ (.A(_03100_),
    .B(_02825_),
    .Y(_03102_));
 sky130_fd_sc_hd__nand3_1 _09830_ (.A(net85),
    .B(_03101_),
    .C(_03102_),
    .Y(_03104_));
 sky130_fd_sc_hd__a21bo_1 _09831_ (.A1(_02813_),
    .A2(_03099_),
    .B1_N(_03104_),
    .X(_03105_));
 sky130_fd_sc_hd__or2_1 _09832_ (.A(_02856_),
    .B(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__nand2_1 _09833_ (.A(_03105_),
    .B(_02856_),
    .Y(_03107_));
 sky130_fd_sc_hd__nand2_1 _09834_ (.A(_03106_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__or2_1 _09835_ (.A(_03098_),
    .B(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__nand2_1 _09836_ (.A(_03108_),
    .B(_03098_),
    .Y(_03110_));
 sky130_fd_sc_hd__nand2_1 _09837_ (.A(_03109_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__buf_6 _09838_ (.A(_02441_),
    .X(_03112_));
 sky130_fd_sc_hd__nor3_4 _09839_ (.A(_02764_),
    .B(_03083_),
    .C(_03065_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand3_2 _09840_ (.A(_03113_),
    .B(_02898_),
    .C(_03089_),
    .Y(_03115_));
 sky130_fd_sc_hd__nor3_1 _09841_ (.A(\sq.out[8] ),
    .B(_03112_),
    .C(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__buf_6 _09842_ (.A(_03090_),
    .X(_03117_));
 sky130_fd_sc_hd__xor2_1 _09843_ (.A(\sq.out[7] ),
    .B(\sq.out[6] ),
    .X(_03118_));
 sky130_fd_sc_hd__a21oi_1 _09844_ (.A1(_03117_),
    .A2(_03112_),
    .B1(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__nand2_1 _09845_ (.A(_03117_),
    .B(_03118_),
    .Y(_03120_));
 sky130_fd_sc_hd__nand2_1 _09846_ (.A(_03115_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__nand2_1 _09847_ (.A(_03121_),
    .B(\sq.out[8] ),
    .Y(_03122_));
 sky130_fd_sc_hd__nand3_1 _09848_ (.A(_03115_),
    .B(_03120_),
    .C(_02498_),
    .Y(_03123_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_03122_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__nor2_2 _09850_ (.A(\sq.out[6] ),
    .B(_03090_),
    .Y(_03126_));
 sky130_fd_sc_hd__nand2_1 _09851_ (.A(_03126_),
    .B(\sq.out[7] ),
    .Y(_03127_));
 sky130_fd_sc_hd__nand2_1 _09852_ (.A(_03124_),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__o21ai_1 _09853_ (.A1(_03116_),
    .A2(_03119_),
    .B1(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_1 _09854_ (.A(_03126_),
    .B(_03112_),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_1 _09855_ (.A(net85),
    .B(_02778_),
    .Y(_03131_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(_03130_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__nand2_1 _09857_ (.A(_03132_),
    .B(\sq.out[9] ),
    .Y(_03133_));
 sky130_fd_sc_hd__nand3_1 _09858_ (.A(_03130_),
    .B(_02495_),
    .C(_03131_),
    .Y(_03134_));
 sky130_fd_sc_hd__nand2_1 _09859_ (.A(_03133_),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(_03135_),
    .B(_03122_),
    .Y(_03137_));
 sky130_fd_sc_hd__nand3b_1 _09861_ (.A_N(_03122_),
    .B(_03133_),
    .C(_03134_),
    .Y(_03138_));
 sky130_fd_sc_hd__nand3_1 _09862_ (.A(_03129_),
    .B(_03137_),
    .C(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__nand2_1 _09863_ (.A(_03139_),
    .B(_03137_),
    .Y(_03140_));
 sky130_fd_sc_hd__or2_1 _09864_ (.A(_02769_),
    .B(_03090_),
    .X(_03141_));
 sky130_fd_sc_hd__a21o_1 _09865_ (.A1(_02782_),
    .A2(_02784_),
    .B1(_02788_),
    .X(_03142_));
 sky130_fd_sc_hd__nand3_1 _09866_ (.A(net85),
    .B(_02789_),
    .C(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2_1 _09867_ (.A(_03141_),
    .B(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__nand2_1 _09868_ (.A(_03144_),
    .B(_02345_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand3_2 _09869_ (.A(_03141_),
    .B(\sq.out[11] ),
    .C(_03143_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand2_1 _09870_ (.A(_03145_),
    .B(_03146_),
    .Y(_03148_));
 sky130_fd_sc_hd__inv_2 _09871_ (.A(_02788_),
    .Y(_03149_));
 sky130_fd_sc_hd__a21boi_1 _09872_ (.A1(_02781_),
    .A2(_02787_),
    .B1_N(_02786_),
    .Y(_03150_));
 sky130_fd_sc_hd__o21ai_1 _09873_ (.A1(_03149_),
    .A2(_03150_),
    .B1(_03090_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand3b_1 _09874_ (.A_N(_02780_),
    .B(_03113_),
    .C(_03089_),
    .Y(_03152_));
 sky130_fd_sc_hd__nand3_1 _09875_ (.A(_03151_),
    .B(_03152_),
    .C(\sq.out[10] ),
    .Y(_03153_));
 sky130_fd_sc_hd__nand2_1 _09876_ (.A(_03148_),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__nand3b_1 _09877_ (.A_N(_03153_),
    .B(_03145_),
    .C(_03146_),
    .Y(_03155_));
 sky130_fd_sc_hd__nand2_1 _09878_ (.A(_03154_),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__inv_2 _09879_ (.A(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__nand2_1 _09880_ (.A(_03151_),
    .B(_03152_),
    .Y(_03159_));
 sky130_fd_sc_hd__nand2_1 _09881_ (.A(_03159_),
    .B(_02504_),
    .Y(_03160_));
 sky130_fd_sc_hd__nand2_1 _09882_ (.A(_03160_),
    .B(_03153_),
    .Y(_03161_));
 sky130_fd_sc_hd__or2_1 _09883_ (.A(_03133_),
    .B(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(_03161_),
    .B(_03133_),
    .Y(_03163_));
 sky130_fd_sc_hd__and2_1 _09885_ (.A(_03162_),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__nand3_1 _09886_ (.A(_03140_),
    .B(_03157_),
    .C(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__o21a_1 _09887_ (.A1(_03163_),
    .A2(_03156_),
    .B1(_03154_),
    .X(_03166_));
 sky130_fd_sc_hd__nand2_2 _09888_ (.A(_03165_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand2_1 _09889_ (.A(_02789_),
    .B(_02782_),
    .Y(_03168_));
 sky130_fd_sc_hd__or2_1 _09890_ (.A(_02804_),
    .B(_03168_),
    .X(_03170_));
 sky130_fd_sc_hd__nand2_1 _09891_ (.A(_03168_),
    .B(_02804_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _09892_ (.A(_03170_),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand2_1 _09893_ (.A(_03099_),
    .B(_02798_),
    .Y(_03173_));
 sky130_fd_sc_hd__o21ai_2 _09894_ (.A1(_03172_),
    .A2(_03099_),
    .B1(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__or2_1 _09895_ (.A(_02826_),
    .B(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__nand2_1 _09896_ (.A(_03097_),
    .B(_00844_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand2_1 _09897_ (.A(_03098_),
    .B(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__or2_1 _09898_ (.A(_03175_),
    .B(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__nand2_1 _09899_ (.A(_03177_),
    .B(_03175_),
    .Y(_03179_));
 sky130_fd_sc_hd__nand2_1 _09900_ (.A(_03178_),
    .B(_03179_),
    .Y(_03181_));
 sky130_fd_sc_hd__nand2_1 _09901_ (.A(_03174_),
    .B(_02826_),
    .Y(_03182_));
 sky130_fd_sc_hd__nand2_1 _09902_ (.A(_03175_),
    .B(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__or2_1 _09903_ (.A(_03146_),
    .B(_03183_),
    .X(_03184_));
 sky130_fd_sc_hd__nand2_1 _09904_ (.A(_03183_),
    .B(_03146_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_1 _09905_ (.A(_03184_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__nor2_1 _09906_ (.A(_03181_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_1 _09907_ (.A(_03167_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__o21a_1 _09908_ (.A1(_03185_),
    .A2(_03181_),
    .B1(_03179_),
    .X(_03189_));
 sky130_fd_sc_hd__nand2_1 _09909_ (.A(_03188_),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__xor2_1 _09910_ (.A(_03111_),
    .B(_03190_),
    .X(_03192_));
 sky130_fd_sc_hd__buf_6 _09911_ (.A(_03117_),
    .X(\sq.out[5] ));
 sky130_fd_sc_hd__nand2_1 _09912_ (.A(\sq.out[5] ),
    .B(_03066_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand2b_1 _09913_ (.A_N(_03193_),
    .B(_03073_),
    .Y(_03194_));
 sky130_fd_sc_hd__o21ai_1 _09914_ (.A1(_03077_),
    .A2(_03194_),
    .B1(_03079_),
    .Y(_03195_));
 sky130_fd_sc_hd__nand2_1 _09915_ (.A(_03113_),
    .B(_03088_),
    .Y(_03196_));
 sky130_fd_sc_hd__or2_1 _09916_ (.A(_03087_),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__nand2_1 _09917_ (.A(_03196_),
    .B(_03087_),
    .Y(_03198_));
 sky130_fd_sc_hd__and2_1 _09918_ (.A(_03197_),
    .B(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__and3_1 _09919_ (.A(_03195_),
    .B(_03196_),
    .C(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__nand2_1 _09920_ (.A(_03197_),
    .B(_03085_),
    .Y(_03202_));
 sky130_fd_sc_hd__nand2_1 _09921_ (.A(_03200_),
    .B(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__buf_8 _09922_ (.A(_03099_),
    .X(_03204_));
 sky130_fd_sc_hd__or2_1 _09923_ (.A(_03065_),
    .B(_03204_),
    .X(_03205_));
 sky130_fd_sc_hd__or2_1 _09924_ (.A(_02756_),
    .B(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__or2_1 _09925_ (.A(_02758_),
    .B(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__or2_1 _09926_ (.A(_02754_),
    .B(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__xor2_2 _09927_ (.A(_02762_),
    .B(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__xor2_1 _09928_ (.A(_03068_),
    .B(_03193_),
    .X(_03210_));
 sky130_fd_sc_hd__a21o_1 _09929_ (.A1(_03066_),
    .A2(_03068_),
    .B1(_03072_),
    .X(_03211_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(_03194_),
    .B(_03211_),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_1 _09931_ (.A(_03077_),
    .B(_03194_),
    .Y(_03214_));
 sky130_fd_sc_hd__nor3_1 _09932_ (.A(_03210_),
    .B(_03213_),
    .C(_03214_),
    .Y(_03215_));
 sky130_fd_sc_hd__nand2_1 _09933_ (.A(_03209_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__nor2_2 _09934_ (.A(_03203_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__inv_2 _09935_ (.A(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__or2b_1 _09936_ (.A(_02837_),
    .B_N(_02861_),
    .X(_03219_));
 sky130_fd_sc_hd__a21o_1 _09937_ (.A1(_02835_),
    .A2(_02836_),
    .B1(_02861_),
    .X(_03220_));
 sky130_fd_sc_hd__nand2_1 _09938_ (.A(_03219_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__nand2_1 _09939_ (.A(_03099_),
    .B(_02850_),
    .Y(_03222_));
 sky130_fd_sc_hd__o21ai_2 _09940_ (.A1(_03221_),
    .A2(_03099_),
    .B1(_03222_),
    .Y(_03224_));
 sky130_fd_sc_hd__or2_1 _09941_ (.A(_02843_),
    .B(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__nand2_1 _09942_ (.A(_03224_),
    .B(_02843_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand2_1 _09943_ (.A(_03225_),
    .B(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__or2_1 _09944_ (.A(_03227_),
    .B(_03106_),
    .X(_03228_));
 sky130_fd_sc_hd__nand2_1 _09945_ (.A(_03106_),
    .B(_03227_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _09946_ (.A(_03228_),
    .B(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__nor2_1 _09947_ (.A(_03230_),
    .B(_03111_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _09948_ (.A(_03190_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__o21a_1 _09949_ (.A1(_03110_),
    .A2(_03230_),
    .B1(_03229_),
    .X(_03233_));
 sky130_fd_sc_hd__nand2_1 _09950_ (.A(_03232_),
    .B(_03233_),
    .Y(_03235_));
 sky130_fd_sc_hd__nand2_1 _09951_ (.A(_02866_),
    .B(_02890_),
    .Y(_03236_));
 sky130_fd_sc_hd__or2_1 _09952_ (.A(_02890_),
    .B(_02866_),
    .X(_03237_));
 sky130_fd_sc_hd__nand3_1 _09953_ (.A(_03117_),
    .B(_03236_),
    .C(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand2_1 _09954_ (.A(_03099_),
    .B(_02869_),
    .Y(_03239_));
 sky130_fd_sc_hd__nand2_1 _09955_ (.A(_03238_),
    .B(_03239_),
    .Y(_03240_));
 sky130_fd_sc_hd__inv_2 _09956_ (.A(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _09957_ (.A(_03241_),
    .B(\sq.out[17] ),
    .Y(_03242_));
 sky130_fd_sc_hd__nand2_1 _09958_ (.A(_03240_),
    .B(_02877_),
    .Y(_03243_));
 sky130_fd_sc_hd__nand2_1 _09959_ (.A(_03242_),
    .B(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand2_1 _09960_ (.A(_03220_),
    .B(_02860_),
    .Y(_03246_));
 sky130_fd_sc_hd__xor2_1 _09961_ (.A(_02855_),
    .B(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(_03204_),
    .B(_02841_),
    .Y(_03248_));
 sky130_fd_sc_hd__o21ai_2 _09963_ (.A1(_03247_),
    .A2(_03204_),
    .B1(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hd__or2_1 _09964_ (.A(_00092_),
    .B(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__or2_1 _09965_ (.A(_03244_),
    .B(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__nand2_1 _09966_ (.A(_03250_),
    .B(_03244_),
    .Y(_03252_));
 sky130_fd_sc_hd__nand2_1 _09967_ (.A(_03251_),
    .B(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__inv_2 _09968_ (.A(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand2_1 _09969_ (.A(_03249_),
    .B(_00092_),
    .Y(_03255_));
 sky130_fd_sc_hd__nand2_1 _09970_ (.A(_03250_),
    .B(_03255_),
    .Y(_03257_));
 sky130_fd_sc_hd__or2_1 _09971_ (.A(_03225_),
    .B(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__nand2_1 _09972_ (.A(_03257_),
    .B(_03225_),
    .Y(_03259_));
 sky130_fd_sc_hd__nand2_1 _09973_ (.A(_03258_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__inv_2 _09974_ (.A(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand3_1 _09975_ (.A(_03235_),
    .B(_03254_),
    .C(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__inv_2 _09976_ (.A(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__a21bo_1 _09977_ (.A1(_02926_),
    .A2(_02964_),
    .B1_N(_02965_),
    .X(_03264_));
 sky130_fd_sc_hd__xor2_1 _09978_ (.A(_02959_),
    .B(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__nand2_1 _09979_ (.A(_03117_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__o21ai_1 _09980_ (.A1(_02932_),
    .A2(_03117_),
    .B1(_03266_),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_1 _09981_ (.A(_03268_),
    .B(\sq.out[22] ),
    .Y(_03269_));
 sky130_fd_sc_hd__a21bo_1 _09982_ (.A1(_02926_),
    .A2(_02967_),
    .B1_N(_02986_),
    .X(_03270_));
 sky130_fd_sc_hd__nand2_1 _09983_ (.A(_03270_),
    .B(_02948_),
    .Y(_03271_));
 sky130_fd_sc_hd__or2_1 _09984_ (.A(_02948_),
    .B(_03270_),
    .X(_03272_));
 sky130_fd_sc_hd__nand3_1 _09985_ (.A(_03117_),
    .B(_03271_),
    .C(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__nand2_1 _09986_ (.A(_03099_),
    .B(_02940_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_1 _09987_ (.A(_03273_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__inv_2 _09988_ (.A(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_1 _09989_ (.A(_03276_),
    .B(\sq.out[23] ),
    .Y(_03277_));
 sky130_fd_sc_hd__nand2_1 _09990_ (.A(_03275_),
    .B(_01993_),
    .Y(_03279_));
 sky130_fd_sc_hd__nand2_1 _09991_ (.A(_03277_),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__or2_1 _09992_ (.A(_03269_),
    .B(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__nand2_1 _09993_ (.A(_03280_),
    .B(_03269_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_1 _09994_ (.A(_03281_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__inv_2 _09995_ (.A(_03268_),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_03284_),
    .B(_02009_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _09997_ (.A(_03285_),
    .B(_03269_),
    .Y(_03286_));
 sky130_fd_sc_hd__xor2_1 _09998_ (.A(_02966_),
    .B(_02926_),
    .X(_03287_));
 sky130_fd_sc_hd__or2_1 _09999_ (.A(_03287_),
    .B(_03095_),
    .X(_03288_));
 sky130_fd_sc_hd__nand2_1 _10000_ (.A(_03099_),
    .B(_02960_),
    .Y(_03290_));
 sky130_fd_sc_hd__nand2_1 _10001_ (.A(_03288_),
    .B(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__inv_2 _10002_ (.A(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__nand2_1 _10003_ (.A(_03292_),
    .B(\sq.out[21] ),
    .Y(_03293_));
 sky130_fd_sc_hd__or2_1 _10004_ (.A(_03286_),
    .B(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__nand2_1 _10005_ (.A(_03293_),
    .B(_03286_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand2_1 _10006_ (.A(_03294_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__or2_1 _10007_ (.A(_03283_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__xor2_1 _10008_ (.A(_02910_),
    .B(_02893_),
    .X(_03298_));
 sky130_fd_sc_hd__or2_1 _10009_ (.A(_03298_),
    .B(_03099_),
    .X(_03299_));
 sky130_fd_sc_hd__nand2_1 _10010_ (.A(_03204_),
    .B(_02903_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand2_1 _10011_ (.A(_03299_),
    .B(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand2b_1 _10012_ (.A_N(_03302_),
    .B(\sq.out[19] ),
    .Y(_03303_));
 sky130_fd_sc_hd__a21bo_1 _10013_ (.A1(_02893_),
    .A2(_02908_),
    .B1_N(_02909_),
    .X(_03304_));
 sky130_fd_sc_hd__xnor2_1 _10014_ (.A(_02922_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(_02915_),
    .A1(_03305_),
    .S(net85),
    .X(_03306_));
 sky130_fd_sc_hd__or2_1 _10016_ (.A(_01730_),
    .B(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__nand2_1 _10017_ (.A(_03306_),
    .B(_01730_),
    .Y(_03308_));
 sky130_fd_sc_hd__nand2_1 _10018_ (.A(_03307_),
    .B(_03308_),
    .Y(_03309_));
 sky130_fd_sc_hd__or2_1 _10019_ (.A(_03303_),
    .B(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__nand2_1 _10020_ (.A(_03309_),
    .B(_03303_),
    .Y(_03312_));
 sky130_fd_sc_hd__nand2_1 _10021_ (.A(_03310_),
    .B(_03312_),
    .Y(_03313_));
 sky130_fd_sc_hd__inv_2 _10022_ (.A(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__nand2_1 _10023_ (.A(_03291_),
    .B(_02927_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand2_1 _10024_ (.A(_03293_),
    .B(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__or2_1 _10025_ (.A(_03316_),
    .B(_03307_),
    .X(_03317_));
 sky130_fd_sc_hd__nand2_1 _10026_ (.A(_03307_),
    .B(_03316_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2_1 _10027_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__inv_2 _10028_ (.A(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__nand2_1 _10029_ (.A(_03314_),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__nor2_1 _10030_ (.A(_03297_),
    .B(_03321_),
    .Y(_03323_));
 sky130_fd_sc_hd__nand2_1 _10031_ (.A(_03236_),
    .B(_02888_),
    .Y(_03324_));
 sky130_fd_sc_hd__or2_1 _10032_ (.A(_02883_),
    .B(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__nand2_1 _10033_ (.A(_03324_),
    .B(_02883_),
    .Y(_03326_));
 sky130_fd_sc_hd__nand2_1 _10034_ (.A(_03325_),
    .B(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__nand2_1 _10035_ (.A(_03204_),
    .B(_02875_),
    .Y(_03328_));
 sky130_fd_sc_hd__o21ai_1 _10036_ (.A1(_03327_),
    .A2(_03204_),
    .B1(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__or2_1 _10037_ (.A(_01712_),
    .B(_03329_),
    .X(_03330_));
 sky130_fd_sc_hd__nand2_1 _10038_ (.A(_03329_),
    .B(_01712_),
    .Y(_03331_));
 sky130_fd_sc_hd__nand2_1 _10039_ (.A(_03330_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__or2_1 _10040_ (.A(_03242_),
    .B(_03332_),
    .X(_03334_));
 sky130_fd_sc_hd__nand2_1 _10041_ (.A(_03332_),
    .B(_03242_),
    .Y(_03335_));
 sky130_fd_sc_hd__nand2_1 _10042_ (.A(_03334_),
    .B(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_1 _10043_ (.A(_03302_),
    .B(_05140_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand2_1 _10044_ (.A(_03303_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__or2_1 _10045_ (.A(_03330_),
    .B(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__nand2_1 _10046_ (.A(_03338_),
    .B(_03330_),
    .Y(_03340_));
 sky130_fd_sc_hd__nand2_1 _10047_ (.A(_03339_),
    .B(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__nor2_1 _10048_ (.A(_03336_),
    .B(_03341_),
    .Y(_03342_));
 sky130_fd_sc_hd__nand3_1 _10049_ (.A(_03263_),
    .B(_03323_),
    .C(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__o21a_1 _10050_ (.A1(_03312_),
    .A2(_03319_),
    .B1(_03318_),
    .X(_03345_));
 sky130_fd_sc_hd__o21a_1 _10051_ (.A1(_03295_),
    .A2(_03283_),
    .B1(_03282_),
    .X(_03346_));
 sky130_fd_sc_hd__o21ai_1 _10052_ (.A1(_03259_),
    .A2(_03253_),
    .B1(_03252_),
    .Y(_03347_));
 sky130_fd_sc_hd__o21ai_1 _10053_ (.A1(_03335_),
    .A2(_03341_),
    .B1(_03340_),
    .Y(_03348_));
 sky130_fd_sc_hd__a21o_1 _10054_ (.A1(_03347_),
    .A2(_03342_),
    .B1(_03348_),
    .X(_03349_));
 sky130_fd_sc_hd__nand2_1 _10055_ (.A(_03349_),
    .B(_03323_),
    .Y(_03350_));
 sky130_fd_sc_hd__o211a_1 _10056_ (.A1(_03297_),
    .A2(_03345_),
    .B1(_03346_),
    .C1(_03350_),
    .X(_03351_));
 sky130_fd_sc_hd__nand2_4 _10057_ (.A(_03343_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand2_1 _10058_ (.A(_03271_),
    .B(_02946_),
    .Y(_03353_));
 sky130_fd_sc_hd__or2_1 _10059_ (.A(_02982_),
    .B(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__nand2_1 _10060_ (.A(_03353_),
    .B(_02982_),
    .Y(_03356_));
 sky130_fd_sc_hd__a21o_1 _10061_ (.A1(_03354_),
    .A2(_03356_),
    .B1(_03204_),
    .X(_03357_));
 sky130_fd_sc_hd__o21ai_2 _10062_ (.A1(_02975_),
    .A2(_03117_),
    .B1(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__xor2_1 _10063_ (.A(_03007_),
    .B(_02989_),
    .X(_03359_));
 sky130_fd_sc_hd__or2_1 _10064_ (.A(_02992_),
    .B(_03117_),
    .X(_03360_));
 sky130_fd_sc_hd__o21ai_2 _10065_ (.A1(_03204_),
    .A2(_03359_),
    .B1(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__and3_1 _10066_ (.A(_03358_),
    .B(_03361_),
    .C(_02071_),
    .X(_03362_));
 sky130_fd_sc_hd__buf_6 _10067_ (.A(_02071_),
    .X(\sq.out[24] ));
 sky130_fd_sc_hd__a21o_1 _10068_ (.A1(_03358_),
    .A2(\sq.out[24] ),
    .B1(_03361_),
    .X(_03363_));
 sky130_fd_sc_hd__or2b_1 _10069_ (.A(_03362_),
    .B_N(_03363_),
    .X(_03364_));
 sky130_fd_sc_hd__xor2_1 _10070_ (.A(_01081_),
    .B(_03358_),
    .X(_03366_));
 sky130_fd_sc_hd__or2_1 _10071_ (.A(_03277_),
    .B(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__nand2_1 _10072_ (.A(_03366_),
    .B(_03277_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _10073_ (.A(_03367_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__nor2_1 _10074_ (.A(_03364_),
    .B(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__a21bo_1 _10075_ (.A1(_02989_),
    .A2(_03004_),
    .B1_N(_03006_),
    .X(_03371_));
 sky130_fd_sc_hd__xor2_1 _10076_ (.A(_03001_),
    .B(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__buf_6 _10077_ (.A(_03204_),
    .X(_03373_));
 sky130_fd_sc_hd__nand2_1 _10078_ (.A(_03373_),
    .B(_02998_),
    .Y(_03374_));
 sky130_fd_sc_hd__o21ai_1 _10079_ (.A1(_03372_),
    .A2(_03373_),
    .B1(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__nor2_1 _10080_ (.A(_03375_),
    .B(_03361_),
    .Y(_03377_));
 sky130_fd_sc_hd__nand2_1 _10081_ (.A(_03361_),
    .B(_03375_),
    .Y(_03378_));
 sky130_fd_sc_hd__inv_2 _10082_ (.A(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__nor2_1 _10083_ (.A(_03377_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__a21o_1 _10084_ (.A1(_02989_),
    .A2(_03008_),
    .B1(_03030_),
    .X(_03381_));
 sky130_fd_sc_hd__or2b_1 _10085_ (.A(_03025_),
    .B_N(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__or2b_1 _10086_ (.A(_03381_),
    .B_N(_03025_),
    .X(_03383_));
 sky130_fd_sc_hd__and2_1 _10087_ (.A(_03373_),
    .B(_03022_),
    .X(_03384_));
 sky130_fd_sc_hd__a31o_1 _10088_ (.A1(\sq.out[5] ),
    .A2(_03382_),
    .A3(_03383_),
    .B1(_03384_),
    .X(_03385_));
 sky130_fd_sc_hd__clkinvlp_2 _10089_ (.A(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__and3_1 _10090_ (.A(_03370_),
    .B(_03380_),
    .C(_03386_),
    .X(_03388_));
 sky130_fd_sc_hd__nand2_4 _10091_ (.A(_03352_),
    .B(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__o21a_1 _10092_ (.A1(_03362_),
    .A2(_03368_),
    .B1(_03363_),
    .X(_03390_));
 sky130_fd_sc_hd__o211a_1 _10093_ (.A1(_03377_),
    .A2(_03390_),
    .B1(_03378_),
    .C1(_03386_),
    .X(_03391_));
 sky130_fd_sc_hd__and3_1 _10094_ (.A(_03029_),
    .B(_03031_),
    .C(_03032_),
    .X(_03392_));
 sky130_fd_sc_hd__nand3_1 _10095_ (.A(_03117_),
    .B(_03049_),
    .C(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nor2_1 _10096_ (.A(_03039_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hd__or2_1 _10097_ (.A(_03045_),
    .B(_03394_),
    .X(_03395_));
 sky130_fd_sc_hd__nand2_1 _10098_ (.A(_03394_),
    .B(_03045_),
    .Y(_03396_));
 sky130_fd_sc_hd__and2_1 _10099_ (.A(_03395_),
    .B(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__nand2_1 _10100_ (.A(_03393_),
    .B(_03039_),
    .Y(_03399_));
 sky130_fd_sc_hd__and2b_1 _10101_ (.A_N(_03394_),
    .B(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__nand3_1 _10102_ (.A(\sq.out[5] ),
    .B(_03024_),
    .C(_03382_),
    .Y(_03401_));
 sky130_fd_sc_hd__xor2_1 _10103_ (.A(_03016_),
    .B(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__a21o_1 _10104_ (.A1(\sq.out[5] ),
    .A2(_03392_),
    .B1(_03049_),
    .X(_03403_));
 sky130_fd_sc_hd__nand2_1 _10105_ (.A(_03403_),
    .B(_03393_),
    .Y(_03404_));
 sky130_fd_sc_hd__inv_2 _10106_ (.A(_03404_),
    .Y(_03405_));
 sky130_fd_sc_hd__and4_1 _10107_ (.A(_03397_),
    .B(_03400_),
    .C(_03402_),
    .D(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__nand2_1 _10108_ (.A(_03391_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__inv_2 _10109_ (.A(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__or3b_1 _10110_ (.A(_03051_),
    .B(_03204_),
    .C_N(_03029_),
    .X(_03410_));
 sky130_fd_sc_hd__nor2_1 _10111_ (.A(_03063_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__and2_1 _10112_ (.A(_03411_),
    .B(_03058_),
    .X(_03412_));
 sky130_fd_sc_hd__nand2_1 _10113_ (.A(_03412_),
    .B(_03056_),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_2 _10114_ (.A(_03054_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand2_1 _10115_ (.A(_03205_),
    .B(_02756_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_1 _10116_ (.A(_03206_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_1 _10117_ (.A(_03206_),
    .B(_02758_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _10118_ (.A(_03207_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__nand2_1 _10119_ (.A(_03207_),
    .B(_02754_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_1 _10120_ (.A(_03208_),
    .B(_03419_),
    .Y(_03421_));
 sky130_fd_sc_hd__or3_1 _10121_ (.A(_03416_),
    .B(_03418_),
    .C(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__xor2_1 _10122_ (.A(_03044_),
    .B(_03396_),
    .X(_03423_));
 sky130_fd_sc_hd__inv_2 _10123_ (.A(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__nor2_1 _10124_ (.A(_03058_),
    .B(_03411_),
    .Y(_03425_));
 sky130_fd_sc_hd__nor2_1 _10125_ (.A(_03425_),
    .B(_03412_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _10126_ (.A(_03410_),
    .B(_03063_),
    .Y(_03427_));
 sky130_fd_sc_hd__and2b_1 _10127_ (.A_N(_03411_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__nand2_1 _10128_ (.A(_03426_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__or2_1 _10129_ (.A(_03056_),
    .B(_03412_),
    .X(_03430_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(_03430_),
    .B(_03413_),
    .Y(_03432_));
 sky130_fd_sc_hd__or3_1 _10131_ (.A(_03424_),
    .B(_03429_),
    .C(_03432_),
    .X(_03433_));
 sky130_fd_sc_hd__nor3_2 _10132_ (.A(_03414_),
    .B(_03422_),
    .C(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand3_4 _10133_ (.A(_03389_),
    .B(_03408_),
    .C(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__nor2_8 _10134_ (.A(_03218_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__buf_6 _10135_ (.A(_03436_),
    .X(_03437_));
 sky130_fd_sc_hd__buf_6 _10136_ (.A(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__buf_8 _10137_ (.A(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__nand2_1 _10138_ (.A(_03438_),
    .B(_03105_),
    .Y(_03440_));
 sky130_fd_sc_hd__o21ai_1 _10139_ (.A1(_03192_),
    .A2(_03439_),
    .B1(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__or2_4 _10140_ (.A(_02843_),
    .B(_03441_),
    .X(_03443_));
 sky130_fd_sc_hd__nand2_1 _10141_ (.A(_03441_),
    .B(_02843_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _10142_ (.A(_03443_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__a21bo_1 _10143_ (.A1(_03167_),
    .A2(_03184_),
    .B1_N(_03185_),
    .X(_03446_));
 sky130_fd_sc_hd__xor2_1 _10144_ (.A(_03181_),
    .B(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__nand2_1 _10145_ (.A(net97),
    .B(_03097_),
    .Y(_03448_));
 sky130_fd_sc_hd__o21ai_2 _10146_ (.A1(_03447_),
    .A2(net97),
    .B1(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__nor2_1 _10147_ (.A(_02856_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__inv_2 _10148_ (.A(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2_1 _10149_ (.A(_03445_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__nand3_1 _10150_ (.A(_03443_),
    .B(_03450_),
    .C(_03444_),
    .Y(_03454_));
 sky130_fd_sc_hd__nand2_1 _10151_ (.A(_03452_),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__o21bai_1 _10152_ (.A1(_03218_),
    .A2(_03435_),
    .B1_N(_03118_),
    .Y(_03456_));
 sky130_fd_sc_hd__nand2_1 _10153_ (.A(_03437_),
    .B(_03115_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_1 _10154_ (.A(_03456_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_03458_),
    .B(_02498_),
    .Y(_03459_));
 sky130_fd_sc_hd__nand3_1 _10156_ (.A(_03456_),
    .B(_03457_),
    .C(\sq.out[8] ),
    .Y(_03460_));
 sky130_fd_sc_hd__nand2_1 _10157_ (.A(_03459_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__nand2_1 _10158_ (.A(_03373_),
    .B(\sq.out[6] ),
    .Y(_03462_));
 sky130_fd_sc_hd__nand2_1 _10159_ (.A(\sq.out[5] ),
    .B(_02898_),
    .Y(_03463_));
 sky130_fd_sc_hd__nand2_1 _10160_ (.A(_03462_),
    .B(_03463_),
    .Y(_03465_));
 sky130_fd_sc_hd__o21bai_1 _10161_ (.A1(_03218_),
    .A2(_03435_),
    .B1_N(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__inv_2 _10162_ (.A(_03435_),
    .Y(_03467_));
 sky130_fd_sc_hd__nand3_1 _10163_ (.A(_03467_),
    .B(\sq.out[5] ),
    .C(_03217_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand3_1 _10164_ (.A(_03466_),
    .B(_03468_),
    .C(\sq.out[7] ),
    .Y(_03469_));
 sky130_fd_sc_hd__nand2_1 _10165_ (.A(_03461_),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_1 _10166_ (.A(_03466_),
    .B(_03468_),
    .Y(_03471_));
 sky130_fd_sc_hd__nor2_1 _10167_ (.A(_03112_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand3_1 _10168_ (.A(_03472_),
    .B(_03459_),
    .C(_03460_),
    .Y(_03473_));
 sky130_fd_sc_hd__nand2_1 _10169_ (.A(_03471_),
    .B(_03112_),
    .Y(_03474_));
 sky130_fd_sc_hd__inv_2 _10170_ (.A(_03463_),
    .Y(_03476_));
 sky130_fd_sc_hd__nor2_1 _10171_ (.A(\sq.out[5] ),
    .B(_03438_),
    .Y(_03477_));
 sky130_fd_sc_hd__nor2_1 _10172_ (.A(_03476_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__nand3_1 _10173_ (.A(_03474_),
    .B(_03469_),
    .C(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__nand3_1 _10174_ (.A(_03470_),
    .B(_03473_),
    .C(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2_1 _10175_ (.A(_03480_),
    .B(_03470_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand2b_1 _10176_ (.A_N(_03121_),
    .B(net86),
    .Y(_03482_));
 sky130_fd_sc_hd__or2b_1 _10177_ (.A(_03116_),
    .B_N(_03128_),
    .X(_03483_));
 sky130_fd_sc_hd__xnor2_1 _10178_ (.A(_03119_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__o21bai_1 _10179_ (.A1(_03218_),
    .A2(_03435_),
    .B1_N(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(_03482_),
    .B(_03485_),
    .Y(_03487_));
 sky130_fd_sc_hd__nand2_1 _10181_ (.A(_03487_),
    .B(_02495_),
    .Y(_03488_));
 sky130_fd_sc_hd__nand3_1 _10182_ (.A(_03482_),
    .B(_03485_),
    .C(\sq.out[9] ),
    .Y(_03489_));
 sky130_fd_sc_hd__nand2_1 _10183_ (.A(_03488_),
    .B(_03489_),
    .Y(_03490_));
 sky130_fd_sc_hd__nand2_1 _10184_ (.A(_03490_),
    .B(_03460_),
    .Y(_03491_));
 sky130_fd_sc_hd__nand3b_1 _10185_ (.A_N(_03460_),
    .B(_03488_),
    .C(_03489_),
    .Y(_03492_));
 sky130_fd_sc_hd__nand2_1 _10186_ (.A(_03491_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__inv_2 _10187_ (.A(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2_1 _10188_ (.A(_03481_),
    .B(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__nand2_1 _10189_ (.A(_03495_),
    .B(_03491_),
    .Y(_03496_));
 sky130_fd_sc_hd__inv_6 _10190_ (.A(_03436_),
    .Y(_03498_));
 sky130_fd_sc_hd__or2_1 _10191_ (.A(_03132_),
    .B(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__buf_6 _10192_ (.A(_03498_),
    .X(\sq.out[4] ));
 sky130_fd_sc_hd__a21o_1 _10193_ (.A1(_03137_),
    .A2(_03138_),
    .B1(_03129_),
    .X(_03500_));
 sky130_fd_sc_hd__nand3_1 _10194_ (.A(\sq.out[4] ),
    .B(_03139_),
    .C(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__nand2_1 _10195_ (.A(_03499_),
    .B(_03501_),
    .Y(_03502_));
 sky130_fd_sc_hd__nand2_1 _10196_ (.A(_03502_),
    .B(_02504_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand3_2 _10197_ (.A(_03499_),
    .B(\sq.out[10] ),
    .C(_03501_),
    .Y(_03504_));
 sky130_fd_sc_hd__nand2_1 _10198_ (.A(_03503_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand2_1 _10199_ (.A(_03505_),
    .B(_03489_),
    .Y(_03506_));
 sky130_fd_sc_hd__nand3b_1 _10200_ (.A_N(_03489_),
    .B(_03503_),
    .C(_03504_),
    .Y(_03508_));
 sky130_fd_sc_hd__nand2_1 _10201_ (.A(_03506_),
    .B(_03508_),
    .Y(_03509_));
 sky130_fd_sc_hd__or2_1 _10202_ (.A(_03164_),
    .B(_03140_),
    .X(_03510_));
 sky130_fd_sc_hd__nand2_1 _10203_ (.A(_03140_),
    .B(_03164_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(_03510_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_1 _10205_ (.A(_03436_),
    .B(_03159_),
    .Y(_03513_));
 sky130_fd_sc_hd__o21ai_2 _10206_ (.A1(_03512_),
    .A2(net86),
    .B1(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__nor2_1 _10207_ (.A(_02345_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__inv_2 _10208_ (.A(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_1 _10209_ (.A(_03514_),
    .B(_02345_),
    .Y(_03517_));
 sky130_fd_sc_hd__nand2_1 _10210_ (.A(_03516_),
    .B(_03517_),
    .Y(_03519_));
 sky130_fd_sc_hd__nor2_1 _10211_ (.A(_03504_),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__inv_2 _10212_ (.A(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__nand2_1 _10213_ (.A(_03519_),
    .B(_03504_),
    .Y(_03522_));
 sky130_fd_sc_hd__nand2_1 _10214_ (.A(_03521_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__nor2_1 _10215_ (.A(_03509_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__nand2_1 _10216_ (.A(_03496_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__o21a_1 _10217_ (.A1(_03520_),
    .A2(_03506_),
    .B1(_03522_),
    .X(_03526_));
 sky130_fd_sc_hd__nand2_1 _10218_ (.A(_03525_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__xor2_1 _10219_ (.A(_03186_),
    .B(_03167_),
    .X(_03528_));
 sky130_fd_sc_hd__nand2_1 _10220_ (.A(net86),
    .B(_03174_),
    .Y(_03530_));
 sky130_fd_sc_hd__o21ai_2 _10221_ (.A1(_03528_),
    .A2(net86),
    .B1(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__nor2_1 _10222_ (.A(_00844_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__inv_2 _10223_ (.A(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__nand2_1 _10224_ (.A(_03531_),
    .B(_00844_),
    .Y(_03534_));
 sky130_fd_sc_hd__nand2_1 _10225_ (.A(_03533_),
    .B(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _10226_ (.A(_03511_),
    .B(_03163_),
    .Y(_03536_));
 sky130_fd_sc_hd__xor2_1 _10227_ (.A(_03156_),
    .B(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__nand2_1 _10228_ (.A(net86),
    .B(_03144_),
    .Y(_03538_));
 sky130_fd_sc_hd__o21ai_2 _10229_ (.A1(_03537_),
    .A2(_03437_),
    .B1(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__or2_1 _10230_ (.A(_02826_),
    .B(_03539_),
    .X(_03541_));
 sky130_fd_sc_hd__nand2_1 _10231_ (.A(_03535_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nor2_1 _10232_ (.A(_03541_),
    .B(_03535_),
    .Y(_03543_));
 sky130_fd_sc_hd__inv_2 _10233_ (.A(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__nand2_1 _10234_ (.A(_03539_),
    .B(_02826_),
    .Y(_03545_));
 sky130_fd_sc_hd__nand2_1 _10235_ (.A(_03541_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand2_1 _10236_ (.A(_03546_),
    .B(_03516_),
    .Y(_03547_));
 sky130_fd_sc_hd__nand3_1 _10237_ (.A(_03541_),
    .B(_03515_),
    .C(_03545_),
    .Y(_03548_));
 sky130_fd_sc_hd__nand2_1 _10238_ (.A(_03547_),
    .B(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__inv_4 _10239_ (.A(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__o21ai_1 _10240_ (.A1(_03543_),
    .A2(_03547_),
    .B1(_03542_),
    .Y(_03552_));
 sky130_fd_sc_hd__a41o_1 _10241_ (.A1(_03527_),
    .A2(_03542_),
    .A3(_03544_),
    .A4(_03550_),
    .B1(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__nand2_1 _10242_ (.A(_03449_),
    .B(_02856_),
    .Y(_03554_));
 sky130_fd_sc_hd__nand2_1 _10243_ (.A(_03451_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nand2_1 _10244_ (.A(_03555_),
    .B(_03533_),
    .Y(_03556_));
 sky130_fd_sc_hd__nand3_1 _10245_ (.A(_03451_),
    .B(_03532_),
    .C(_03554_),
    .Y(_03557_));
 sky130_fd_sc_hd__nand2_1 _10246_ (.A(_03556_),
    .B(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__clkinvlp_2 _10247_ (.A(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__nand2_1 _10248_ (.A(_03553_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__nand2_1 _10249_ (.A(_03560_),
    .B(_03556_),
    .Y(_03561_));
 sky130_fd_sc_hd__or2_1 _10250_ (.A(_03455_),
    .B(_03561_),
    .X(_03563_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(_03561_),
    .B(_03455_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand2_1 _10252_ (.A(_03563_),
    .B(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__nor2_1 _10253_ (.A(_03217_),
    .B(_03435_),
    .Y(_03566_));
 sky130_fd_sc_hd__nand2_1 _10254_ (.A(_03566_),
    .B(_03209_),
    .Y(_03567_));
 sky130_fd_sc_hd__or2_1 _10255_ (.A(_03210_),
    .B(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__or2_1 _10256_ (.A(_03213_),
    .B(_03568_),
    .X(_03569_));
 sky130_fd_sc_hd__nand2_1 _10257_ (.A(_03568_),
    .B(_03213_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand2_1 _10258_ (.A(_03569_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__nand2_1 _10259_ (.A(_03567_),
    .B(_03210_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2_1 _10260_ (.A(_03568_),
    .B(_03572_),
    .Y(_03574_));
 sky130_fd_sc_hd__inv_2 _10261_ (.A(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__or2_1 _10262_ (.A(_03209_),
    .B(_03566_),
    .X(_03576_));
 sky130_fd_sc_hd__and2_1 _10263_ (.A(_03576_),
    .B(_03567_),
    .X(_03577_));
 sky130_fd_sc_hd__nand2_1 _10264_ (.A(_03575_),
    .B(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__nand3_2 _10265_ (.A(_03498_),
    .B(_03389_),
    .C(_03408_),
    .Y(_03579_));
 sky130_fd_sc_hd__or2_1 _10266_ (.A(_03433_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__or2_1 _10267_ (.A(_03414_),
    .B(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__or2_1 _10268_ (.A(_03416_),
    .B(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__or2_1 _10269_ (.A(_03418_),
    .B(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__xnor2_2 _10270_ (.A(_03421_),
    .B(_03583_),
    .Y(_03585_));
 sky130_fd_sc_hd__nor3_2 _10271_ (.A(_03571_),
    .B(_03578_),
    .C(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__inv_1 _10272_ (.A(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__and2_1 _10273_ (.A(_03195_),
    .B(_03196_),
    .X(_03588_));
 sky130_fd_sc_hd__or3_1 _10274_ (.A(_03216_),
    .B(_03217_),
    .C(_03435_),
    .X(_03589_));
 sky130_fd_sc_hd__xor2_1 _10275_ (.A(_03588_),
    .B(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__a21bo_1 _10276_ (.A1(_03569_),
    .A2(_03214_),
    .B1_N(_03589_),
    .X(_03591_));
 sky130_fd_sc_hd__or2_1 _10277_ (.A(_03590_),
    .B(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(_03235_),
    .B(_03261_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_1 _10279_ (.A(_03593_),
    .B(_03259_),
    .Y(_03594_));
 sky130_fd_sc_hd__or2_1 _10280_ (.A(_03254_),
    .B(_03594_),
    .X(_03596_));
 sky130_fd_sc_hd__nand2_1 _10281_ (.A(_03594_),
    .B(_03254_),
    .Y(_03597_));
 sky130_fd_sc_hd__a21o_1 _10282_ (.A1(_03596_),
    .A2(_03597_),
    .B1(_03437_),
    .X(_03598_));
 sky130_fd_sc_hd__nand2_1 _10283_ (.A(_03438_),
    .B(_03241_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _10284_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__nand2_1 _10285_ (.A(_03600_),
    .B(\sq.out[18] ),
    .Y(_03601_));
 sky130_fd_sc_hd__inv_2 _10286_ (.A(_03336_),
    .Y(_03602_));
 sky130_fd_sc_hd__or2_1 _10287_ (.A(_03347_),
    .B(_03263_),
    .X(_03603_));
 sky130_fd_sc_hd__or2_1 _10288_ (.A(_03602_),
    .B(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__nand2_1 _10289_ (.A(_03603_),
    .B(_03602_),
    .Y(_03605_));
 sky130_fd_sc_hd__nand2_1 _10290_ (.A(_03604_),
    .B(_03605_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(_03437_),
    .B(_03329_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21ai_4 _10292_ (.A1(_03607_),
    .A2(net97),
    .B1(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__nor2_1 _10293_ (.A(_05140_),
    .B(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand2_1 _10294_ (.A(_03609_),
    .B(_05140_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand2b_1 _10295_ (.A_N(_03610_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__or2_1 _10296_ (.A(_03601_),
    .B(_03612_),
    .X(_03613_));
 sky130_fd_sc_hd__nand2_1 _10297_ (.A(_03612_),
    .B(_03601_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand2_1 _10298_ (.A(_03613_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__or2_1 _10299_ (.A(_03261_),
    .B(_03235_),
    .X(_03616_));
 sky130_fd_sc_hd__nand2_1 _10300_ (.A(_03616_),
    .B(_03593_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _10301_ (.A(_03438_),
    .B(_03249_),
    .Y(_03619_));
 sky130_fd_sc_hd__o21ai_2 _10302_ (.A1(_03618_),
    .A2(_03438_),
    .B1(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__or2_1 _10303_ (.A(_02877_),
    .B(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__inv_2 _10304_ (.A(_03600_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand2_1 _10305_ (.A(_03622_),
    .B(_01712_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2_1 _10306_ (.A(_03623_),
    .B(_03601_),
    .Y(_03624_));
 sky130_fd_sc_hd__or2_1 _10307_ (.A(_03621_),
    .B(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__nand2_1 _10308_ (.A(_03624_),
    .B(_03621_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand2_1 _10309_ (.A(_03625_),
    .B(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__nor2_1 _10310_ (.A(_03615_),
    .B(_03627_),
    .Y(_03629_));
 sky130_fd_sc_hd__clkinvlp_2 _10311_ (.A(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__nand3_1 _10312_ (.A(_03559_),
    .B(_03452_),
    .C(_03454_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_1 _10313_ (.A(_03544_),
    .B(_03542_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand2b_1 _10314_ (.A_N(_03632_),
    .B(_03550_),
    .Y(_03633_));
 sky130_fd_sc_hd__nor2_1 _10315_ (.A(_03631_),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__nand2_1 _10316_ (.A(_03527_),
    .B(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__nor2_1 _10317_ (.A(_03558_),
    .B(_03455_),
    .Y(_03636_));
 sky130_fd_sc_hd__o21ai_1 _10318_ (.A1(_03556_),
    .A2(_03455_),
    .B1(_03452_),
    .Y(_03637_));
 sky130_fd_sc_hd__a21oi_1 _10319_ (.A1(_03552_),
    .A2(_03636_),
    .B1(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__nand2_1 _10320_ (.A(_03638_),
    .B(_03635_),
    .Y(_03640_));
 sky130_fd_sc_hd__nand2_1 _10321_ (.A(_03620_),
    .B(_02877_),
    .Y(_03641_));
 sky130_fd_sc_hd__nand2_1 _10322_ (.A(_03621_),
    .B(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__a21bo_1 _10323_ (.A1(_03190_),
    .A2(_03109_),
    .B1_N(_03110_),
    .X(_03643_));
 sky130_fd_sc_hd__nand2_1 _10324_ (.A(_03643_),
    .B(_03230_),
    .Y(_03644_));
 sky130_fd_sc_hd__or2_1 _10325_ (.A(_03230_),
    .B(_03643_),
    .X(_03645_));
 sky130_fd_sc_hd__a21oi_1 _10326_ (.A1(_03644_),
    .A2(_03645_),
    .B1(_03438_),
    .Y(_03646_));
 sky130_fd_sc_hd__a21o_1 _10327_ (.A1(_03224_),
    .A2(_03438_),
    .B1(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__or2_1 _10328_ (.A(_00092_),
    .B(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__nor2_1 _10329_ (.A(_03642_),
    .B(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__nand2_1 _10330_ (.A(_03648_),
    .B(_03642_),
    .Y(_03651_));
 sky130_fd_sc_hd__or2b_1 _10331_ (.A(_03649_),
    .B_N(_03651_),
    .X(_03652_));
 sky130_fd_sc_hd__inv_2 _10332_ (.A(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__nand2_1 _10333_ (.A(_03647_),
    .B(_00092_),
    .Y(_03654_));
 sky130_fd_sc_hd__nand2_1 _10334_ (.A(_03648_),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__or2_1 _10335_ (.A(_03443_),
    .B(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__nand2_1 _10336_ (.A(_03655_),
    .B(_03443_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand2_1 _10337_ (.A(_03656_),
    .B(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__inv_2 _10338_ (.A(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand3_2 _10339_ (.A(_03640_),
    .B(_03653_),
    .C(_03659_),
    .Y(_03660_));
 sky130_fd_sc_hd__nor2_4 _10340_ (.A(_03630_),
    .B(_03660_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand3_1 _10341_ (.A(\sq.out[4] ),
    .B(_03389_),
    .C(_03391_),
    .Y(_03663_));
 sky130_fd_sc_hd__nor2b_1 _10342_ (.A(_03663_),
    .B_N(_03402_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand2_1 _10343_ (.A(_03664_),
    .B(_03405_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2b_1 _10344_ (.A_N(_03665_),
    .B(_03400_),
    .Y(_03666_));
 sky130_fd_sc_hd__a21o_1 _10345_ (.A1(_03664_),
    .A2(_03405_),
    .B1(_03400_),
    .X(_03667_));
 sky130_fd_sc_hd__nand2_1 _10346_ (.A(_03666_),
    .B(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__inv_4 _10347_ (.A(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__or2_1 _10348_ (.A(_03405_),
    .B(_03664_),
    .X(_03670_));
 sky130_fd_sc_hd__and2_1 _10349_ (.A(_03670_),
    .B(_03665_),
    .X(_03671_));
 sky130_fd_sc_hd__xor2_1 _10350_ (.A(_03402_),
    .B(_03663_),
    .X(_03673_));
 sky130_fd_sc_hd__a21bo_1 _10351_ (.A1(_03352_),
    .A2(_03370_),
    .B1_N(_03390_),
    .X(_03674_));
 sky130_fd_sc_hd__nand2_1 _10352_ (.A(_03674_),
    .B(_03380_),
    .Y(_03675_));
 sky130_fd_sc_hd__and3_1 _10353_ (.A(\sq.out[4] ),
    .B(_03378_),
    .C(_03675_),
    .X(_03676_));
 sky130_fd_sc_hd__xor2_1 _10354_ (.A(_03385_),
    .B(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__nor2_1 _10355_ (.A(_03673_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__nand3_1 _10356_ (.A(_03669_),
    .B(_03671_),
    .C(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__a21o_1 _10357_ (.A1(_03263_),
    .A2(_03342_),
    .B1(_03349_),
    .X(_03680_));
 sky130_fd_sc_hd__or2b_1 _10358_ (.A(_03321_),
    .B_N(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__a21o_1 _10359_ (.A1(_03681_),
    .A2(_03345_),
    .B1(_03296_),
    .X(_03682_));
 sky130_fd_sc_hd__nand2_1 _10360_ (.A(_03682_),
    .B(_03295_),
    .Y(_03684_));
 sky130_fd_sc_hd__xor2_1 _10361_ (.A(_03283_),
    .B(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__nand2_1 _10362_ (.A(_03685_),
    .B(\sq.out[4] ),
    .Y(_03686_));
 sky130_fd_sc_hd__nand2_1 _10363_ (.A(_03439_),
    .B(_03276_),
    .Y(_03687_));
 sky130_fd_sc_hd__nand2_1 _10364_ (.A(_03686_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__nand2_1 _10365_ (.A(_03688_),
    .B(\sq.out[24] ),
    .Y(_03689_));
 sky130_fd_sc_hd__xor2_1 _10366_ (.A(_03369_),
    .B(_03352_),
    .X(_03690_));
 sky130_fd_sc_hd__nor2_1 _10367_ (.A(_03690_),
    .B(_03438_),
    .Y(_03691_));
 sky130_fd_sc_hd__o21ba_1 _10368_ (.A1(_03358_),
    .A2(\sq.out[4] ),
    .B1_N(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__nand2_1 _10369_ (.A(_03689_),
    .B(_03692_),
    .Y(_03693_));
 sky130_fd_sc_hd__inv_2 _10370_ (.A(_03692_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand3_1 _10371_ (.A(_03688_),
    .B(\sq.out[24] ),
    .C(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand2_1 _10372_ (.A(_03693_),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand3_1 _10373_ (.A(_03686_),
    .B(_01081_),
    .C(_03687_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand2_1 _10374_ (.A(_03689_),
    .B(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__nand3_1 _10375_ (.A(_03681_),
    .B(_03296_),
    .C(_03345_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand3_1 _10376_ (.A(_03682_),
    .B(_03498_),
    .C(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__nand2_1 _10377_ (.A(net97),
    .B(_03284_),
    .Y(_03702_));
 sky130_fd_sc_hd__nand2_1 _10378_ (.A(_03701_),
    .B(_03702_),
    .Y(_03703_));
 sky130_fd_sc_hd__or2_1 _10379_ (.A(_01993_),
    .B(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__nand2_1 _10380_ (.A(_03699_),
    .B(_03704_),
    .Y(_03706_));
 sky130_fd_sc_hd__nand3b_1 _10381_ (.A_N(_03704_),
    .B(_03689_),
    .C(_03698_),
    .Y(_03707_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(_03706_),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__nor2_1 _10383_ (.A(_03697_),
    .B(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__or2_1 _10384_ (.A(_03380_),
    .B(_03674_),
    .X(_03710_));
 sky130_fd_sc_hd__and2_1 _10385_ (.A(_03439_),
    .B(_03375_),
    .X(_03711_));
 sky130_fd_sc_hd__a31o_1 _10386_ (.A1(_03710_),
    .A2(\sq.out[4] ),
    .A3(_03675_),
    .B1(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__a21bo_1 _10387_ (.A1(_03352_),
    .A2(_03367_),
    .B1_N(_03368_),
    .X(_03713_));
 sky130_fd_sc_hd__xor2_1 _10388_ (.A(_03364_),
    .B(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__nand2_1 _10389_ (.A(_03439_),
    .B(_03361_),
    .Y(_03715_));
 sky130_fd_sc_hd__o21ai_2 _10390_ (.A1(_03439_),
    .A2(_03714_),
    .B1(_03715_),
    .Y(_03717_));
 sky130_fd_sc_hd__or2_1 _10391_ (.A(_03717_),
    .B(_03695_),
    .X(_03718_));
 sky130_fd_sc_hd__nand2_1 _10392_ (.A(_03695_),
    .B(_03717_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _10393_ (.A(_03718_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__nor2_1 _10394_ (.A(_03712_),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__nand2_1 _10395_ (.A(_03709_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__nor2_1 _10396_ (.A(_03679_),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__nand2_1 _10397_ (.A(_03680_),
    .B(_03314_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2_1 _10398_ (.A(_03724_),
    .B(_03312_),
    .Y(_03725_));
 sky130_fd_sc_hd__or2_1 _10399_ (.A(_03320_),
    .B(_03725_),
    .X(_03726_));
 sky130_fd_sc_hd__nand2_1 _10400_ (.A(_03725_),
    .B(_03320_),
    .Y(_03728_));
 sky130_fd_sc_hd__a21o_1 _10401_ (.A1(_03726_),
    .A2(_03728_),
    .B1(net97),
    .X(_03729_));
 sky130_fd_sc_hd__nand2_1 _10402_ (.A(_03438_),
    .B(_03292_),
    .Y(_03730_));
 sky130_fd_sc_hd__nand2_1 _10403_ (.A(_03729_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__inv_2 _10404_ (.A(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_1 _10405_ (.A(_03732_),
    .B(_02009_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand2_1 _10406_ (.A(_03731_),
    .B(\sq.out[22] ),
    .Y(_03734_));
 sky130_fd_sc_hd__or2_1 _10407_ (.A(_03314_),
    .B(_03680_),
    .X(_03735_));
 sky130_fd_sc_hd__nand2_1 _10408_ (.A(_03735_),
    .B(_03724_),
    .Y(_03736_));
 sky130_fd_sc_hd__nand2_1 _10409_ (.A(_03436_),
    .B(_03306_),
    .Y(_03737_));
 sky130_fd_sc_hd__o21ai_2 _10410_ (.A1(_03736_),
    .A2(_03436_),
    .B1(_03737_),
    .Y(_03739_));
 sky130_fd_sc_hd__nor2_1 _10411_ (.A(_02927_),
    .B(_03739_),
    .Y(_03740_));
 sky130_fd_sc_hd__a21o_1 _10412_ (.A1(_03733_),
    .A2(_03734_),
    .B1(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__nand3_1 _10413_ (.A(_03733_),
    .B(_03734_),
    .C(_03740_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _10414_ (.A(_03741_),
    .B(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand2_1 _10415_ (.A(_03703_),
    .B(_01993_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_1 _10416_ (.A(_03704_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__nor2_1 _10417_ (.A(_03734_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__nand2_1 _10418_ (.A(_03745_),
    .B(_03734_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand2b_1 _10419_ (.A_N(_03746_),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__nor2_1 _10420_ (.A(_03743_),
    .B(_03748_),
    .Y(_03750_));
 sky130_fd_sc_hd__nand2_1 _10421_ (.A(_03605_),
    .B(_03335_),
    .Y(_03751_));
 sky130_fd_sc_hd__xor2_1 _10422_ (.A(_03341_),
    .B(_03751_),
    .X(_03752_));
 sky130_fd_sc_hd__nor2_1 _10423_ (.A(_03302_),
    .B(_03498_),
    .Y(_03753_));
 sky130_fd_sc_hd__a21oi_2 _10424_ (.A1(\sq.out[4] ),
    .A2(_03752_),
    .B1(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__or2_1 _10425_ (.A(_01730_),
    .B(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__and2_1 _10426_ (.A(_03739_),
    .B(_02927_),
    .X(_03756_));
 sky130_fd_sc_hd__or2_1 _10427_ (.A(_03740_),
    .B(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__nor2_1 _10428_ (.A(_03755_),
    .B(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_1 _10429_ (.A(_03757_),
    .B(_03755_),
    .Y(_03759_));
 sky130_fd_sc_hd__nand2b_1 _10430_ (.A_N(_03758_),
    .B(_03759_),
    .Y(_03761_));
 sky130_fd_sc_hd__nand2_1 _10431_ (.A(_03754_),
    .B(_01730_),
    .Y(_03762_));
 sky130_fd_sc_hd__nand2_1 _10432_ (.A(_03755_),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand2b_1 _10433_ (.A_N(_03763_),
    .B(_03610_),
    .Y(_03764_));
 sky130_fd_sc_hd__o21ai_1 _10434_ (.A1(_05140_),
    .A2(_03609_),
    .B1(_03763_),
    .Y(_03765_));
 sky130_fd_sc_hd__nand2_1 _10435_ (.A(_03764_),
    .B(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__nor2_1 _10436_ (.A(_03761_),
    .B(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__nand2_1 _10437_ (.A(_03750_),
    .B(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__inv_2 _10438_ (.A(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__nand3_2 _10439_ (.A(_03662_),
    .B(_03723_),
    .C(_03769_),
    .Y(_03770_));
 sky130_fd_sc_hd__o21ai_1 _10440_ (.A1(_03649_),
    .A2(_03657_),
    .B1(_03651_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand2_1 _10441_ (.A(_03772_),
    .B(_03629_),
    .Y(_03773_));
 sky130_fd_sc_hd__o21a_1 _10442_ (.A1(_03626_),
    .A2(_03615_),
    .B1(_03614_),
    .X(_03774_));
 sky130_fd_sc_hd__nand2_1 _10443_ (.A(_03773_),
    .B(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_1 _10444_ (.A(_03769_),
    .B(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__o21ai_1 _10445_ (.A1(_03758_),
    .A2(_03765_),
    .B1(_03759_),
    .Y(_03777_));
 sky130_fd_sc_hd__o21ai_1 _10446_ (.A1(_03746_),
    .A2(_03741_),
    .B1(_03747_),
    .Y(_03778_));
 sky130_fd_sc_hd__a21oi_1 _10447_ (.A1(_03750_),
    .A2(_03777_),
    .B1(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__nand2_2 _10448_ (.A(_03776_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__o21ai_1 _10449_ (.A1(_03697_),
    .A2(_03706_),
    .B1(_03693_),
    .Y(_03781_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_03781_),
    .B(_03721_),
    .Y(_03783_));
 sky130_fd_sc_hd__a21oi_1 _10451_ (.A1(_03695_),
    .A2(_03717_),
    .B1(_03712_),
    .Y(_03784_));
 sky130_fd_sc_hd__nand3b_1 _10452_ (.A_N(_03679_),
    .B(_03783_),
    .C(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__a21oi_2 _10453_ (.A1(_03780_),
    .A2(_03723_),
    .B1(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__nand2_1 _10454_ (.A(_03582_),
    .B(_03418_),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _10455_ (.A(_03583_),
    .B(_03787_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _10456_ (.A(_03581_),
    .B(_03416_),
    .Y(_03789_));
 sky130_fd_sc_hd__nand2_1 _10457_ (.A(_03582_),
    .B(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__or2_1 _10458_ (.A(_03424_),
    .B(_03579_),
    .X(_03791_));
 sky130_fd_sc_hd__nor2b_1 _10459_ (.A(_03791_),
    .B_N(_03428_),
    .Y(_03792_));
 sky130_fd_sc_hd__nand2_1 _10460_ (.A(_03792_),
    .B(_03426_),
    .Y(_03794_));
 sky130_fd_sc_hd__xnor2_1 _10461_ (.A(_03432_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _10462_ (.A(_03580_),
    .B(_03414_),
    .Y(_03796_));
 sky130_fd_sc_hd__and2_1 _10463_ (.A(_03581_),
    .B(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__nor3b_1 _10464_ (.A(_03790_),
    .B(_03795_),
    .C_N(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hd__or2_1 _10465_ (.A(_03426_),
    .B(_03792_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2_1 _10466_ (.A(_03799_),
    .B(_03794_),
    .Y(_03800_));
 sky130_fd_sc_hd__and2b_1 _10467_ (.A_N(_03428_),
    .B(_03791_),
    .X(_03801_));
 sky130_fd_sc_hd__nor2_1 _10468_ (.A(_03801_),
    .B(_03792_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _10469_ (.A(_03579_),
    .B(_03424_),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _10470_ (.A(_03791_),
    .B(_03803_),
    .Y(_03805_));
 sky130_fd_sc_hd__inv_2 _10471_ (.A(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_1 _10472_ (.A(_03802_),
    .B(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__xnor2_2 _10473_ (.A(_03397_),
    .B(_03666_),
    .Y(_03808_));
 sky130_fd_sc_hd__nor3b_1 _10474_ (.A(_03800_),
    .B(_03807_),
    .C_N(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__and3b_1 _10475_ (.A_N(_03788_),
    .B(_03798_),
    .C(_03809_),
    .X(_03810_));
 sky130_fd_sc_hd__nand3_2 _10476_ (.A(_03770_),
    .B(_03786_),
    .C(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__nor3_2 _10477_ (.A(_03587_),
    .B(_03592_),
    .C(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hd__a41o_1 _10478_ (.A1(_03566_),
    .A2(_03588_),
    .A3(_03209_),
    .A4(_03215_),
    .B1(_03199_),
    .X(_03813_));
 sky130_fd_sc_hd__or2b_1 _10479_ (.A(_03589_),
    .B_N(_03200_),
    .X(_03814_));
 sky130_fd_sc_hd__nand2_1 _10480_ (.A(_03813_),
    .B(_03814_),
    .Y(_03816_));
 sky130_fd_sc_hd__inv_1 _10481_ (.A(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__inv_2 _10482_ (.A(_03202_),
    .Y(_03818_));
 sky130_fd_sc_hd__nand2_2 _10483_ (.A(_03814_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__nand3_2 _10484_ (.A(_03812_),
    .B(_03817_),
    .C(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__buf_6 _10485_ (.A(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__buf_6 _10486_ (.A(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__mux2_2 _10487_ (.A0(_03441_),
    .A1(_03565_),
    .S(_03822_),
    .X(_03823_));
 sky130_fd_sc_hd__or2_1 _10488_ (.A(_00092_),
    .B(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__nand2_1 _10489_ (.A(_03823_),
    .B(_00092_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2_1 _10490_ (.A(_03824_),
    .B(_03825_),
    .Y(_03827_));
 sky130_fd_sc_hd__or2_1 _10491_ (.A(_03559_),
    .B(_03553_),
    .X(_03828_));
 sky130_fd_sc_hd__clkinvlp_2 _10492_ (.A(_03819_),
    .Y(_03829_));
 sky130_fd_sc_hd__nor2_2 _10493_ (.A(_03587_),
    .B(_03811_),
    .Y(_03830_));
 sky130_fd_sc_hd__clkinvlp_2 _10494_ (.A(_03592_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand3_2 _10495_ (.A(_03830_),
    .B(_03817_),
    .C(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__nor2_4 _10496_ (.A(_03829_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__buf_6 _10497_ (.A(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__and2_1 _10498_ (.A(net95),
    .B(_03449_),
    .X(_03835_));
 sky130_fd_sc_hd__a31o_1 _10499_ (.A1(_03822_),
    .A2(_03560_),
    .A3(_03828_),
    .B1(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__or2_1 _10500_ (.A(_02843_),
    .B(_03836_),
    .X(_03838_));
 sky130_fd_sc_hd__nand2_1 _10501_ (.A(_03827_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__nand2_1 _10502_ (.A(_03640_),
    .B(_03659_),
    .Y(_03840_));
 sky130_fd_sc_hd__or2_1 _10503_ (.A(_03659_),
    .B(_03640_),
    .X(_03841_));
 sky130_fd_sc_hd__nand3_1 _10504_ (.A(_03822_),
    .B(_03840_),
    .C(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__buf_6 _10505_ (.A(_03834_),
    .X(_03843_));
 sky130_fd_sc_hd__nand2_1 _10506_ (.A(_03843_),
    .B(_03647_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _10507_ (.A(_03842_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__or2_1 _10508_ (.A(_02877_),
    .B(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__nand2_1 _10509_ (.A(_03845_),
    .B(_02877_),
    .Y(_03847_));
 sky130_fd_sc_hd__nand2_1 _10510_ (.A(_03846_),
    .B(_03847_),
    .Y(_03849_));
 sky130_fd_sc_hd__or2_1 _10511_ (.A(_03849_),
    .B(_03824_),
    .X(_03850_));
 sky130_fd_sc_hd__nand2_1 _10512_ (.A(_03824_),
    .B(_03849_),
    .Y(_03851_));
 sky130_fd_sc_hd__nand2_1 _10513_ (.A(_03850_),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__o21ai_1 _10514_ (.A1(_03839_),
    .A2(_03852_),
    .B1(_03851_),
    .Y(_03853_));
 sky130_fd_sc_hd__inv_2 _10515_ (.A(_03811_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand3_1 _10516_ (.A(_03854_),
    .B(_03586_),
    .C(_03831_),
    .Y(_03855_));
 sky130_fd_sc_hd__nor2_1 _10517_ (.A(_03816_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__nand3_2 _10518_ (.A(_03856_),
    .B(_03439_),
    .C(_03819_),
    .Y(_03857_));
 sky130_fd_sc_hd__nor3_1 _10519_ (.A(\sq.out[6] ),
    .B(_03373_),
    .C(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__buf_6 _10520_ (.A(_03821_),
    .X(\sq.out[3] ));
 sky130_fd_sc_hd__and2b_1 _10521_ (.A_N(_03477_),
    .B(_03468_),
    .X(_03860_));
 sky130_fd_sc_hd__inv_2 _10522_ (.A(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__a21oi_1 _10523_ (.A1(\sq.out[3] ),
    .A2(_03373_),
    .B1(_03861_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _10524_ (.A(_03821_),
    .B(_03861_),
    .Y(_03863_));
 sky130_fd_sc_hd__nand2_1 _10525_ (.A(_03857_),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__nand2_1 _10526_ (.A(_03864_),
    .B(\sq.out[6] ),
    .Y(_03865_));
 sky130_fd_sc_hd__nand3_1 _10527_ (.A(_03857_),
    .B(_03863_),
    .C(_02898_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _10528_ (.A(_03865_),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__or2_1 _10529_ (.A(_03373_),
    .B(_03857_),
    .X(_03868_));
 sky130_fd_sc_hd__nand2_1 _10530_ (.A(_03867_),
    .B(_03868_),
    .Y(_03870_));
 sky130_fd_sc_hd__o21ai_1 _10531_ (.A1(_03858_),
    .A2(_03862_),
    .B1(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__nand3_1 _10532_ (.A(_03834_),
    .B(_03373_),
    .C(_03439_),
    .Y(_03872_));
 sky130_fd_sc_hd__nand2_1 _10533_ (.A(_03821_),
    .B(_03465_),
    .Y(_03873_));
 sky130_fd_sc_hd__nand2_2 _10534_ (.A(_03872_),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nand2_2 _10535_ (.A(_03874_),
    .B(\sq.out[7] ),
    .Y(_03875_));
 sky130_fd_sc_hd__nand3_1 _10536_ (.A(_03872_),
    .B(_03112_),
    .C(_03873_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _10537_ (.A(_03875_),
    .B(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _10538_ (.A(_03877_),
    .B(_03865_),
    .Y(_03878_));
 sky130_fd_sc_hd__nand3b_1 _10539_ (.A_N(_03865_),
    .B(_03875_),
    .C(_03876_),
    .Y(_03879_));
 sky130_fd_sc_hd__nand3_2 _10540_ (.A(_03871_),
    .B(_03878_),
    .C(_03879_),
    .Y(_03881_));
 sky130_fd_sc_hd__nand2_2 _10541_ (.A(_03881_),
    .B(_03878_),
    .Y(_03882_));
 sky130_fd_sc_hd__a21oi_1 _10542_ (.A1(_03470_),
    .A2(_03473_),
    .B1(_03479_),
    .Y(_03883_));
 sky130_fd_sc_hd__nand3b_1 _10543_ (.A_N(_03883_),
    .B(_03821_),
    .C(_03480_),
    .Y(_03884_));
 sky130_fd_sc_hd__nand2_1 _10544_ (.A(_03834_),
    .B(_03458_),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _10545_ (.A(_03884_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand2_1 _10546_ (.A(_03886_),
    .B(_02495_),
    .Y(_03887_));
 sky130_fd_sc_hd__nand3_2 _10547_ (.A(_03884_),
    .B(\sq.out[9] ),
    .C(_03885_),
    .Y(_03888_));
 sky130_fd_sc_hd__nand2_1 _10548_ (.A(_03833_),
    .B(_03471_),
    .Y(_03889_));
 sky130_fd_sc_hd__a21oi_1 _10549_ (.A1(_03474_),
    .A2(_03469_),
    .B1(_03478_),
    .Y(_03890_));
 sky130_fd_sc_hd__or2b_1 _10550_ (.A(_03890_),
    .B_N(_03479_),
    .X(_03892_));
 sky130_fd_sc_hd__nand2_1 _10551_ (.A(_03820_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_1 _10552_ (.A(_03889_),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__nor2_1 _10553_ (.A(_02498_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__a21o_1 _10554_ (.A1(_03887_),
    .A2(_03888_),
    .B1(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__nand3_1 _10555_ (.A(_03887_),
    .B(_03888_),
    .C(_03895_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_1 _10556_ (.A(_03896_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__inv_2 _10557_ (.A(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _10558_ (.A(_03894_),
    .B(_02498_),
    .Y(_03900_));
 sky130_fd_sc_hd__nand2b_1 _10559_ (.A_N(_03895_),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__nor2_1 _10560_ (.A(_03875_),
    .B(_03901_),
    .Y(_03903_));
 sky130_fd_sc_hd__nand2_1 _10561_ (.A(_03901_),
    .B(_03875_),
    .Y(_03904_));
 sky130_fd_sc_hd__and2b_1 _10562_ (.A_N(_03903_),
    .B(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__nand3_1 _10563_ (.A(_03882_),
    .B(_03899_),
    .C(_03905_),
    .Y(_03906_));
 sky130_fd_sc_hd__o21a_1 _10564_ (.A1(_03904_),
    .A2(_03898_),
    .B1(_03896_),
    .X(_03907_));
 sky130_fd_sc_hd__nand2_1 _10565_ (.A(_03906_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__or2_1 _10566_ (.A(_03494_),
    .B(_03481_),
    .X(_03909_));
 sky130_fd_sc_hd__nand3_1 _10567_ (.A(_03821_),
    .B(_03495_),
    .C(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _10568_ (.A(_03833_),
    .B(_03487_),
    .Y(_03911_));
 sky130_fd_sc_hd__nand2_1 _10569_ (.A(_03910_),
    .B(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__or2_1 _10570_ (.A(_02504_),
    .B(_03912_),
    .X(_03914_));
 sky130_fd_sc_hd__or2b_1 _10571_ (.A(_03496_),
    .B_N(_03509_),
    .X(_03915_));
 sky130_fd_sc_hd__a21o_1 _10572_ (.A1(_03495_),
    .A2(_03491_),
    .B1(_03509_),
    .X(_03916_));
 sky130_fd_sc_hd__nand2_1 _10573_ (.A(_03915_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__nand2_1 _10574_ (.A(_03833_),
    .B(_03502_),
    .Y(_03918_));
 sky130_fd_sc_hd__o21ai_2 _10575_ (.A1(_03917_),
    .A2(_03833_),
    .B1(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__or2_1 _10576_ (.A(_02345_),
    .B(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__nand2_1 _10577_ (.A(_03919_),
    .B(_02345_),
    .Y(_03921_));
 sky130_fd_sc_hd__nand2_1 _10578_ (.A(_03920_),
    .B(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__or2_1 _10579_ (.A(_03914_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__nand2_1 _10580_ (.A(_03922_),
    .B(_03914_),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _10581_ (.A(_03923_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__inv_2 _10582_ (.A(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2_1 _10583_ (.A(_03912_),
    .B(_02504_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand2_1 _10584_ (.A(_03914_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__or2_1 _10585_ (.A(_03888_),
    .B(_03929_),
    .X(_03930_));
 sky130_fd_sc_hd__nand2_1 _10586_ (.A(_03929_),
    .B(_03888_),
    .Y(_03931_));
 sky130_fd_sc_hd__nand2_1 _10587_ (.A(_03930_),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__inv_2 _10588_ (.A(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__nand3_1 _10589_ (.A(_03908_),
    .B(_03927_),
    .C(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__o21a_1 _10590_ (.A1(_03931_),
    .A2(_03926_),
    .B1(_03925_),
    .X(_03936_));
 sky130_fd_sc_hd__nand2_2 _10591_ (.A(_03934_),
    .B(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__nand2_1 _10592_ (.A(_03916_),
    .B(_03506_),
    .Y(_03938_));
 sky130_fd_sc_hd__xor2_1 _10593_ (.A(_03523_),
    .B(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__nand2_1 _10594_ (.A(_03834_),
    .B(_03514_),
    .Y(_03940_));
 sky130_fd_sc_hd__o21ai_2 _10595_ (.A1(_03939_),
    .A2(_03843_),
    .B1(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__or2_1 _10596_ (.A(_02826_),
    .B(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__nand2_1 _10597_ (.A(_03941_),
    .B(_02826_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _10598_ (.A(_03942_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__or2_1 _10599_ (.A(_03920_),
    .B(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__nand2_1 _10600_ (.A(_03944_),
    .B(_03920_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _10601_ (.A(_03945_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(_03527_),
    .B(_03550_),
    .Y(_03949_));
 sky130_fd_sc_hd__or2_1 _10603_ (.A(_03550_),
    .B(_03527_),
    .X(_03950_));
 sky130_fd_sc_hd__and2_1 _10604_ (.A(_03833_),
    .B(_03539_),
    .X(_03951_));
 sky130_fd_sc_hd__a31o_1 _10605_ (.A1(_03821_),
    .A2(_03949_),
    .A3(_03950_),
    .B1(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__or2_1 _10606_ (.A(_00844_),
    .B(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__nand2_1 _10607_ (.A(_03952_),
    .B(_00844_),
    .Y(_03954_));
 sky130_fd_sc_hd__nand2_1 _10608_ (.A(_03953_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__or2_1 _10609_ (.A(_03942_),
    .B(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__nand2_1 _10610_ (.A(_03955_),
    .B(_03942_),
    .Y(_03958_));
 sky130_fd_sc_hd__nand2_1 _10611_ (.A(_03956_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__nor2_1 _10612_ (.A(_03948_),
    .B(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_1 _10613_ (.A(_03937_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__o21a_1 _10614_ (.A1(_03947_),
    .A2(_03959_),
    .B1(_03958_),
    .X(_03962_));
 sky130_fd_sc_hd__nand2_1 _10615_ (.A(_03961_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__nand2_1 _10616_ (.A(_03949_),
    .B(_03547_),
    .Y(_03964_));
 sky130_fd_sc_hd__xor2_1 _10617_ (.A(_03632_),
    .B(_03964_),
    .X(_03965_));
 sky130_fd_sc_hd__nand2_1 _10618_ (.A(_03843_),
    .B(_03531_),
    .Y(_03966_));
 sky130_fd_sc_hd__o21ai_2 _10619_ (.A1(_03965_),
    .A2(_03843_),
    .B1(_03966_),
    .Y(_03967_));
 sky130_fd_sc_hd__or2_1 _10620_ (.A(_02856_),
    .B(_03967_),
    .X(_03969_));
 sky130_fd_sc_hd__nand2_1 _10621_ (.A(_03967_),
    .B(_02856_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _10622_ (.A(_03969_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__or2_1 _10623_ (.A(_03971_),
    .B(_03953_),
    .X(_03972_));
 sky130_fd_sc_hd__nand2_1 _10624_ (.A(_03953_),
    .B(_03971_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _10625_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _10626_ (.A(_03836_),
    .B(_02843_),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_1 _10627_ (.A(_03838_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__or2_1 _10628_ (.A(_03969_),
    .B(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__nand2_1 _10629_ (.A(_03976_),
    .B(_03969_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_1 _10630_ (.A(_03977_),
    .B(_03978_),
    .Y(_03980_));
 sky130_fd_sc_hd__nor2_1 _10631_ (.A(_03974_),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_1 _10632_ (.A(_03963_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__o21a_1 _10633_ (.A1(_03973_),
    .A2(_03980_),
    .B1(_03978_),
    .X(_03983_));
 sky130_fd_sc_hd__nand2_1 _10634_ (.A(_03982_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__clkinvlp_2 _10635_ (.A(_03852_),
    .Y(_03985_));
 sky130_fd_sc_hd__or2_1 _10636_ (.A(_03838_),
    .B(_03827_),
    .X(_03986_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(_03986_),
    .B(_03839_),
    .Y(_03987_));
 sky130_fd_sc_hd__clkinvlp_2 _10638_ (.A(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand3_2 _10639_ (.A(_03984_),
    .B(_03985_),
    .C(_03988_),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2b_1 _10640_ (.A_N(_03853_),
    .B(_03989_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _10641_ (.A(_03840_),
    .B(_03657_),
    .Y(_03992_));
 sky130_fd_sc_hd__or2_1 _10642_ (.A(_03652_),
    .B(_03992_),
    .X(_03993_));
 sky130_fd_sc_hd__nand2_1 _10643_ (.A(_03992_),
    .B(_03652_),
    .Y(_03994_));
 sky130_fd_sc_hd__nand2_1 _10644_ (.A(_03993_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__mux2_1 _10645_ (.A0(_03620_),
    .A1(_03995_),
    .S(_03821_),
    .X(_03996_));
 sky130_fd_sc_hd__or2_1 _10646_ (.A(_01712_),
    .B(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__nand2_1 _10647_ (.A(_03996_),
    .B(_01712_),
    .Y(_03998_));
 sky130_fd_sc_hd__nand2_1 _10648_ (.A(_03997_),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__or2_1 _10649_ (.A(_03846_),
    .B(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__nand2_1 _10650_ (.A(_03999_),
    .B(_03846_),
    .Y(_04002_));
 sky130_fd_sc_hd__nand2_1 _10651_ (.A(_04000_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__or2b_1 _10652_ (.A(_03991_),
    .B_N(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__nand2b_1 _10653_ (.A_N(_04003_),
    .B(_03991_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand2_1 _10654_ (.A(_04004_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_1 _10655_ (.A(_03832_),
    .B(_03829_),
    .Y(_04007_));
 sky130_fd_sc_hd__inv_1 _10656_ (.A(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__nand2b_1 _10657_ (.A_N(_03772_),
    .B(_03660_),
    .Y(_04009_));
 sky130_fd_sc_hd__xor2_1 _10658_ (.A(_03627_),
    .B(_04009_),
    .X(_04010_));
 sky130_fd_sc_hd__or2_1 _10659_ (.A(_04010_),
    .B(net95),
    .X(_04011_));
 sky130_fd_sc_hd__nand2_1 _10660_ (.A(_03834_),
    .B(_03622_),
    .Y(_04013_));
 sky130_fd_sc_hd__nand2_1 _10661_ (.A(_04011_),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__inv_2 _10662_ (.A(_04014_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand2_1 _10663_ (.A(_04015_),
    .B(\sq.out[19] ),
    .Y(_04016_));
 sky130_fd_sc_hd__nand2_1 _10664_ (.A(_04014_),
    .B(_05140_),
    .Y(_04017_));
 sky130_fd_sc_hd__nand2_1 _10665_ (.A(_04016_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__or2_1 _10666_ (.A(_04018_),
    .B(_03997_),
    .X(_04019_));
 sky130_fd_sc_hd__nand2_1 _10667_ (.A(_03997_),
    .B(_04018_),
    .Y(_04020_));
 sky130_fd_sc_hd__nand2_1 _10668_ (.A(_04019_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__nor2_1 _10669_ (.A(_04021_),
    .B(_04003_),
    .Y(_04022_));
 sky130_fd_sc_hd__inv_2 _10670_ (.A(_04022_),
    .Y(_04024_));
 sky130_fd_sc_hd__nor2_4 _10671_ (.A(_04024_),
    .B(_03989_),
    .Y(_04025_));
 sky130_fd_sc_hd__inv_2 _10672_ (.A(_03720_),
    .Y(_04026_));
 sky130_fd_sc_hd__or2_1 _10673_ (.A(_03697_),
    .B(_03708_),
    .X(_04027_));
 sky130_fd_sc_hd__a21oi_2 _10674_ (.A1(_03662_),
    .A2(_03769_),
    .B1(_03780_),
    .Y(_04028_));
 sky130_fd_sc_hd__o21bai_1 _10675_ (.A1(_04027_),
    .A2(_04028_),
    .B1_N(_03781_),
    .Y(_04029_));
 sky130_fd_sc_hd__a21oi_1 _10676_ (.A1(_04026_),
    .A2(_04029_),
    .B1(_03843_),
    .Y(_04030_));
 sky130_fd_sc_hd__or2_1 _10677_ (.A(_04026_),
    .B(_04029_),
    .X(_04031_));
 sky130_fd_sc_hd__a22o_1 _10678_ (.A1(_03717_),
    .A2(_03843_),
    .B1(_04030_),
    .B2(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__o21ai_1 _10679_ (.A1(_03708_),
    .A2(_04028_),
    .B1(_03706_),
    .Y(_04033_));
 sky130_fd_sc_hd__xor2_1 _10680_ (.A(_03697_),
    .B(_04033_),
    .X(_04035_));
 sky130_fd_sc_hd__nand2_1 _10681_ (.A(_03843_),
    .B(_03695_),
    .Y(_04036_));
 sky130_fd_sc_hd__o21ai_2 _10682_ (.A1(_03843_),
    .A2(_04035_),
    .B1(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__or2_1 _10683_ (.A(_03708_),
    .B(_04028_),
    .X(_04038_));
 sky130_fd_sc_hd__nand2_1 _10684_ (.A(_04028_),
    .B(_03708_),
    .Y(_04039_));
 sky130_fd_sc_hd__nor2_1 _10685_ (.A(_03688_),
    .B(_03822_),
    .Y(_04040_));
 sky130_fd_sc_hd__a31o_2 _10686_ (.A1(_03822_),
    .A2(_04038_),
    .A3(_04039_),
    .B1(_04040_),
    .X(_04041_));
 sky130_fd_sc_hd__or2_1 _10687_ (.A(_04037_),
    .B(_04041_),
    .X(_04042_));
 sky130_fd_sc_hd__nand2_1 _10688_ (.A(_04041_),
    .B(_04037_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand2_1 _10689_ (.A(_04042_),
    .B(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__or2_1 _10690_ (.A(_04032_),
    .B(_04044_),
    .X(_04046_));
 sky130_fd_sc_hd__or2_1 _10691_ (.A(_03775_),
    .B(_03662_),
    .X(_04047_));
 sky130_fd_sc_hd__a21o_1 _10692_ (.A1(_04047_),
    .A2(_03767_),
    .B1(_03777_),
    .X(_04048_));
 sky130_fd_sc_hd__a21bo_1 _10693_ (.A1(_04048_),
    .A2(_03742_),
    .B1_N(_03741_),
    .X(_04049_));
 sky130_fd_sc_hd__xor2_1 _10694_ (.A(_03748_),
    .B(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__nand2_1 _10695_ (.A(_04050_),
    .B(_03822_),
    .Y(_04051_));
 sky130_fd_sc_hd__o21ai_2 _10696_ (.A1(_03703_),
    .A2(\sq.out[3] ),
    .B1(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__nand2_1 _10697_ (.A(_04052_),
    .B(\sq.out[24] ),
    .Y(_04053_));
 sky130_fd_sc_hd__nand2b_1 _10698_ (.A_N(_04053_),
    .B(_04041_),
    .Y(_04054_));
 sky130_fd_sc_hd__a21o_1 _10699_ (.A1(_04052_),
    .A2(\sq.out[24] ),
    .B1(_04041_),
    .X(_04055_));
 sky130_fd_sc_hd__nand2_1 _10700_ (.A(_04054_),
    .B(_04055_),
    .Y(_04057_));
 sky130_fd_sc_hd__xor2_1 _10701_ (.A(_03743_),
    .B(_04048_),
    .X(_04058_));
 sky130_fd_sc_hd__or2_1 _10702_ (.A(_03833_),
    .B(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__nand2_1 _10703_ (.A(net95),
    .B(_03732_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _10704_ (.A(_04059_),
    .B(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__inv_2 _10705_ (.A(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__nand2_1 _10706_ (.A(_04062_),
    .B(\sq.out[23] ),
    .Y(_04063_));
 sky130_fd_sc_hd__or2_1 _10707_ (.A(\sq.out[24] ),
    .B(_04052_),
    .X(_04064_));
 sky130_fd_sc_hd__nand2_1 _10708_ (.A(_04064_),
    .B(_04053_),
    .Y(_04065_));
 sky130_fd_sc_hd__or2_1 _10709_ (.A(_04063_),
    .B(_04065_),
    .X(_04066_));
 sky130_fd_sc_hd__nand2_1 _10710_ (.A(_04065_),
    .B(_04063_),
    .Y(_04068_));
 sky130_fd_sc_hd__nand2_1 _10711_ (.A(_04066_),
    .B(_04068_),
    .Y(_04069_));
 sky130_fd_sc_hd__nor2_1 _10712_ (.A(_04057_),
    .B(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__nor2b_1 _10713_ (.A(_04046_),
    .B_N(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__o2111a_1 _10714_ (.A1(_03722_),
    .A2(_04028_),
    .B1(_03783_),
    .C1(_03784_),
    .D1(_03821_),
    .X(_04072_));
 sky130_fd_sc_hd__nand2b_1 _10715_ (.A_N(_03677_),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__nor2_1 _10716_ (.A(_03673_),
    .B(_04073_),
    .Y(_04074_));
 sky130_fd_sc_hd__or2_1 _10717_ (.A(_03671_),
    .B(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__nand2_1 _10718_ (.A(_04074_),
    .B(_03671_),
    .Y(_04076_));
 sky130_fd_sc_hd__and2_1 _10719_ (.A(_04075_),
    .B(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_04073_),
    .B(_03673_),
    .Y(_04079_));
 sky130_fd_sc_hd__and2b_1 _10721_ (.A_N(_04074_),
    .B(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__nand2_1 _10722_ (.A(_04030_),
    .B(_03719_),
    .Y(_04081_));
 sky130_fd_sc_hd__xnor2_1 _10723_ (.A(_03712_),
    .B(_04081_),
    .Y(_04082_));
 sky130_fd_sc_hd__or2b_1 _10724_ (.A(_04072_),
    .B_N(_03677_),
    .X(_04083_));
 sky130_fd_sc_hd__nand2_1 _10725_ (.A(_04083_),
    .B(_04073_),
    .Y(_04084_));
 sky130_fd_sc_hd__nor2_1 _10726_ (.A(_04082_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__and3_1 _10727_ (.A(_04077_),
    .B(_04080_),
    .C(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__nand2_1 _10728_ (.A(_04071_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__clkinvlp_2 _10729_ (.A(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__xor2_1 _10730_ (.A(_03766_),
    .B(_04047_),
    .X(_04090_));
 sky130_fd_sc_hd__or2_1 _10731_ (.A(_04090_),
    .B(net95),
    .X(_04091_));
 sky130_fd_sc_hd__nand2_1 _10732_ (.A(net95),
    .B(_03754_),
    .Y(_04092_));
 sky130_fd_sc_hd__nand2_1 _10733_ (.A(_04091_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__inv_2 _10734_ (.A(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2_1 _10735_ (.A(_04094_),
    .B(\sq.out[21] ),
    .Y(_04095_));
 sky130_fd_sc_hd__a21bo_1 _10736_ (.A1(_04047_),
    .A2(_03764_),
    .B1_N(_03765_),
    .X(_04096_));
 sky130_fd_sc_hd__xor2_1 _10737_ (.A(_03761_),
    .B(_04096_),
    .X(_04097_));
 sky130_fd_sc_hd__nand2_1 _10738_ (.A(_04097_),
    .B(_03822_),
    .Y(_04098_));
 sky130_fd_sc_hd__o21ai_2 _10739_ (.A1(_03739_),
    .A2(_03822_),
    .B1(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__inv_2 _10740_ (.A(_04099_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_1 _10741_ (.A(_04101_),
    .B(_02009_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand2_1 _10742_ (.A(_04099_),
    .B(\sq.out[22] ),
    .Y(_04103_));
 sky130_fd_sc_hd__nand2_1 _10743_ (.A(_04102_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__or2_1 _10744_ (.A(_04095_),
    .B(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__nand2_1 _10745_ (.A(_04104_),
    .B(_04095_),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_1 _10746_ (.A(_04105_),
    .B(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _10747_ (.A(_04061_),
    .B(_01993_),
    .Y(_04108_));
 sky130_fd_sc_hd__nand2_1 _10748_ (.A(_04063_),
    .B(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__or2_1 _10749_ (.A(_04103_),
    .B(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__nand2_1 _10750_ (.A(_04109_),
    .B(_04103_),
    .Y(_04112_));
 sky130_fd_sc_hd__nand2_1 _10751_ (.A(_04110_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__nor2_1 _10752_ (.A(_04107_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__a21bo_1 _10753_ (.A1(_04009_),
    .A2(_03625_),
    .B1_N(_03626_),
    .X(_04115_));
 sky130_fd_sc_hd__xor2_1 _10754_ (.A(_03615_),
    .B(_04115_),
    .X(_04116_));
 sky130_fd_sc_hd__nand2_1 _10755_ (.A(_03822_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__o21ai_2 _10756_ (.A1(_03609_),
    .A2(_03822_),
    .B1(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__inv_2 _10757_ (.A(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _10758_ (.A(_04119_),
    .B(_01730_),
    .Y(_04120_));
 sky130_fd_sc_hd__nand2_1 _10759_ (.A(_04118_),
    .B(\sq.out[20] ),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _10760_ (.A(_04120_),
    .B(_04121_),
    .Y(_04123_));
 sky130_fd_sc_hd__or2_1 _10761_ (.A(_04016_),
    .B(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__nand2_1 _10762_ (.A(_04123_),
    .B(_04016_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _10763_ (.A(_04124_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_1 _10764_ (.A(_04093_),
    .B(_02927_),
    .Y(_04127_));
 sky130_fd_sc_hd__nand2_1 _10765_ (.A(_04095_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__or2_1 _10766_ (.A(_04121_),
    .B(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__nand2_1 _10767_ (.A(_04128_),
    .B(_04121_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _10768_ (.A(_04129_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__nor2_1 _10769_ (.A(_04126_),
    .B(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__nand2_1 _10770_ (.A(_04114_),
    .B(_04132_),
    .Y(_04134_));
 sky130_fd_sc_hd__inv_4 _10771_ (.A(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand3_4 _10772_ (.A(_04025_),
    .B(_04088_),
    .C(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hd__o21ai_1 _10773_ (.A1(_04002_),
    .A2(_04021_),
    .B1(_04020_),
    .Y(_04137_));
 sky130_fd_sc_hd__a21o_1 _10774_ (.A1(_03853_),
    .A2(_04022_),
    .B1(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__o21ai_1 _10775_ (.A1(_04125_),
    .A2(_04131_),
    .B1(_04130_),
    .Y(_04139_));
 sky130_fd_sc_hd__o21ai_1 _10776_ (.A1(_04106_),
    .A2(_04113_),
    .B1(_04112_),
    .Y(_04140_));
 sky130_fd_sc_hd__a21o_1 _10777_ (.A1(_04114_),
    .A2(_04139_),
    .B1(_04140_),
    .X(_04141_));
 sky130_fd_sc_hd__a21oi_2 _10778_ (.A1(_04138_),
    .A2(_04135_),
    .B1(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__o21a_1 _10779_ (.A1(_04057_),
    .A2(_04068_),
    .B1(_04055_),
    .X(_04143_));
 sky130_fd_sc_hd__a21oi_1 _10780_ (.A1(_04041_),
    .A2(_04037_),
    .B1(_04032_),
    .Y(_04145_));
 sky130_fd_sc_hd__o21ai_1 _10781_ (.A1(_04046_),
    .A2(_04143_),
    .B1(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__or2b_1 _10782_ (.A(_04146_),
    .B_N(_04086_),
    .X(_04147_));
 sky130_fd_sc_hd__o21ba_4 _10783_ (.A1(_04087_),
    .A2(_04142_),
    .B1_N(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__and3_1 _10784_ (.A(_03821_),
    .B(_03770_),
    .C(_03786_),
    .X(_04149_));
 sky130_fd_sc_hd__nand2_1 _10785_ (.A(_04149_),
    .B(_03809_),
    .Y(_04150_));
 sky130_fd_sc_hd__nor2_1 _10786_ (.A(_03795_),
    .B(_04150_),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_1 _10787_ (.A(_04151_),
    .B(_03797_),
    .Y(_04152_));
 sky130_fd_sc_hd__or2_1 _10788_ (.A(_03790_),
    .B(_04152_),
    .X(_04153_));
 sky130_fd_sc_hd__nand2_1 _10789_ (.A(_04152_),
    .B(_03790_),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _10790_ (.A(_04153_),
    .B(_04154_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_1 _10791_ (.A(_04149_),
    .B(_03808_),
    .Y(_04157_));
 sky130_fd_sc_hd__nor2_1 _10792_ (.A(_03805_),
    .B(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__nor2_1 _10793_ (.A(_03807_),
    .B(_04157_),
    .Y(_04159_));
 sky130_fd_sc_hd__o21bai_2 _10794_ (.A1(_03802_),
    .A2(_04158_),
    .B1_N(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__or2_1 _10795_ (.A(_03808_),
    .B(_04149_),
    .X(_04161_));
 sky130_fd_sc_hd__nand2_1 _10796_ (.A(_04161_),
    .B(_04157_),
    .Y(_04162_));
 sky130_fd_sc_hd__nand2_1 _10797_ (.A(_04157_),
    .B(_03805_),
    .Y(_04163_));
 sky130_fd_sc_hd__nor2b_1 _10798_ (.A(_04158_),
    .B_N(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2b_1 _10799_ (.A_N(_04162_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__xor2_2 _10800_ (.A(_03669_),
    .B(_04076_),
    .X(_04167_));
 sky130_fd_sc_hd__nor3_1 _10801_ (.A(_04160_),
    .B(_04165_),
    .C(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__xor2_1 _10802_ (.A(_03800_),
    .B(_04159_),
    .X(_04169_));
 sky130_fd_sc_hd__or2_1 _10803_ (.A(_03797_),
    .B(_04151_),
    .X(_04170_));
 sky130_fd_sc_hd__and2_1 _10804_ (.A(_04170_),
    .B(_04152_),
    .X(_04171_));
 sky130_fd_sc_hd__nand2_1 _10805_ (.A(_04150_),
    .B(_03795_),
    .Y(_04172_));
 sky130_fd_sc_hd__and2b_1 _10806_ (.A_N(_04151_),
    .B(_04172_),
    .X(_04173_));
 sky130_fd_sc_hd__and3b_1 _10807_ (.A_N(_04169_),
    .B(_04171_),
    .C(_04173_),
    .X(_04174_));
 sky130_fd_sc_hd__and3b_1 _10808_ (.A_N(_04156_),
    .B(_04168_),
    .C(_04174_),
    .X(_04175_));
 sky130_fd_sc_hd__nand2_1 _10809_ (.A(\sq.out[3] ),
    .B(_03830_),
    .Y(_04176_));
 sky130_fd_sc_hd__or2_1 _10810_ (.A(_03591_),
    .B(_04176_),
    .X(_04178_));
 sky130_fd_sc_hd__nand2_1 _10811_ (.A(_04176_),
    .B(_03591_),
    .Y(_04179_));
 sky130_fd_sc_hd__nand2_1 _10812_ (.A(_04178_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__nand2_1 _10813_ (.A(\sq.out[3] ),
    .B(_03854_),
    .Y(_04181_));
 sky130_fd_sc_hd__nor2_1 _10814_ (.A(_03585_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand2_1 _10815_ (.A(_04182_),
    .B(_03577_),
    .Y(_04183_));
 sky130_fd_sc_hd__or2_1 _10816_ (.A(_03574_),
    .B(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__xor2_1 _10817_ (.A(_03571_),
    .B(_04184_),
    .X(_04185_));
 sky130_fd_sc_hd__nand2_1 _10818_ (.A(_04178_),
    .B(_03590_),
    .Y(_04186_));
 sky130_fd_sc_hd__nand2_1 _10819_ (.A(\sq.out[3] ),
    .B(_03812_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand2_1 _10820_ (.A(_04186_),
    .B(_04187_),
    .Y(_04189_));
 sky130_fd_sc_hd__clkinvlp_2 _10821_ (.A(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__and3b_1 _10822_ (.A_N(_04180_),
    .B(_04185_),
    .C(_04190_),
    .X(_04191_));
 sky130_fd_sc_hd__xor2_2 _10823_ (.A(_03788_),
    .B(_04153_),
    .X(_04192_));
 sky130_fd_sc_hd__xor2_1 _10824_ (.A(_03817_),
    .B(_04187_),
    .X(_04193_));
 sky130_fd_sc_hd__inv_2 _10825_ (.A(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__or2_1 _10826_ (.A(_03577_),
    .B(_04182_),
    .X(_04195_));
 sky130_fd_sc_hd__nand2_1 _10827_ (.A(_04181_),
    .B(_03585_),
    .Y(_04196_));
 sky130_fd_sc_hd__and2b_1 _10828_ (.A_N(_04182_),
    .B(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__and4_1 _10829_ (.A(_04195_),
    .B(_04197_),
    .C(_03575_),
    .D(_04183_),
    .X(_04198_));
 sky130_fd_sc_hd__and4_1 _10830_ (.A(_04191_),
    .B(_04192_),
    .C(_04194_),
    .D(_04198_),
    .X(_04200_));
 sky130_fd_sc_hd__and2_1 _10831_ (.A(_04175_),
    .B(_04200_),
    .X(_04201_));
 sky130_fd_sc_hd__nand3_4 _10832_ (.A(_04136_),
    .B(_04148_),
    .C(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__nor2_8 _10833_ (.A(_04008_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hd__buf_8 _10834_ (.A(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__nand2_1 _10835_ (.A(net121),
    .B(_03996_),
    .Y(_04205_));
 sky130_fd_sc_hd__o21ai_2 _10836_ (.A1(_04006_),
    .A2(net121),
    .B1(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__or2_1 _10837_ (.A(_05140_),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__nand2_1 _10838_ (.A(_04206_),
    .B(_05140_),
    .Y(_04208_));
 sky130_fd_sc_hd__nand2_1 _10839_ (.A(_04207_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__inv_2 _10840_ (.A(_04202_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2_4 _10841_ (.A(_04211_),
    .B(_04007_),
    .Y(_04212_));
 sky130_fd_sc_hd__buf_6 _10842_ (.A(_04212_),
    .X(\sq.out[2] ));
 sky130_fd_sc_hd__and2_1 _10843_ (.A(_03984_),
    .B(_03988_),
    .X(_04213_));
 sky130_fd_sc_hd__nand2b_1 _10844_ (.A_N(_04213_),
    .B(_03839_),
    .Y(_04214_));
 sky130_fd_sc_hd__or2_1 _10845_ (.A(_03985_),
    .B(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__nand2_1 _10846_ (.A(_04214_),
    .B(_03985_),
    .Y(_04216_));
 sky130_fd_sc_hd__buf_8 _10847_ (.A(_04203_),
    .X(_04217_));
 sky130_fd_sc_hd__a21o_1 _10848_ (.A1(_04215_),
    .A2(_04216_),
    .B1(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__o21ai_2 _10849_ (.A1(_03845_),
    .A2(\sq.out[2] ),
    .B1(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__or2_1 _10850_ (.A(\sq.out[18] ),
    .B(_04219_),
    .X(_04221_));
 sky130_fd_sc_hd__nand2_1 _10851_ (.A(_04219_),
    .B(\sq.out[18] ),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_1 _10852_ (.A(_04221_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__nor2_1 _10853_ (.A(_04209_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__clkinvlp_2 _10854_ (.A(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__xnor2_1 _10855_ (.A(_03905_),
    .B(_03882_),
    .Y(_04226_));
 sky130_fd_sc_hd__nand2_1 _10856_ (.A(_04204_),
    .B(_03894_),
    .Y(_04227_));
 sky130_fd_sc_hd__o21ai_2 _10857_ (.A1(_04226_),
    .A2(_04204_),
    .B1(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__nor2_1 _10858_ (.A(_02495_),
    .B(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _10859_ (.A(_04228_),
    .B(_02495_),
    .Y(_04230_));
 sky130_fd_sc_hd__or2b_1 _10860_ (.A(_04229_),
    .B_N(_04230_),
    .X(_04232_));
 sky130_fd_sc_hd__o21ai_1 _10861_ (.A1(_04008_),
    .A2(_04202_),
    .B1(\sq.out[3] ),
    .Y(_04233_));
 sky130_fd_sc_hd__nand2_1 _10862_ (.A(_04233_),
    .B(_03439_),
    .Y(_04234_));
 sky130_fd_sc_hd__nand2_1 _10863_ (.A(_04234_),
    .B(\sq.out[5] ),
    .Y(_04235_));
 sky130_fd_sc_hd__buf_6 _10864_ (.A(_04217_),
    .X(_04236_));
 sky130_fd_sc_hd__nand2_1 _10865_ (.A(_04236_),
    .B(_03843_),
    .Y(_04237_));
 sky130_fd_sc_hd__nand2_1 _10866_ (.A(_04235_),
    .B(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hd__nand3_1 _10867_ (.A(_04204_),
    .B(_03439_),
    .C(_03843_),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_1 _10868_ (.A(_04212_),
    .B(_03861_),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_1 _10869_ (.A(_04239_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__nand2_1 _10870_ (.A(_04241_),
    .B(\sq.out[6] ),
    .Y(_04243_));
 sky130_fd_sc_hd__nand3_2 _10871_ (.A(_04239_),
    .B(_04240_),
    .C(_02898_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_1 _10872_ (.A(_04243_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__or2b_1 _10873_ (.A(_03858_),
    .B_N(_03870_),
    .X(_04246_));
 sky130_fd_sc_hd__xnor2_1 _10874_ (.A(_03862_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__o21bai_1 _10875_ (.A1(_04008_),
    .A2(_04202_),
    .B1_N(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__inv_2 _10876_ (.A(_03864_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_1 _10877_ (.A(_04217_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__nand2_1 _10878_ (.A(_04248_),
    .B(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hd__nand2_1 _10879_ (.A(_04251_),
    .B(_03112_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _10880_ (.A(_04244_),
    .B(_04252_),
    .Y(_04254_));
 sky130_fd_sc_hd__o21bai_1 _10881_ (.A1(_04238_),
    .A2(_04245_),
    .B1_N(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__a21oi_1 _10882_ (.A1(_03878_),
    .A2(_03879_),
    .B1(_03871_),
    .Y(_04256_));
 sky130_fd_sc_hd__and2b_1 _10883_ (.A_N(_04256_),
    .B(_03881_),
    .X(_04257_));
 sky130_fd_sc_hd__nand2_1 _10884_ (.A(_04212_),
    .B(_04257_),
    .Y(_04258_));
 sky130_fd_sc_hd__o21ai_2 _10885_ (.A1(_03874_),
    .A2(_04212_),
    .B1(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__xor2_1 _10886_ (.A(\sq.out[8] ),
    .B(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__inv_2 _10887_ (.A(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__or2_1 _10888_ (.A(_03112_),
    .B(_04251_),
    .X(_04262_));
 sky130_fd_sc_hd__nand3_2 _10889_ (.A(_04255_),
    .B(_04261_),
    .C(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__nor2_2 _10890_ (.A(_04232_),
    .B(_04263_),
    .Y(_04265_));
 sky130_fd_sc_hd__xor2_1 _10891_ (.A(_03948_),
    .B(_03937_),
    .X(_04266_));
 sky130_fd_sc_hd__or2_1 _10892_ (.A(_04266_),
    .B(_04203_),
    .X(_04267_));
 sky130_fd_sc_hd__nand2_1 _10893_ (.A(_04217_),
    .B(_03941_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_1 _10894_ (.A(_04267_),
    .B(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__nand2_1 _10895_ (.A(_04269_),
    .B(_00844_),
    .Y(_04270_));
 sky130_fd_sc_hd__nand3_1 _10896_ (.A(_04267_),
    .B(\sq.out[13] ),
    .C(_04268_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand2_1 _10897_ (.A(_04270_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__inv_2 _10898_ (.A(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__nand2_1 _10899_ (.A(_03908_),
    .B(_03933_),
    .Y(_04274_));
 sky130_fd_sc_hd__nand2_1 _10900_ (.A(_04274_),
    .B(_03931_),
    .Y(_04276_));
 sky130_fd_sc_hd__or2_1 _10901_ (.A(_03927_),
    .B(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__nand2_1 _10902_ (.A(_04276_),
    .B(_03927_),
    .Y(_04278_));
 sky130_fd_sc_hd__nand3_1 _10903_ (.A(_04212_),
    .B(_04277_),
    .C(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand2_1 _10904_ (.A(_04217_),
    .B(_03919_),
    .Y(_04280_));
 sky130_fd_sc_hd__nand2_1 _10905_ (.A(_04279_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2_1 _10906_ (.A(_04281_),
    .B(_02826_),
    .Y(_04282_));
 sky130_fd_sc_hd__nand3_1 _10907_ (.A(_04279_),
    .B(\sq.out[12] ),
    .C(_04280_),
    .Y(_04283_));
 sky130_fd_sc_hd__nand2_1 _10908_ (.A(_04282_),
    .B(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__inv_2 _10909_ (.A(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__nand2_1 _10910_ (.A(_04273_),
    .B(_04285_),
    .Y(_04287_));
 sky130_fd_sc_hd__xor2_1 _10911_ (.A(_03974_),
    .B(_03963_),
    .X(_04288_));
 sky130_fd_sc_hd__or2_1 _10912_ (.A(_04288_),
    .B(_04203_),
    .X(_04289_));
 sky130_fd_sc_hd__nand2_1 _10913_ (.A(_04217_),
    .B(_03967_),
    .Y(_04290_));
 sky130_fd_sc_hd__nand2_1 _10914_ (.A(_04289_),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__nand2_1 _10915_ (.A(_04291_),
    .B(_02843_),
    .Y(_04292_));
 sky130_fd_sc_hd__nand3_1 _10916_ (.A(_04289_),
    .B(\sq.out[15] ),
    .C(_04290_),
    .Y(_04293_));
 sky130_fd_sc_hd__nand2_1 _10917_ (.A(_04292_),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__a21bo_1 _10918_ (.A1(_03937_),
    .A2(_03945_),
    .B1_N(_03947_),
    .X(_04295_));
 sky130_fd_sc_hd__xor2_1 _10919_ (.A(_03959_),
    .B(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__or2_1 _10920_ (.A(_04296_),
    .B(_04203_),
    .X(_04298_));
 sky130_fd_sc_hd__nand2_1 _10921_ (.A(_04217_),
    .B(_03952_),
    .Y(_04299_));
 sky130_fd_sc_hd__nand2_1 _10922_ (.A(_04298_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__nand2_1 _10923_ (.A(_04300_),
    .B(_02856_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand3_1 _10924_ (.A(_04298_),
    .B(\sq.out[14] ),
    .C(_04299_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_1 _10925_ (.A(_04301_),
    .B(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__nor2_1 _10926_ (.A(_04294_),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__inv_2 _10927_ (.A(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__nor2_1 _10928_ (.A(_04287_),
    .B(_04305_),
    .Y(_04306_));
 sky130_fd_sc_hd__or2_1 _10929_ (.A(_03933_),
    .B(_03908_),
    .X(_04307_));
 sky130_fd_sc_hd__nand3_1 _10930_ (.A(\sq.out[2] ),
    .B(_04274_),
    .C(_04307_),
    .Y(_04309_));
 sky130_fd_sc_hd__nand2_1 _10931_ (.A(_04204_),
    .B(_03912_),
    .Y(_04310_));
 sky130_fd_sc_hd__nand2_1 _10932_ (.A(_04309_),
    .B(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand2_1 _10933_ (.A(_04311_),
    .B(_02345_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand3_1 _10934_ (.A(_04309_),
    .B(\sq.out[11] ),
    .C(_04310_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _10935_ (.A(_04312_),
    .B(_04313_),
    .Y(_04314_));
 sky130_fd_sc_hd__a21bo_1 _10936_ (.A1(_03882_),
    .A2(_03905_),
    .B1_N(_03904_),
    .X(_04315_));
 sky130_fd_sc_hd__or2_1 _10937_ (.A(_03899_),
    .B(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__nand2_1 _10938_ (.A(_04315_),
    .B(_03899_),
    .Y(_04317_));
 sky130_fd_sc_hd__nand3_1 _10939_ (.A(\sq.out[2] ),
    .B(_04316_),
    .C(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__nand2_1 _10940_ (.A(_04204_),
    .B(_03886_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand2_1 _10941_ (.A(_04318_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__nand2_1 _10942_ (.A(_04321_),
    .B(_02504_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand3_1 _10943_ (.A(_04318_),
    .B(\sq.out[10] ),
    .C(_04320_),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2_1 _10944_ (.A(_04322_),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hd__nor2_1 _10945_ (.A(_04314_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__nand3_1 _10946_ (.A(_04265_),
    .B(_04306_),
    .C(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand2_1 _10947_ (.A(_04259_),
    .B(_02498_),
    .Y(_04327_));
 sky130_fd_sc_hd__o21ai_1 _10948_ (.A1(_04229_),
    .A2(_04327_),
    .B1(_04230_),
    .Y(_04328_));
 sky130_fd_sc_hd__nand2_1 _10949_ (.A(_04328_),
    .B(_04325_),
    .Y(_04329_));
 sky130_fd_sc_hd__and2_1 _10950_ (.A(_04321_),
    .B(_02504_),
    .X(_04331_));
 sky130_fd_sc_hd__a21boi_1 _10951_ (.A1(_04331_),
    .A2(_04313_),
    .B1_N(_04312_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand2_1 _10952_ (.A(_04329_),
    .B(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__o21a_1 _10953_ (.A1(_04301_),
    .A2(_04294_),
    .B1(_04292_),
    .X(_04334_));
 sky130_fd_sc_hd__inv_2 _10954_ (.A(_04271_),
    .Y(_04335_));
 sky130_fd_sc_hd__o21ai_1 _10955_ (.A1(_04282_),
    .A2(_04335_),
    .B1(_04270_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _10956_ (.A(_04336_),
    .B(_04304_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_1 _10957_ (.A(_04334_),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__a21oi_1 _10958_ (.A1(_04306_),
    .A2(_04333_),
    .B1(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__nand2_1 _10959_ (.A(_04326_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__or2_1 _10960_ (.A(_03988_),
    .B(_03984_),
    .X(_04342_));
 sky130_fd_sc_hd__or2b_1 _10961_ (.A(_04213_),
    .B_N(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__nand2_1 _10962_ (.A(_04236_),
    .B(_03823_),
    .Y(_04344_));
 sky130_fd_sc_hd__o21ai_2 _10963_ (.A1(_04343_),
    .A2(_04236_),
    .B1(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__or2_1 _10964_ (.A(_02877_),
    .B(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__nand2_1 _10965_ (.A(_04345_),
    .B(_02877_),
    .Y(_04347_));
 sky130_fd_sc_hd__nand2_1 _10966_ (.A(_04346_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hd__clkinvlp_2 _10967_ (.A(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__a21bo_1 _10968_ (.A1(_03963_),
    .A2(_03972_),
    .B1_N(_03973_),
    .X(_04350_));
 sky130_fd_sc_hd__xnor2_1 _10969_ (.A(_03980_),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(_04351_),
    .A1(_03836_),
    .S(_04217_),
    .X(_04353_));
 sky130_fd_sc_hd__or2_1 _10971_ (.A(_00092_),
    .B(_04353_),
    .X(_04354_));
 sky130_fd_sc_hd__nand2_1 _10972_ (.A(_04353_),
    .B(_00092_),
    .Y(_04355_));
 sky130_fd_sc_hd__nand2_1 _10973_ (.A(_04354_),
    .B(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__inv_2 _10974_ (.A(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__nand3_2 _10975_ (.A(_04340_),
    .B(_04349_),
    .C(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__nor2_4 _10976_ (.A(_04225_),
    .B(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__a21bo_1 _10977_ (.A1(_04025_),
    .A2(_04135_),
    .B1_N(_04142_),
    .X(_04360_));
 sky130_fd_sc_hd__or2b_1 _10978_ (.A(_04360_),
    .B_N(_04069_),
    .X(_04361_));
 sky130_fd_sc_hd__or2b_1 _10979_ (.A(_04069_),
    .B_N(_04360_),
    .X(_04362_));
 sky130_fd_sc_hd__nand2_1 _10980_ (.A(_04361_),
    .B(_04362_),
    .Y(_04364_));
 sky130_fd_sc_hd__mux2_1 _10981_ (.A0(_04364_),
    .A1(_04052_),
    .S(_04236_),
    .X(_04365_));
 sky130_fd_sc_hd__inv_2 _10982_ (.A(_04132_),
    .Y(_04366_));
 sky130_fd_sc_hd__nor2_1 _10983_ (.A(_04138_),
    .B(_04025_),
    .Y(_04367_));
 sky130_fd_sc_hd__o21bai_1 _10984_ (.A1(_04366_),
    .A2(_04367_),
    .B1_N(_04139_),
    .Y(_04368_));
 sky130_fd_sc_hd__nand2b_1 _10985_ (.A_N(_04107_),
    .B(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__nand2_1 _10986_ (.A(_04369_),
    .B(_04106_),
    .Y(_04370_));
 sky130_fd_sc_hd__xor2_1 _10987_ (.A(_04113_),
    .B(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__nand2_1 _10988_ (.A(_04371_),
    .B(\sq.out[2] ),
    .Y(_04372_));
 sky130_fd_sc_hd__nand2_1 _10989_ (.A(net121),
    .B(_04062_),
    .Y(_04373_));
 sky130_fd_sc_hd__nand2_2 _10990_ (.A(_04372_),
    .B(_04373_),
    .Y(_04375_));
 sky130_fd_sc_hd__inv_2 _10991_ (.A(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand2_1 _10992_ (.A(_04376_),
    .B(_01081_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(_04375_),
    .B(\sq.out[24] ),
    .Y(_04378_));
 sky130_fd_sc_hd__nand2_1 _10994_ (.A(_04377_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__or2_1 _10995_ (.A(_04365_),
    .B(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__a21oi_1 _10996_ (.A1(_04360_),
    .A2(_04071_),
    .B1(_04146_),
    .Y(_04381_));
 sky130_fd_sc_hd__nand2_1 _10997_ (.A(_04381_),
    .B(_04212_),
    .Y(_04382_));
 sky130_fd_sc_hd__inv_2 _10998_ (.A(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__or2_1 _10999_ (.A(_04082_),
    .B(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__nand2_1 _11000_ (.A(_04383_),
    .B(_04082_),
    .Y(_04386_));
 sky130_fd_sc_hd__a21o_1 _11001_ (.A1(_04384_),
    .A2(_04386_),
    .B1(_04084_),
    .X(_04387_));
 sky130_fd_sc_hd__a21bo_1 _11002_ (.A1(_04360_),
    .A2(_04070_),
    .B1_N(_04143_),
    .X(_04388_));
 sky130_fd_sc_hd__inv_2 _11003_ (.A(_04044_),
    .Y(_04389_));
 sky130_fd_sc_hd__nand2_1 _11004_ (.A(_04388_),
    .B(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand3_1 _11005_ (.A(_04390_),
    .B(_04043_),
    .C(\sq.out[2] ),
    .Y(_04391_));
 sky130_fd_sc_hd__xor2_1 _11006_ (.A(_04032_),
    .B(_04391_),
    .X(_04392_));
 sky130_fd_sc_hd__nor2b_1 _11007_ (.A(_04387_),
    .B_N(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__a31o_1 _11008_ (.A1(_04381_),
    .A2(\sq.out[2] ),
    .A3(_04085_),
    .B1(_04080_),
    .X(_04394_));
 sky130_fd_sc_hd__nand3_1 _11009_ (.A(_04383_),
    .B(_04080_),
    .C(_04085_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2_1 _11010_ (.A(_04394_),
    .B(_04395_),
    .Y(_04397_));
 sky130_fd_sc_hd__inv_2 _11011_ (.A(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__and2_1 _11012_ (.A(_04393_),
    .B(_04398_),
    .X(_04399_));
 sky130_fd_sc_hd__or2_1 _11013_ (.A(_04389_),
    .B(_04388_),
    .X(_04400_));
 sky130_fd_sc_hd__and2_1 _11014_ (.A(_04236_),
    .B(_04037_),
    .X(_04401_));
 sky130_fd_sc_hd__a31o_1 _11015_ (.A1(_04400_),
    .A2(\sq.out[2] ),
    .A3(_04390_),
    .B1(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__inv_2 _11016_ (.A(_04057_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_1 _11017_ (.A(_04362_),
    .B(_04068_),
    .Y(_04404_));
 sky130_fd_sc_hd__o21ai_1 _11018_ (.A1(_04403_),
    .A2(_04404_),
    .B1(\sq.out[2] ),
    .Y(_04405_));
 sky130_fd_sc_hd__a21oi_1 _11019_ (.A1(_04403_),
    .A2(_04404_),
    .B1(_04405_),
    .Y(_04406_));
 sky130_fd_sc_hd__a21o_1 _11020_ (.A1(_04041_),
    .A2(_04236_),
    .B1(_04406_),
    .X(_04408_));
 sky130_fd_sc_hd__nor2_1 _11021_ (.A(_04402_),
    .B(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__nand2_1 _11022_ (.A(_04399_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nor2_1 _11023_ (.A(_04380_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__xnor2_1 _11024_ (.A(_04126_),
    .B(_04367_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand2_1 _11025_ (.A(_04236_),
    .B(_04119_),
    .Y(_04413_));
 sky130_fd_sc_hd__o21ai_2 _11026_ (.A1(_04412_),
    .A2(_04236_),
    .B1(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__or2_1 _11027_ (.A(_02927_),
    .B(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__nand2_1 _11028_ (.A(_04414_),
    .B(_02927_),
    .Y(_04416_));
 sky130_fd_sc_hd__nand2_1 _11029_ (.A(_04415_),
    .B(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__nand2_1 _11030_ (.A(_04005_),
    .B(_04002_),
    .Y(_04419_));
 sky130_fd_sc_hd__xor2_1 _11031_ (.A(_04021_),
    .B(_04419_),
    .X(_04420_));
 sky130_fd_sc_hd__mux2_4 _11032_ (.A0(_04420_),
    .A1(_04015_),
    .S(_04217_),
    .X(_04421_));
 sky130_fd_sc_hd__or2_1 _11033_ (.A(\sq.out[20] ),
    .B(_04421_),
    .X(_04422_));
 sky130_fd_sc_hd__nand2_1 _11034_ (.A(_04421_),
    .B(\sq.out[20] ),
    .Y(_04423_));
 sky130_fd_sc_hd__nand2_1 _11035_ (.A(_04422_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__nor2_1 _11036_ (.A(_04417_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hd__o21ai_1 _11037_ (.A1(_04126_),
    .A2(_04367_),
    .B1(_04125_),
    .Y(_04426_));
 sky130_fd_sc_hd__xor2_1 _11038_ (.A(_04131_),
    .B(_04426_),
    .X(_04427_));
 sky130_fd_sc_hd__nand2_1 _11039_ (.A(_04427_),
    .B(_04212_),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_1 _11040_ (.A(_04217_),
    .B(_04094_),
    .Y(_04430_));
 sky130_fd_sc_hd__nand2_1 _11041_ (.A(_04428_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__inv_2 _11042_ (.A(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__nand2_1 _11043_ (.A(_04432_),
    .B(_02009_),
    .Y(_04433_));
 sky130_fd_sc_hd__nand2_1 _11044_ (.A(_04431_),
    .B(\sq.out[22] ),
    .Y(_04434_));
 sky130_fd_sc_hd__nand2_1 _11045_ (.A(_04433_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__or2b_1 _11046_ (.A(_04368_),
    .B_N(_04107_),
    .X(_04436_));
 sky130_fd_sc_hd__nand2_1 _11047_ (.A(_04436_),
    .B(_04369_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _11048_ (.A(net121),
    .B(_04101_),
    .Y(_04438_));
 sky130_fd_sc_hd__o21ai_2 _11049_ (.A1(net121),
    .A2(_04437_),
    .B1(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__inv_2 _11050_ (.A(_04439_),
    .Y(_04441_));
 sky130_fd_sc_hd__nand2_1 _11051_ (.A(_04441_),
    .B(\sq.out[23] ),
    .Y(_04442_));
 sky130_fd_sc_hd__nand2_1 _11052_ (.A(_04439_),
    .B(_01993_),
    .Y(_04443_));
 sky130_fd_sc_hd__nand2_1 _11053_ (.A(_04442_),
    .B(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__nor2_1 _11054_ (.A(_04435_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__and2_4 _11055_ (.A(_04425_),
    .B(_04445_),
    .X(_04446_));
 sky130_fd_sc_hd__nand3_4 _11056_ (.A(_04359_),
    .B(_04411_),
    .C(_04446_),
    .Y(_04447_));
 sky130_fd_sc_hd__o21ai_1 _11057_ (.A1(_04348_),
    .A2(_04355_),
    .B1(_04347_),
    .Y(_04448_));
 sky130_fd_sc_hd__o21ai_1 _11058_ (.A1(_04209_),
    .A2(_04221_),
    .B1(_04208_),
    .Y(_04449_));
 sky130_fd_sc_hd__a21o_1 _11059_ (.A1(_04448_),
    .A2(_04224_),
    .B1(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__nand2_1 _11060_ (.A(_04446_),
    .B(_04450_),
    .Y(_04452_));
 sky130_fd_sc_hd__o21ai_1 _11061_ (.A1(_04417_),
    .A2(_04422_),
    .B1(_04416_),
    .Y(_04453_));
 sky130_fd_sc_hd__o21ai_1 _11062_ (.A1(_04433_),
    .A2(_04444_),
    .B1(_04443_),
    .Y(_04454_));
 sky130_fd_sc_hd__a21oi_1 _11063_ (.A1(_04453_),
    .A2(_04445_),
    .B1(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__nand2_2 _11064_ (.A(_04452_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__o21a_1 _11065_ (.A1(_04365_),
    .A2(_04377_),
    .B1(_04409_),
    .X(_04457_));
 sky130_fd_sc_hd__nand2_1 _11066_ (.A(_04457_),
    .B(_04399_),
    .Y(_04458_));
 sky130_fd_sc_hd__a21oi_4 _11067_ (.A1(_04456_),
    .A2(_04411_),
    .B1(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2_1 _11068_ (.A(_04136_),
    .B(_04148_),
    .Y(_04460_));
 sky130_fd_sc_hd__or2_4 _11069_ (.A(_04460_),
    .B(_04203_),
    .X(_04461_));
 sky130_fd_sc_hd__inv_2 _11070_ (.A(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_1 _11071_ (.A(_04463_),
    .B(_04168_),
    .Y(_04464_));
 sky130_fd_sc_hd__nor2_2 _11072_ (.A(_04169_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__or2_1 _11073_ (.A(_04173_),
    .B(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__nand2_1 _11074_ (.A(_04465_),
    .B(_04173_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _11075_ (.A(_04466_),
    .B(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand2b_2 _11076_ (.A_N(_04467_),
    .B(_04171_),
    .Y(_04469_));
 sky130_fd_sc_hd__a21o_1 _11077_ (.A1(_04465_),
    .A2(_04173_),
    .B1(_04171_),
    .X(_04470_));
 sky130_fd_sc_hd__nand2_1 _11078_ (.A(_04469_),
    .B(_04470_),
    .Y(_04471_));
 sky130_fd_sc_hd__or2_1 _11079_ (.A(_04468_),
    .B(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__xnor2_1 _11080_ (.A(_04077_),
    .B(_04395_),
    .Y(_04474_));
 sky130_fd_sc_hd__inv_4 _11081_ (.A(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__or2_1 _11082_ (.A(_04167_),
    .B(_04461_),
    .X(_04476_));
 sky130_fd_sc_hd__nor2_2 _11083_ (.A(_04162_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__and2_1 _11084_ (.A(_04476_),
    .B(_04162_),
    .X(_04478_));
 sky130_fd_sc_hd__nor2_2 _11085_ (.A(_04477_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__nand2_1 _11086_ (.A(_04461_),
    .B(_04167_),
    .Y(_04480_));
 sky130_fd_sc_hd__nand2_1 _11087_ (.A(_04476_),
    .B(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hd__clkinvlp_2 _11088_ (.A(_04481_),
    .Y(_04482_));
 sky130_fd_sc_hd__nand2_1 _11089_ (.A(_04479_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__or2_1 _11090_ (.A(_04164_),
    .B(_04477_),
    .X(_04485_));
 sky130_fd_sc_hd__nand2_1 _11091_ (.A(_04477_),
    .B(_04164_),
    .Y(_04486_));
 sky130_fd_sc_hd__nand2_1 _11092_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__nor3_2 _11093_ (.A(_04475_),
    .B(_04483_),
    .C(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__and2_1 _11094_ (.A(_04464_),
    .B(_04169_),
    .X(_04489_));
 sky130_fd_sc_hd__or2_1 _11095_ (.A(_04465_),
    .B(_04489_),
    .X(_04490_));
 sky130_fd_sc_hd__xnor2_1 _11096_ (.A(_04160_),
    .B(_04486_),
    .Y(_04491_));
 sky130_fd_sc_hd__nor2_2 _11097_ (.A(_04490_),
    .B(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__nand3b_4 _11098_ (.A_N(_04472_),
    .B(_04488_),
    .C(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hd__and4_1 _11099_ (.A(_04463_),
    .B(_04192_),
    .C(_04198_),
    .D(_04175_),
    .X(_04494_));
 sky130_fd_sc_hd__nand2_1 _11100_ (.A(_04494_),
    .B(_04185_),
    .Y(_04496_));
 sky130_fd_sc_hd__or2_1 _11101_ (.A(_04180_),
    .B(_04496_),
    .X(_04497_));
 sky130_fd_sc_hd__nand2_1 _11102_ (.A(_04496_),
    .B(_04180_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand3_1 _11103_ (.A(_04497_),
    .B(_04190_),
    .C(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__nand2_1 _11104_ (.A(_04183_),
    .B(_03574_),
    .Y(_04500_));
 sky130_fd_sc_hd__nand2_1 _11105_ (.A(_04184_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand2_1 _11106_ (.A(_04463_),
    .B(_04175_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand3b_4 _11107_ (.A_N(_04502_),
    .B(_04192_),
    .C(_04197_),
    .Y(_04503_));
 sky130_fd_sc_hd__and2_1 _11108_ (.A(_04195_),
    .B(_04183_),
    .X(_04504_));
 sky130_fd_sc_hd__or2b_4 _11109_ (.A(_04503_),
    .B_N(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__xor2_4 _11110_ (.A(_04501_),
    .B(_04505_),
    .X(_04507_));
 sky130_fd_sc_hd__or2_1 _11111_ (.A(_04185_),
    .B(_04494_),
    .X(_04508_));
 sky130_fd_sc_hd__nand2_1 _11112_ (.A(_04508_),
    .B(_04496_),
    .Y(_04509_));
 sky130_fd_sc_hd__inv_2 _11113_ (.A(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand2_1 _11114_ (.A(_04507_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_1 _11115_ (.A(_04499_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__xor2_2 _11116_ (.A(_04156_),
    .B(_04469_),
    .X(_04513_));
 sky130_fd_sc_hd__inv_2 _11117_ (.A(_04192_),
    .Y(_04514_));
 sky130_fd_sc_hd__or2_1 _11118_ (.A(_04514_),
    .B(_04502_),
    .X(_04515_));
 sky130_fd_sc_hd__nand2_1 _11119_ (.A(_04502_),
    .B(_04514_),
    .Y(_04516_));
 sky130_fd_sc_hd__and4_1 _11120_ (.A(_04515_),
    .B(_04197_),
    .C(_04504_),
    .D(_04516_),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_2 _11121_ (.A(_04513_),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__inv_4 _11122_ (.A(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _11123_ (.A(_04512_),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__nor2_4 _11124_ (.A(_04493_),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__nand3_4 _11125_ (.A(_04447_),
    .B(_04459_),
    .C(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__inv_2 _11126_ (.A(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__nand2_2 _11127_ (.A(_04494_),
    .B(_04191_),
    .Y(_04525_));
 sky130_fd_sc_hd__xor2_4 _11128_ (.A(_04194_),
    .B(_04525_),
    .X(_04526_));
 sky130_fd_sc_hd__clkinvlp_2 _11129_ (.A(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand2_2 _11130_ (.A(_04202_),
    .B(_04008_),
    .Y(_04529_));
 sky130_fd_sc_hd__nand3_2 _11131_ (.A(_04524_),
    .B(_04527_),
    .C(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__buf_6 _11132_ (.A(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__and2_1 _11133_ (.A(_04233_),
    .B(_04237_),
    .X(_04532_));
 sky130_fd_sc_hd__nand2_1 _11134_ (.A(_04531_),
    .B(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__nor2_4 _11135_ (.A(_04526_),
    .B(_04523_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand3_2 _11136_ (.A(_04534_),
    .B(_04236_),
    .C(_04529_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2_1 _11137_ (.A(_04533_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__nand2_1 _11138_ (.A(_04536_),
    .B(\sq.out[4] ),
    .Y(_04537_));
 sky130_fd_sc_hd__nand3_1 _11139_ (.A(_04533_),
    .B(_03439_),
    .C(_04535_),
    .Y(_04538_));
 sky130_fd_sc_hd__inv_2 _11140_ (.A(_04530_),
    .Y(_04540_));
 sky130_fd_sc_hd__buf_6 _11141_ (.A(_04540_),
    .X(_04541_));
 sky130_fd_sc_hd__nand2_1 _11142_ (.A(_04541_),
    .B(\sq.out[3] ),
    .Y(_04542_));
 sky130_fd_sc_hd__nand3_1 _11143_ (.A(_04537_),
    .B(_04538_),
    .C(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__nand2_1 _11144_ (.A(_04543_),
    .B(_04538_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _11145_ (.A(\sq.out[3] ),
    .B(\sq.out[4] ),
    .Y(_04545_));
 sky130_fd_sc_hd__nand2_1 _11146_ (.A(_03857_),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__nand2_1 _11147_ (.A(_04531_),
    .B(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__nand3_1 _11148_ (.A(_04534_),
    .B(_04237_),
    .C(_04529_),
    .Y(_04548_));
 sky130_fd_sc_hd__nand2_1 _11149_ (.A(_04547_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__nand2_1 _11150_ (.A(_04549_),
    .B(_03373_),
    .Y(_04551_));
 sky130_fd_sc_hd__nand3_1 _11151_ (.A(_04547_),
    .B(\sq.out[5] ),
    .C(_04548_),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_1 _11152_ (.A(_04551_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__inv_2 _11153_ (.A(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hd__nand2_1 _11154_ (.A(_04544_),
    .B(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__nand2_1 _11155_ (.A(_04555_),
    .B(_04551_),
    .Y(_04556_));
 sky130_fd_sc_hd__nand2_1 _11156_ (.A(_04234_),
    .B(_04237_),
    .Y(_04557_));
 sky130_fd_sc_hd__xor2_1 _11157_ (.A(_03373_),
    .B(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__nor2_1 _11158_ (.A(_04546_),
    .B(_04236_),
    .Y(_04559_));
 sky130_fd_sc_hd__o22ai_2 _11159_ (.A1(_04558_),
    .A2(_04541_),
    .B1(_04559_),
    .B2(_04548_),
    .Y(_04560_));
 sky130_fd_sc_hd__or2_1 _11160_ (.A(_02898_),
    .B(_04560_),
    .X(_04562_));
 sky130_fd_sc_hd__nand2_1 _11161_ (.A(_04556_),
    .B(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hd__nand2_1 _11162_ (.A(_04560_),
    .B(_02898_),
    .Y(_04564_));
 sky130_fd_sc_hd__nand2_1 _11163_ (.A(_04563_),
    .B(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__or2_1 _11164_ (.A(_04238_),
    .B(_04245_),
    .X(_04566_));
 sky130_fd_sc_hd__nand2_1 _11165_ (.A(_04245_),
    .B(_04238_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand3_1 _11166_ (.A(_04531_),
    .B(_04566_),
    .C(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__o21ai_1 _11167_ (.A1(_04241_),
    .A2(net101),
    .B1(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__or2_1 _11168_ (.A(_03112_),
    .B(_04569_),
    .X(_04570_));
 sky130_fd_sc_hd__nand2_1 _11169_ (.A(_04569_),
    .B(_03112_),
    .Y(_04571_));
 sky130_fd_sc_hd__nand2_1 _11170_ (.A(_04570_),
    .B(_04571_),
    .Y(_04573_));
 sky130_fd_sc_hd__inv_2 _11171_ (.A(_04573_),
    .Y(_04574_));
 sky130_fd_sc_hd__nand2_1 _11172_ (.A(_04565_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hd__nand2_1 _11173_ (.A(_04566_),
    .B(_04244_),
    .Y(_04576_));
 sky130_fd_sc_hd__a21oi_1 _11174_ (.A1(_04262_),
    .A2(_04252_),
    .B1(_04576_),
    .Y(_04577_));
 sky130_fd_sc_hd__and3_1 _11175_ (.A(_04576_),
    .B(_04262_),
    .C(_04252_),
    .X(_04578_));
 sky130_fd_sc_hd__nand2_1 _11176_ (.A(_04541_),
    .B(_04251_),
    .Y(_04579_));
 sky130_fd_sc_hd__o31ai_2 _11177_ (.A1(_04577_),
    .A2(_04578_),
    .A3(_04541_),
    .B1(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__nand2_1 _11178_ (.A(_04580_),
    .B(_02498_),
    .Y(_04581_));
 sky130_fd_sc_hd__nand2_1 _11179_ (.A(_04581_),
    .B(_04571_),
    .Y(_04582_));
 sky130_fd_sc_hd__inv_2 _11180_ (.A(_04582_),
    .Y(_04584_));
 sky130_fd_sc_hd__nand2_1 _11181_ (.A(_04575_),
    .B(_04584_),
    .Y(_04585_));
 sky130_fd_sc_hd__a21o_1 _11182_ (.A1(_04255_),
    .A2(_04262_),
    .B1(_04261_),
    .X(_04586_));
 sky130_fd_sc_hd__nand2_1 _11183_ (.A(_04586_),
    .B(_04263_),
    .Y(_04587_));
 sky130_fd_sc_hd__nand2_1 _11184_ (.A(_04540_),
    .B(_04259_),
    .Y(_04588_));
 sky130_fd_sc_hd__o21ai_1 _11185_ (.A1(_04587_),
    .A2(_04540_),
    .B1(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__or2_1 _11186_ (.A(_02495_),
    .B(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__nand2_1 _11187_ (.A(_04589_),
    .B(_02495_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand2_1 _11188_ (.A(_04590_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__inv_2 _11189_ (.A(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__o21ai_1 _11190_ (.A1(_02498_),
    .A2(_04580_),
    .B1(_04593_),
    .Y(_04595_));
 sky130_fd_sc_hd__inv_2 _11191_ (.A(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__nand2_1 _11192_ (.A(_04585_),
    .B(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _11193_ (.A(_04597_),
    .B(_04591_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_1 _11194_ (.A(_04263_),
    .B(_04327_),
    .Y(_04599_));
 sky130_fd_sc_hd__xor2_1 _11195_ (.A(_04232_),
    .B(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__buf_6 _11196_ (.A(_04541_),
    .X(_04601_));
 sky130_fd_sc_hd__nand2_1 _11197_ (.A(_04601_),
    .B(_04228_),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_1 _11198_ (.A1(_04600_),
    .A2(_04601_),
    .B1(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__or2_1 _11199_ (.A(_02504_),
    .B(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__nand2_1 _11200_ (.A(_04598_),
    .B(_04604_),
    .Y(_04606_));
 sky130_fd_sc_hd__nand2_1 _11201_ (.A(_04603_),
    .B(_02504_),
    .Y(_04607_));
 sky130_fd_sc_hd__nand2_1 _11202_ (.A(_04606_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__buf_6 _11203_ (.A(_04531_),
    .X(_04609_));
 sky130_fd_sc_hd__or2_1 _11204_ (.A(_04328_),
    .B(_04265_),
    .X(_04610_));
 sky130_fd_sc_hd__or2b_1 _11205_ (.A(_04324_),
    .B_N(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__or2b_1 _11206_ (.A(_04610_),
    .B_N(_04324_),
    .X(_04612_));
 sky130_fd_sc_hd__nand3_1 _11207_ (.A(_04609_),
    .B(_04611_),
    .C(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand2_1 _11208_ (.A(_04601_),
    .B(_04321_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2_1 _11209_ (.A(_04613_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__clkinvlp_2 _11210_ (.A(_04615_),
    .Y(_04617_));
 sky130_fd_sc_hd__nand2_1 _11211_ (.A(_04611_),
    .B(_04322_),
    .Y(_04618_));
 sky130_fd_sc_hd__nand2_1 _11212_ (.A(_04618_),
    .B(_04314_),
    .Y(_04619_));
 sky130_fd_sc_hd__or2_1 _11213_ (.A(_04314_),
    .B(_04618_),
    .X(_04620_));
 sky130_fd_sc_hd__a21o_1 _11214_ (.A1(_04619_),
    .A2(_04620_),
    .B1(_04541_),
    .X(_04621_));
 sky130_fd_sc_hd__nand2_1 _11215_ (.A(_04601_),
    .B(_04311_),
    .Y(_04622_));
 sky130_fd_sc_hd__nand2_1 _11216_ (.A(_04621_),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__or2_1 _11217_ (.A(_02826_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__nand2_1 _11218_ (.A(_04623_),
    .B(_02826_),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_1 _11219_ (.A(_04624_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__nand2_1 _11220_ (.A(_04615_),
    .B(_02345_),
    .Y(_04628_));
 sky130_fd_sc_hd__nand2b_1 _11221_ (.A_N(_04626_),
    .B(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__a21oi_1 _11222_ (.A1(\sq.out[11] ),
    .A2(_04617_),
    .B1(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _11223_ (.A(_04608_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__o21a_1 _11224_ (.A1(_04628_),
    .A2(_04626_),
    .B1(_04625_),
    .X(_04632_));
 sky130_fd_sc_hd__nand2_1 _11225_ (.A(_04631_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__a21o_1 _11226_ (.A1(_04265_),
    .A2(_04325_),
    .B1(_04333_),
    .X(_04634_));
 sky130_fd_sc_hd__nand2_1 _11227_ (.A(_04634_),
    .B(_04285_),
    .Y(_04635_));
 sky130_fd_sc_hd__nand2_1 _11228_ (.A(_04635_),
    .B(_04282_),
    .Y(_04636_));
 sky130_fd_sc_hd__nand2_1 _11229_ (.A(_04636_),
    .B(_04272_),
    .Y(_04637_));
 sky130_fd_sc_hd__or2_1 _11230_ (.A(_04272_),
    .B(_04636_),
    .X(_04639_));
 sky130_fd_sc_hd__a21o_1 _11231_ (.A1(_04637_),
    .A2(_04639_),
    .B1(_04541_),
    .X(_04640_));
 sky130_fd_sc_hd__nand2_1 _11232_ (.A(_04541_),
    .B(_04269_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand2_1 _11233_ (.A(_04640_),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__or2_1 _11234_ (.A(_02856_),
    .B(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__nand2_1 _11235_ (.A(_04642_),
    .B(_02856_),
    .Y(_04644_));
 sky130_fd_sc_hd__nand2_1 _11236_ (.A(_04643_),
    .B(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__or2_1 _11237_ (.A(_04285_),
    .B(_04634_),
    .X(_04646_));
 sky130_fd_sc_hd__and3_1 _11238_ (.A(_04534_),
    .B(_04281_),
    .C(_04529_),
    .X(_04647_));
 sky130_fd_sc_hd__a31o_1 _11239_ (.A1(net101),
    .A2(_04635_),
    .A3(_04646_),
    .B1(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__or2_1 _11240_ (.A(_00844_),
    .B(_04648_),
    .X(_04650_));
 sky130_fd_sc_hd__nand2_1 _11241_ (.A(_04648_),
    .B(_00844_),
    .Y(_04651_));
 sky130_fd_sc_hd__nand2_1 _11242_ (.A(_04650_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__inv_2 _11243_ (.A(_04294_),
    .Y(_04653_));
 sky130_fd_sc_hd__a31o_1 _11244_ (.A1(_04634_),
    .A2(_04273_),
    .A3(_04285_),
    .B1(_04336_),
    .X(_04654_));
 sky130_fd_sc_hd__inv_2 _11245_ (.A(_04303_),
    .Y(_04655_));
 sky130_fd_sc_hd__nand2_1 _11246_ (.A(_04654_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__nand2_1 _11247_ (.A(_04656_),
    .B(_04301_),
    .Y(_04657_));
 sky130_fd_sc_hd__or2_1 _11248_ (.A(_04653_),
    .B(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__nand2_1 _11249_ (.A(_04657_),
    .B(_04653_),
    .Y(_04659_));
 sky130_fd_sc_hd__a21o_1 _11250_ (.A1(_04658_),
    .A2(_04659_),
    .B1(_04541_),
    .X(_04661_));
 sky130_fd_sc_hd__o21ai_2 _11251_ (.A1(_04291_),
    .A2(_04609_),
    .B1(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__or2_1 _11252_ (.A(\sq.out[16] ),
    .B(_04662_),
    .X(_04663_));
 sky130_fd_sc_hd__nand2_1 _11253_ (.A(_04662_),
    .B(\sq.out[16] ),
    .Y(_04664_));
 sky130_fd_sc_hd__nand2_1 _11254_ (.A(_04663_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__buf_8 _11255_ (.A(_04609_),
    .X(\sq.out[1] ));
 sky130_fd_sc_hd__or2_1 _11256_ (.A(_04655_),
    .B(_04654_),
    .X(_04666_));
 sky130_fd_sc_hd__nand3_1 _11257_ (.A(\sq.out[1] ),
    .B(_04656_),
    .C(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__nand2_1 _11258_ (.A(_04601_),
    .B(_04300_),
    .Y(_04668_));
 sky130_fd_sc_hd__nand2_1 _11259_ (.A(_04667_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hd__or2_1 _11260_ (.A(_02843_),
    .B(_04669_),
    .X(_04671_));
 sky130_fd_sc_hd__nand2_1 _11261_ (.A(_04669_),
    .B(_02843_),
    .Y(_04672_));
 sky130_fd_sc_hd__nand3b_1 _11262_ (.A_N(_04665_),
    .B(_04671_),
    .C(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__nor3_1 _11263_ (.A(_04645_),
    .B(_04652_),
    .C(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_1 _11264_ (.A(_04633_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__or2_1 _11265_ (.A(_04651_),
    .B(_04645_),
    .X(_04676_));
 sky130_fd_sc_hd__nand2_1 _11266_ (.A(_04676_),
    .B(_04644_),
    .Y(_04677_));
 sky130_fd_sc_hd__inv_2 _11267_ (.A(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__or2_1 _11268_ (.A(_04672_),
    .B(_04665_),
    .X(_04679_));
 sky130_fd_sc_hd__o211a_1 _11269_ (.A1(_04673_),
    .A2(_04678_),
    .B1(_04663_),
    .C1(_04679_),
    .X(_04680_));
 sky130_fd_sc_hd__nand2_1 _11270_ (.A(_04675_),
    .B(_04680_),
    .Y(_04682_));
 sky130_fd_sc_hd__nand2_1 _11271_ (.A(_04340_),
    .B(_04357_),
    .Y(_04683_));
 sky130_fd_sc_hd__nand2_1 _11272_ (.A(_04683_),
    .B(_04355_),
    .Y(_04684_));
 sky130_fd_sc_hd__or2_1 _11273_ (.A(_04349_),
    .B(_04684_),
    .X(_04685_));
 sky130_fd_sc_hd__nand2_1 _11274_ (.A(_04684_),
    .B(_04349_),
    .Y(_04686_));
 sky130_fd_sc_hd__a21o_1 _11275_ (.A1(_04685_),
    .A2(_04686_),
    .B1(_04541_),
    .X(_04687_));
 sky130_fd_sc_hd__or2_1 _11276_ (.A(_04345_),
    .B(net101),
    .X(_04688_));
 sky130_fd_sc_hd__nand2_1 _11277_ (.A(_04687_),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__or2_1 _11278_ (.A(\sq.out[18] ),
    .B(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__nand2_1 _11279_ (.A(_04689_),
    .B(\sq.out[18] ),
    .Y(_04691_));
 sky130_fd_sc_hd__nand2_2 _11280_ (.A(_04690_),
    .B(_04691_),
    .Y(_04693_));
 sky130_fd_sc_hd__inv_2 _11281_ (.A(_04693_),
    .Y(_04694_));
 sky130_fd_sc_hd__or2_1 _11282_ (.A(_04357_),
    .B(_04340_),
    .X(_04695_));
 sky130_fd_sc_hd__nand3_1 _11283_ (.A(_04609_),
    .B(_04683_),
    .C(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__nand2_1 _11284_ (.A(_04601_),
    .B(_04353_),
    .Y(_04697_));
 sky130_fd_sc_hd__nand2_1 _11285_ (.A(_04696_),
    .B(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__or2_1 _11286_ (.A(_02877_),
    .B(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__nand2_1 _11287_ (.A(_04698_),
    .B(_02877_),
    .Y(_04700_));
 sky130_fd_sc_hd__nand2_1 _11288_ (.A(_04699_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__inv_2 _11289_ (.A(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand3_1 _11290_ (.A(_04682_),
    .B(_04694_),
    .C(_04702_),
    .Y(_04704_));
 sky130_fd_sc_hd__inv_2 _11291_ (.A(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__clkinvlp_2 _11292_ (.A(_04425_),
    .Y(_04706_));
 sky130_fd_sc_hd__nor2_1 _11293_ (.A(_04450_),
    .B(_04359_),
    .Y(_04707_));
 sky130_fd_sc_hd__o21bai_1 _11294_ (.A1(_04706_),
    .A2(_04707_),
    .B1_N(_04453_),
    .Y(_04708_));
 sky130_fd_sc_hd__or2b_1 _11295_ (.A(_04708_),
    .B_N(_04435_),
    .X(_04709_));
 sky130_fd_sc_hd__nand3_1 _11296_ (.A(_04708_),
    .B(_04433_),
    .C(_04434_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand3_1 _11297_ (.A(_04709_),
    .B(\sq.out[1] ),
    .C(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_1 _11298_ (.A(_04601_),
    .B(_04432_),
    .Y(_04712_));
 sky130_fd_sc_hd__nand2_1 _11299_ (.A(_04711_),
    .B(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__inv_2 _11300_ (.A(_04713_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand2_1 _11301_ (.A(_04715_),
    .B(\sq.out[23] ),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_1 _11302_ (.A(_04713_),
    .B(_01993_),
    .Y(_04717_));
 sky130_fd_sc_hd__nand2_1 _11303_ (.A(_04716_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__nand2_1 _11304_ (.A(_04710_),
    .B(_04433_),
    .Y(_04719_));
 sky130_fd_sc_hd__xor2_1 _11305_ (.A(_04444_),
    .B(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__nand2_1 _11306_ (.A(_04720_),
    .B(\sq.out[1] ),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _11307_ (.A(_04601_),
    .B(_04441_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _11308_ (.A(_04721_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__or2_1 _11309_ (.A(\sq.out[24] ),
    .B(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__nand2_1 _11310_ (.A(_04723_),
    .B(\sq.out[24] ),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_1 _11311_ (.A(_04724_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__nor2_1 _11312_ (.A(_04718_),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__or2_1 _11313_ (.A(_04414_),
    .B(_04609_),
    .X(_04729_));
 sky130_fd_sc_hd__o21ai_1 _11314_ (.A1(_04424_),
    .A2(_04707_),
    .B1(_04422_),
    .Y(_04730_));
 sky130_fd_sc_hd__xor2_1 _11315_ (.A(_04417_),
    .B(_04730_),
    .X(_04731_));
 sky130_fd_sc_hd__nand2_1 _11316_ (.A(_04731_),
    .B(_04609_),
    .Y(_04732_));
 sky130_fd_sc_hd__nand2_1 _11317_ (.A(_04729_),
    .B(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__inv_2 _11318_ (.A(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__nand2_1 _11319_ (.A(_04734_),
    .B(_02009_),
    .Y(_04735_));
 sky130_fd_sc_hd__nand2_1 _11320_ (.A(_04733_),
    .B(\sq.out[22] ),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_2 _11321_ (.A(_04735_),
    .B(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__or2_1 _11322_ (.A(_04421_),
    .B(_04609_),
    .X(_04739_));
 sky130_fd_sc_hd__or2_1 _11323_ (.A(_04424_),
    .B(_04707_),
    .X(_04740_));
 sky130_fd_sc_hd__nand2_1 _11324_ (.A(_04707_),
    .B(_04424_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand3_1 _11325_ (.A(\sq.out[1] ),
    .B(_04740_),
    .C(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_1 _11326_ (.A(_04739_),
    .B(_04742_),
    .Y(_04743_));
 sky130_fd_sc_hd__or2_1 _11327_ (.A(_02927_),
    .B(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__nand2_1 _11328_ (.A(_04743_),
    .B(_02927_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_1 _11329_ (.A(_04744_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__nor2_1 _11330_ (.A(_04738_),
    .B(_04746_),
    .Y(_04748_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(_04728_),
    .B(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__or2_1 _11332_ (.A(_04206_),
    .B(net101),
    .X(_04750_));
 sky130_fd_sc_hd__or2b_1 _11333_ (.A(_04448_),
    .B_N(_04358_),
    .X(_04751_));
 sky130_fd_sc_hd__a21bo_1 _11334_ (.A1(_04751_),
    .A2(_04222_),
    .B1_N(_04221_),
    .X(_04752_));
 sky130_fd_sc_hd__xor2_1 _11335_ (.A(_04209_),
    .B(_04752_),
    .X(_04753_));
 sky130_fd_sc_hd__nand2_1 _11336_ (.A(_04753_),
    .B(_04609_),
    .Y(_04754_));
 sky130_fd_sc_hd__nand2_1 _11337_ (.A(_04750_),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__inv_2 _11338_ (.A(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand2_1 _11339_ (.A(_04756_),
    .B(_01730_),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _11340_ (.A(_04755_),
    .B(\sq.out[20] ),
    .Y(_04759_));
 sky130_fd_sc_hd__nand2_1 _11341_ (.A(_04757_),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__xor2_1 _11342_ (.A(_04223_),
    .B(_04751_),
    .X(_04761_));
 sky130_fd_sc_hd__or2_1 _11343_ (.A(_04761_),
    .B(_04601_),
    .X(_04762_));
 sky130_fd_sc_hd__or2_1 _11344_ (.A(_04219_),
    .B(net101),
    .X(_04763_));
 sky130_fd_sc_hd__nand2_1 _11345_ (.A(_04762_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__or2_1 _11346_ (.A(_05140_),
    .B(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__nand2_1 _11347_ (.A(_04764_),
    .B(_05140_),
    .Y(_04766_));
 sky130_fd_sc_hd__nand2_1 _11348_ (.A(_04765_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hd__nor2_1 _11349_ (.A(_04760_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand3_1 _11350_ (.A(_04705_),
    .B(_04749_),
    .C(_04768_),
    .Y(_04770_));
 sky130_fd_sc_hd__a21oi_2 _11351_ (.A1(_04359_),
    .A2(_04446_),
    .B1(_04456_),
    .Y(_04771_));
 sky130_fd_sc_hd__o211a_1 _11352_ (.A1(_04380_),
    .A2(_04771_),
    .B1(_04457_),
    .C1(\sq.out[1] ),
    .X(_04772_));
 sky130_fd_sc_hd__nand2_1 _11353_ (.A(_04772_),
    .B(_04393_),
    .Y(_04773_));
 sky130_fd_sc_hd__xor2_1 _11354_ (.A(_04398_),
    .B(_04773_),
    .X(_04774_));
 sky130_fd_sc_hd__o21ai_1 _11355_ (.A1(_04379_),
    .A2(_04771_),
    .B1(_04377_),
    .Y(_04775_));
 sky130_fd_sc_hd__or2b_1 _11356_ (.A(_04365_),
    .B_N(_04775_),
    .X(_04776_));
 sky130_fd_sc_hd__and2_1 _11357_ (.A(_04776_),
    .B(_04609_),
    .X(_04777_));
 sky130_fd_sc_hd__nand2b_1 _11358_ (.A_N(_04408_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__xnor2_1 _11359_ (.A(_04402_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__or2_1 _11360_ (.A(_04601_),
    .B(_04776_),
    .X(_04781_));
 sky130_fd_sc_hd__a21bo_1 _11361_ (.A1(_04609_),
    .A2(_04775_),
    .B1_N(_04365_),
    .X(_04782_));
 sky130_fd_sc_hd__nand2_1 _11362_ (.A(_04781_),
    .B(_04782_),
    .Y(_04783_));
 sky130_fd_sc_hd__inv_2 _11363_ (.A(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__nand2b_1 _11364_ (.A_N(_04777_),
    .B(_04408_),
    .Y(_04785_));
 sky130_fd_sc_hd__nand2_1 _11365_ (.A(_04785_),
    .B(_04778_),
    .Y(_04786_));
 sky130_fd_sc_hd__or2_1 _11366_ (.A(_04784_),
    .B(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__xor2_1 _11367_ (.A(_04392_),
    .B(_04772_),
    .X(_04788_));
 sky130_fd_sc_hd__nand2b_1 _11368_ (.A_N(_04387_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__or4_4 _11369_ (.A(_04774_),
    .B(_04779_),
    .C(_04787_),
    .D(_04789_),
    .X(_04790_));
 sky130_fd_sc_hd__o21a_1 _11370_ (.A1(_04700_),
    .A2(_04693_),
    .B1(_04690_),
    .X(_04792_));
 sky130_fd_sc_hd__or3_1 _11371_ (.A(_04760_),
    .B(_04767_),
    .C(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__o211a_1 _11372_ (.A1(_04760_),
    .A2(_04766_),
    .B1(_04757_),
    .C1(_04793_),
    .X(_04794_));
 sky130_fd_sc_hd__nand2b_1 _11373_ (.A_N(_04794_),
    .B(_04749_),
    .Y(_04795_));
 sky130_fd_sc_hd__o21ai_1 _11374_ (.A1(_04745_),
    .A2(_04738_),
    .B1(_04735_),
    .Y(_04796_));
 sky130_fd_sc_hd__inv_2 _11375_ (.A(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__nand3b_1 _11376_ (.A_N(_04717_),
    .B(_04724_),
    .C(_04726_),
    .Y(_04798_));
 sky130_fd_sc_hd__o311a_1 _11377_ (.A1(_04718_),
    .A2(_04797_),
    .A3(_04727_),
    .B1(_04724_),
    .C1(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__nand2_1 _11378_ (.A(_04795_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__nor2_1 _11379_ (.A(_04790_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__nand2_1 _11380_ (.A(_04770_),
    .B(_04801_),
    .Y(_04803_));
 sky130_fd_sc_hd__or2_1 _11381_ (.A(_04379_),
    .B(_04771_),
    .X(_04804_));
 sky130_fd_sc_hd__nand2_1 _11382_ (.A(_04771_),
    .B(_04379_),
    .Y(_04805_));
 sky130_fd_sc_hd__nor2_1 _11383_ (.A(_04375_),
    .B(\sq.out[1] ),
    .Y(_04806_));
 sky130_fd_sc_hd__a31o_1 _11384_ (.A1(\sq.out[1] ),
    .A2(_04804_),
    .A3(_04805_),
    .B1(_04806_),
    .X(_04807_));
 sky130_fd_sc_hd__or2_1 _11385_ (.A(_04807_),
    .B(_04790_),
    .X(_04808_));
 sky130_fd_sc_hd__nand3_4 _11386_ (.A(_04531_),
    .B(_04447_),
    .C(_04459_),
    .Y(_04809_));
 sky130_fd_sc_hd__nor2_4 _11387_ (.A(_04809_),
    .B(_04493_),
    .Y(_04810_));
 sky130_fd_sc_hd__nand2_2 _11388_ (.A(_04810_),
    .B(_04520_),
    .Y(_04811_));
 sky130_fd_sc_hd__xor2_2 _11389_ (.A(_04507_),
    .B(_04811_),
    .X(_04812_));
 sky130_fd_sc_hd__a31o_1 _11390_ (.A1(_04810_),
    .A2(_04520_),
    .A3(_04507_),
    .B1(_04510_),
    .X(_04814_));
 sky130_fd_sc_hd__or2_1 _11391_ (.A(_04511_),
    .B(_04811_),
    .X(_04815_));
 sky130_fd_sc_hd__nand2_1 _11392_ (.A(_04814_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__or2_1 _11393_ (.A(_04812_),
    .B(_04816_),
    .X(_04817_));
 sky130_fd_sc_hd__nand2_1 _11394_ (.A(_04497_),
    .B(_04498_),
    .Y(_04818_));
 sky130_fd_sc_hd__or2_1 _11395_ (.A(_04818_),
    .B(_04815_),
    .X(_04819_));
 sky130_fd_sc_hd__nand2_1 _11396_ (.A(_04815_),
    .B(_04818_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _11397_ (.A(_04819_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__xor2_1 _11398_ (.A(_04190_),
    .B(_04497_),
    .X(_04822_));
 sky130_fd_sc_hd__xnor2_1 _11399_ (.A(_04822_),
    .B(_04819_),
    .Y(_04823_));
 sky130_fd_sc_hd__or2b_1 _11400_ (.A(_04504_),
    .B_N(_04503_),
    .X(_04825_));
 sky130_fd_sc_hd__nand2_1 _11401_ (.A(_04505_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__a31o_1 _11402_ (.A1(_04463_),
    .A2(_04192_),
    .A3(_04175_),
    .B1(_04197_),
    .X(_04827_));
 sky130_fd_sc_hd__nand2_1 _11403_ (.A(_04827_),
    .B(_04503_),
    .Y(_04828_));
 sky130_fd_sc_hd__nand2_1 _11404_ (.A(_04810_),
    .B(_04513_),
    .Y(_04829_));
 sky130_fd_sc_hd__and2_1 _11405_ (.A(_04515_),
    .B(_04516_),
    .X(_04830_));
 sky130_fd_sc_hd__nand2b_1 _11406_ (.A_N(_04829_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__or2_1 _11407_ (.A(_04828_),
    .B(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__xor2_1 _11408_ (.A(_04826_),
    .B(_04832_),
    .X(_04833_));
 sky130_fd_sc_hd__nand2_1 _11409_ (.A(_04831_),
    .B(_04828_),
    .Y(_04834_));
 sky130_fd_sc_hd__nand2_1 _11410_ (.A(_04832_),
    .B(_04834_),
    .Y(_04836_));
 sky130_fd_sc_hd__or2_1 _11411_ (.A(_04513_),
    .B(_04810_),
    .X(_04837_));
 sky130_fd_sc_hd__nand2_1 _11412_ (.A(_04837_),
    .B(_04829_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21o_1 _11413_ (.A1(_04810_),
    .A2(_04513_),
    .B1(_04830_),
    .X(_04839_));
 sky130_fd_sc_hd__nand2_1 _11414_ (.A(_04831_),
    .B(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hd__or2_1 _11415_ (.A(_04838_),
    .B(_04840_),
    .X(_04841_));
 sky130_fd_sc_hd__nor2_1 _11416_ (.A(_04836_),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__nand2_1 _11417_ (.A(_04833_),
    .B(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__or4_4 _11418_ (.A(_04817_),
    .B(_04821_),
    .C(_04823_),
    .D(_04843_),
    .X(_04844_));
 sky130_fd_sc_hd__nor2_1 _11419_ (.A(_04475_),
    .B(_04809_),
    .Y(_04845_));
 sky130_fd_sc_hd__inv_2 _11420_ (.A(_04845_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_1 _11421_ (.A(_04809_),
    .B(_04475_),
    .Y(_04848_));
 sky130_fd_sc_hd__nand2_1 _11422_ (.A(_04847_),
    .B(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__nor2_1 _11423_ (.A(_04482_),
    .B(_04845_),
    .Y(_04850_));
 sky130_fd_sc_hd__nor2_1 _11424_ (.A(_04481_),
    .B(_04847_),
    .Y(_04851_));
 sky130_fd_sc_hd__or2_1 _11425_ (.A(_04850_),
    .B(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__or2_1 _11426_ (.A(_04849_),
    .B(_04852_),
    .X(_04853_));
 sky130_fd_sc_hd__inv_2 _11427_ (.A(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__nand2_1 _11428_ (.A(_04851_),
    .B(_04479_),
    .Y(_04855_));
 sky130_fd_sc_hd__xnor2_1 _11429_ (.A(_04487_),
    .B(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__inv_2 _11430_ (.A(_04856_),
    .Y(_04858_));
 sky130_fd_sc_hd__or2_1 _11431_ (.A(_04479_),
    .B(_04851_),
    .X(_04859_));
 sky130_fd_sc_hd__nand2_1 _11432_ (.A(_04859_),
    .B(_04855_),
    .Y(_04860_));
 sky130_fd_sc_hd__inv_2 _11433_ (.A(_04860_),
    .Y(_04861_));
 sky130_fd_sc_hd__and3_1 _11434_ (.A(_04854_),
    .B(_04858_),
    .C(_04861_),
    .X(_04862_));
 sky130_fd_sc_hd__inv_2 _11435_ (.A(_04491_),
    .Y(_04863_));
 sky130_fd_sc_hd__nor2b_2 _11436_ (.A(_04809_),
    .B_N(_04488_),
    .Y(_04864_));
 sky130_fd_sc_hd__xor2_2 _11437_ (.A(_04863_),
    .B(_04864_),
    .X(_04865_));
 sky130_fd_sc_hd__clkinvlp_2 _11438_ (.A(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__a21bo_1 _11439_ (.A1(_04864_),
    .A2(_04863_),
    .B1_N(_04490_),
    .X(_04867_));
 sky130_fd_sc_hd__nand2_1 _11440_ (.A(_04864_),
    .B(_04492_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_1 _11441_ (.A(_04867_),
    .B(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__nor2_1 _11442_ (.A(_04866_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__or2_1 _11443_ (.A(_04468_),
    .B(_04869_),
    .X(_04872_));
 sky130_fd_sc_hd__xor2_1 _11444_ (.A(_04471_),
    .B(_04872_),
    .X(_04873_));
 sky130_fd_sc_hd__nand2_1 _11445_ (.A(_04869_),
    .B(_04468_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand2_1 _11446_ (.A(_04872_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__inv_2 _11447_ (.A(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__and4_2 _11448_ (.A(_04862_),
    .B(_04871_),
    .C(_04873_),
    .D(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__nand2b_4 _11449_ (.A_N(_04844_),
    .B(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__a21oi_1 _11450_ (.A1(_04803_),
    .A2(_04808_),
    .B1(_04878_),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _11451_ (.A(\sq.out[1] ),
    .B(_04534_),
    .Y(_04881_));
 sky130_fd_sc_hd__nand2_1 _11452_ (.A(_04523_),
    .B(_04526_),
    .Y(_04882_));
 sky130_fd_sc_hd__nand2_2 _11453_ (.A(_04881_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__clkinvlp_2 _11454_ (.A(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nor2_2 _11455_ (.A(_04529_),
    .B(_04534_),
    .Y(_04885_));
 sky130_fd_sc_hd__inv_2 _11456_ (.A(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand3_2 _11457_ (.A(_04880_),
    .B(_04884_),
    .C(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__buf_6 _11458_ (.A(_04887_),
    .X(_04888_));
 sky130_fd_sc_hd__nand2_1 _11459_ (.A(_04803_),
    .B(_04808_),
    .Y(_04889_));
 sky130_fd_sc_hd__buf_6 _11460_ (.A(_04889_),
    .X(_04891_));
 sky130_fd_sc_hd__nand3_1 _11461_ (.A(_04891_),
    .B(_04862_),
    .C(_04871_),
    .Y(_04892_));
 sky130_fd_sc_hd__inv_2 _11462_ (.A(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand3_1 _11463_ (.A(_04888_),
    .B(_04876_),
    .C(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__and2_1 _11464_ (.A(_04891_),
    .B(_04854_),
    .X(_04895_));
 sky130_fd_sc_hd__nand3_1 _11465_ (.A(_04888_),
    .B(_04861_),
    .C(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__nand2_1 _11466_ (.A(_04894_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__inv_2 _11467_ (.A(_04878_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand3_1 _11468_ (.A(_04891_),
    .B(_04884_),
    .C(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__o21ai_1 _11469_ (.A1(_04885_),
    .A2(_04899_),
    .B1(\sq.out[2] ),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_1 _11470_ (.A(_04900_),
    .B(\sq.out[1] ),
    .Y(_04902_));
 sky130_fd_sc_hd__o31ai_1 _11471_ (.A1(_04883_),
    .A2(_04878_),
    .A3(_04885_),
    .B1(_04889_),
    .Y(_04903_));
 sky130_fd_sc_hd__nand2_1 _11472_ (.A(_04903_),
    .B(_04849_),
    .Y(_04904_));
 sky130_fd_sc_hd__nand2_1 _11473_ (.A(_04902_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__nor2_1 _11474_ (.A(_04897_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__and2_1 _11475_ (.A(_04891_),
    .B(_04862_),
    .X(_04907_));
 sky130_fd_sc_hd__nand3_1 _11476_ (.A(_04887_),
    .B(_04865_),
    .C(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__or2_1 _11477_ (.A(_04849_),
    .B(_04903_),
    .X(_04909_));
 sky130_fd_sc_hd__o311ai_2 _11478_ (.A1(_04883_),
    .A2(_04885_),
    .A3(_04878_),
    .B1(_04862_),
    .C1(_04891_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand2_1 _11479_ (.A(_04910_),
    .B(_04866_),
    .Y(_04911_));
 sky130_fd_sc_hd__nand3_1 _11480_ (.A(_04908_),
    .B(_04909_),
    .C(_04911_),
    .Y(_04913_));
 sky130_fd_sc_hd__inv_2 _11481_ (.A(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand2_1 _11482_ (.A(_04906_),
    .B(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__inv_2 _11483_ (.A(_04843_),
    .Y(_04916_));
 sky130_fd_sc_hd__nand3_2 _11484_ (.A(_04891_),
    .B(_04877_),
    .C(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__inv_2 _11485_ (.A(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__o21ai_1 _11486_ (.A1(_04885_),
    .A2(_04899_),
    .B1(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__nand2_1 _11487_ (.A(_04919_),
    .B(_04812_),
    .Y(_04920_));
 sky130_fd_sc_hd__inv_2 _11488_ (.A(_04812_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand3_1 _11489_ (.A(_04888_),
    .B(_04921_),
    .C(_04918_),
    .Y(_04922_));
 sky130_fd_sc_hd__nand2_1 _11490_ (.A(_04920_),
    .B(_04922_),
    .Y(_04924_));
 sky130_fd_sc_hd__nand3b_1 _11491_ (.A_N(_04841_),
    .B(_04891_),
    .C(_04877_),
    .Y(_04925_));
 sky130_fd_sc_hd__inv_2 _11492_ (.A(_04925_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand2_1 _11493_ (.A(_04888_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand2_1 _11494_ (.A(_04927_),
    .B(_04836_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _11495_ (.A(_04887_),
    .B(_04895_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _11496_ (.A(_04929_),
    .B(_04860_),
    .Y(_04930_));
 sky130_fd_sc_hd__nand2_1 _11497_ (.A(_04928_),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__nor2_1 _11498_ (.A(_04924_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__inv_2 _11499_ (.A(_04838_),
    .Y(_04933_));
 sky130_fd_sc_hd__and2_1 _11500_ (.A(_04891_),
    .B(_04877_),
    .X(_04935_));
 sky130_fd_sc_hd__nand3_1 _11501_ (.A(_04888_),
    .B(_04933_),
    .C(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__o311ai_1 _11502_ (.A1(_04883_),
    .A2(_04844_),
    .A3(_04885_),
    .B1(_04877_),
    .C1(_04891_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand2_1 _11503_ (.A(_04937_),
    .B(_04838_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_1 _11504_ (.A(_04936_),
    .B(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _11505_ (.A(_04888_),
    .B(_04893_),
    .Y(_04940_));
 sky130_fd_sc_hd__nand2_1 _11506_ (.A(_04940_),
    .B(_04875_),
    .Y(_04941_));
 sky130_fd_sc_hd__nor2_1 _11507_ (.A(_04817_),
    .B(_04917_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand3b_1 _11508_ (.A_N(_04821_),
    .B(_04888_),
    .C(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__nand2_1 _11509_ (.A(_04941_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__nor2_1 _11510_ (.A(_04939_),
    .B(_04944_),
    .Y(_04946_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(_04932_),
    .B(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__nor2_4 _11512_ (.A(_04915_),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_1 _11513_ (.A(_04891_),
    .B(_04898_),
    .Y(_04949_));
 sky130_fd_sc_hd__or3_1 _11514_ (.A(_04883_),
    .B(_04886_),
    .C(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__nand2_1 _11515_ (.A(_04888_),
    .B(_04942_),
    .Y(_04951_));
 sky130_fd_sc_hd__nand2_1 _11516_ (.A(_04951_),
    .B(_04821_),
    .Y(_04952_));
 sky130_fd_sc_hd__nand2_1 _11517_ (.A(_04950_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__inv_2 _11518_ (.A(_04800_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _11519_ (.A(_04770_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _11520_ (.A(_04955_),
    .B(_04807_),
    .Y(_04957_));
 sky130_fd_sc_hd__nand2_1 _11521_ (.A(_04957_),
    .B(_04783_),
    .Y(_04958_));
 sky130_fd_sc_hd__nand2_1 _11522_ (.A(_04958_),
    .B(_04786_),
    .Y(_04959_));
 sky130_fd_sc_hd__or4_1 _11523_ (.A(_04840_),
    .B(_04774_),
    .C(_04870_),
    .D(_04789_),
    .X(_04960_));
 sky130_fd_sc_hd__or3b_1 _11524_ (.A(_04823_),
    .B(_04960_),
    .C_N(_04833_),
    .X(_04961_));
 sky130_fd_sc_hd__a2111oi_1 _11525_ (.A1(_04784_),
    .A2(_04807_),
    .B1(_04852_),
    .C1(_04779_),
    .D1(_04816_),
    .Y(_04962_));
 sky130_fd_sc_hd__and4b_1 _11526_ (.A_N(_04961_),
    .B(_04858_),
    .C(_04873_),
    .D(_04962_),
    .X(_04963_));
 sky130_fd_sc_hd__nand2_1 _11527_ (.A(_04959_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__a21oi_1 _11528_ (.A1(_04885_),
    .A2(_04899_),
    .B1(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_1 _11529_ (.A(_04949_),
    .B(_04883_),
    .Y(_04966_));
 sky130_fd_sc_hd__inv_2 _11530_ (.A(_04887_),
    .Y(_04968_));
 sky130_fd_sc_hd__or4_1 _11531_ (.A(_04549_),
    .B(_04569_),
    .C(_04615_),
    .D(_04580_),
    .X(_04969_));
 sky130_fd_sc_hd__or4_1 _11532_ (.A(_04669_),
    .B(_04623_),
    .C(_04642_),
    .D(_04648_),
    .X(_04970_));
 sky130_fd_sc_hd__inv_2 _11533_ (.A(_04535_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand2_1 _11534_ (.A(_04662_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__or4_1 _11535_ (.A(_04603_),
    .B(_04589_),
    .C(_04560_),
    .D(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__or3_1 _11536_ (.A(_04969_),
    .B(_04970_),
    .C(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__nand2_1 _11537_ (.A(_04968_),
    .B(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__nand3_2 _11538_ (.A(_04965_),
    .B(_04966_),
    .C(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__o21ai_1 _11539_ (.A1(_04783_),
    .A2(_04955_),
    .B1(_04957_),
    .Y(_04977_));
 sky130_fd_sc_hd__inv_2 _11540_ (.A(_04977_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand2_1 _11541_ (.A(_04682_),
    .B(_04702_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2_1 _11542_ (.A(_04980_),
    .B(_04700_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2b_1 _11543_ (.A_N(_04981_),
    .B(_04694_),
    .Y(_04982_));
 sky130_fd_sc_hd__nand3_1 _11544_ (.A(_04675_),
    .B(_04701_),
    .C(_04680_),
    .Y(_04983_));
 sky130_fd_sc_hd__nand2_1 _11545_ (.A(_04617_),
    .B(\sq.out[11] ),
    .Y(_04984_));
 sky130_fd_sc_hd__nand2_1 _11546_ (.A(_04984_),
    .B(_04628_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_1 _11547_ (.A(_04604_),
    .B(_04607_),
    .Y(_04986_));
 sky130_fd_sc_hd__or2_1 _11548_ (.A(_04986_),
    .B(_04598_),
    .X(_04987_));
 sky130_fd_sc_hd__and2_1 _11549_ (.A(_04738_),
    .B(_04744_),
    .X(_04988_));
 sky130_fd_sc_hd__a211oi_1 _11550_ (.A1(_04626_),
    .A2(_04984_),
    .B1(_04988_),
    .C1(_04595_),
    .Y(_04990_));
 sky130_fd_sc_hd__nand2_1 _11551_ (.A(_04673_),
    .B(_04677_),
    .Y(_04991_));
 sky130_fd_sc_hd__o211ai_1 _11552_ (.A1(\sq.out[3] ),
    .A2(_04971_),
    .B1(_04564_),
    .C1(_04581_),
    .Y(_04992_));
 sky130_fd_sc_hd__nand3_1 _11553_ (.A(_04574_),
    .B(_04562_),
    .C(_04554_),
    .Y(_04993_));
 sky130_fd_sc_hd__nor3_1 _11554_ (.A(_04543_),
    .B(_04992_),
    .C(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nand3_1 _11555_ (.A(_04990_),
    .B(_04991_),
    .C(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__nand3_1 _11556_ (.A(_04727_),
    .B(\sq.out[23] ),
    .C(_04715_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _11557_ (.A(_04996_),
    .B(_04798_),
    .Y(_04997_));
 sky130_fd_sc_hd__nand2_1 _11558_ (.A(_04997_),
    .B(_04797_),
    .Y(_04998_));
 sky130_fd_sc_hd__o21ai_1 _11559_ (.A1(_04748_),
    .A2(_04796_),
    .B1(_04728_),
    .Y(_04999_));
 sky130_fd_sc_hd__nand2_1 _11560_ (.A(_04998_),
    .B(_04999_),
    .Y(_05001_));
 sky130_fd_sc_hd__inv_2 _11561_ (.A(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hd__nor2_1 _11562_ (.A(_04995_),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__nand2_1 _11563_ (.A(_04598_),
    .B(_04986_),
    .Y(_05004_));
 sky130_fd_sc_hd__nand3_1 _11564_ (.A(_04987_),
    .B(_05003_),
    .C(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__a21oi_1 _11565_ (.A1(_04608_),
    .A2(_04985_),
    .B1(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__a31o_1 _11566_ (.A1(_04606_),
    .A2(_04607_),
    .A3(_04632_),
    .B1(_04674_),
    .X(_05007_));
 sky130_fd_sc_hd__a21o_1 _11567_ (.A1(_04663_),
    .A2(_04664_),
    .B1(_04671_),
    .X(_05008_));
 sky130_fd_sc_hd__nand3_1 _11568_ (.A(_04678_),
    .B(_04679_),
    .C(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__inv_2 _11569_ (.A(_04645_),
    .Y(_05010_));
 sky130_fd_sc_hd__o21ai_1 _11570_ (.A1(_05010_),
    .A2(_04650_),
    .B1(_04676_),
    .Y(_05012_));
 sky130_fd_sc_hd__a21bo_1 _11571_ (.A1(_05009_),
    .A2(_05012_),
    .B1_N(_04632_),
    .X(_05013_));
 sky130_fd_sc_hd__a21o_1 _11572_ (.A1(_05013_),
    .A2(_04629_),
    .B1(_04608_),
    .X(_05014_));
 sky130_fd_sc_hd__nand3_1 _11573_ (.A(_05006_),
    .B(_05007_),
    .C(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__a21oi_1 _11574_ (.A1(_04980_),
    .A2(_04983_),
    .B1(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__nand2_1 _11575_ (.A(_04981_),
    .B(_04693_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand3_1 _11576_ (.A(_04982_),
    .B(_05016_),
    .C(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__clkinvlp_2 _11577_ (.A(_04760_),
    .Y(_05019_));
 sky130_fd_sc_hd__o21a_1 _11578_ (.A1(_04765_),
    .A2(_05019_),
    .B1(_04766_),
    .X(_05020_));
 sky130_fd_sc_hd__nand2_1 _11579_ (.A(_04704_),
    .B(_04792_),
    .Y(_05021_));
 sky130_fd_sc_hd__inv_2 _11580_ (.A(_04767_),
    .Y(_05023_));
 sky130_fd_sc_hd__nand2_1 _11581_ (.A(_05021_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__o21ai_1 _11582_ (.A1(_05020_),
    .A2(_05021_),
    .B1(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hd__inv_2 _11583_ (.A(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nor2_1 _11584_ (.A(_05018_),
    .B(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__clkinvlp_2 _11585_ (.A(_04738_),
    .Y(_05028_));
 sky130_fd_sc_hd__o21a_1 _11586_ (.A1(_04744_),
    .A2(_05028_),
    .B1(_04745_),
    .X(_05029_));
 sky130_fd_sc_hd__nand2_1 _11587_ (.A(_04705_),
    .B(_04768_),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(_05030_),
    .B(_04794_),
    .Y(_05031_));
 sky130_fd_sc_hd__a21oi_1 _11589_ (.A1(_05028_),
    .A2(_04718_),
    .B1(_04746_),
    .Y(_05032_));
 sky130_fd_sc_hd__nand2_1 _11590_ (.A(_05031_),
    .B(_05032_),
    .Y(_05034_));
 sky130_fd_sc_hd__o21ai_1 _11591_ (.A1(_05029_),
    .A2(_05031_),
    .B1(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__a21o_1 _11592_ (.A1(_05024_),
    .A2(_04766_),
    .B1(_05019_),
    .X(_05036_));
 sky130_fd_sc_hd__nand3_2 _11593_ (.A(_05027_),
    .B(_05035_),
    .C(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nor2_2 _11594_ (.A(_04979_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _11595_ (.A(_05038_),
    .B(_04888_),
    .Y(_05039_));
 sky130_fd_sc_hd__a2111o_1 _11596_ (.A1(_04687_),
    .A2(_04688_),
    .B1(_04698_),
    .C1(_04756_),
    .D1(_04764_),
    .X(_05040_));
 sky130_fd_sc_hd__or4_1 _11597_ (.A(_04713_),
    .B(_04743_),
    .C(_04734_),
    .D(_04807_),
    .X(_05041_));
 sky130_fd_sc_hd__a2111o_1 _11598_ (.A1(_04721_),
    .A2(_04722_),
    .B1(_04786_),
    .C1(_05040_),
    .D1(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__a21oi_1 _11599_ (.A1(_04957_),
    .A2(_04784_),
    .B1(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_1 _11600_ (.A(_04968_),
    .B(_05043_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_1 _11601_ (.A(_05039_),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__nand3b_1 _11602_ (.A_N(_04836_),
    .B(_04888_),
    .C(_04926_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_1 _11603_ (.A(_05046_),
    .B(_05047_),
    .Y(_05048_));
 sky130_fd_sc_hd__nor3_4 _11604_ (.A(_04953_),
    .B(_04976_),
    .C(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__inv_2 _11605_ (.A(net146),
    .Y(_05050_));
 sky130_fd_sc_hd__nand3_4 _11606_ (.A(_04948_),
    .B(_05049_),
    .C(net147),
    .Y(_05051_));
 sky130_fd_sc_hd__buf_6 _11607_ (.A(_05051_),
    .X(_05052_));
 sky130_fd_sc_hd__inv_2 _11608_ (.A(net33),
    .Y(_05053_));
 sky130_fd_sc_hd__and2_1 _11609_ (.A(_05053_),
    .B(net34),
    .X(_05054_));
 sky130_fd_sc_hd__inv_2 _11610_ (.A(_05054_),
    .Y(_05056_));
 sky130_fd_sc_hd__nor2_4 _11611_ (.A(net35),
    .B(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hd__buf_6 _11612_ (.A(_05057_),
    .X(_05058_));
 sky130_fd_sc_hd__inv_2 _11613_ (.A(net35),
    .Y(_05059_));
 sky130_fd_sc_hd__or4_1 _11614_ (.A(net34),
    .B(net33),
    .C(_05050_),
    .D(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__clkbuf_4 _11615_ (.A(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__inv_2 _11616_ (.A(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__buf_6 _11617_ (.A(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__a21o_1 _11618_ (.A1(_05052_),
    .A2(_05058_),
    .B1(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__or2_1 _11619_ (.A(_01298_),
    .B(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__nand2_1 _11620_ (.A(_05064_),
    .B(_01298_),
    .Y(_05067_));
 sky130_fd_sc_hd__nor2_1 _11621_ (.A(net34),
    .B(_05053_),
    .Y(_05068_));
 sky130_fd_sc_hd__inv_2 _11622_ (.A(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__nor2_4 _11623_ (.A(net35),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hd__inv_2 _11624_ (.A(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__buf_6 _11625_ (.A(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__nand3_1 _11626_ (.A(_05065_),
    .B(_05067_),
    .C(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_4 _11627_ (.A(_04948_),
    .B(_05049_),
    .Y(_05074_));
 sky130_fd_sc_hd__buf_6 _11628_ (.A(net146),
    .X(_05075_));
 sky130_fd_sc_hd__nand2_2 _11629_ (.A(_05074_),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__buf_6 _11630_ (.A(_05075_),
    .X(_05078_));
 sky130_fd_sc_hd__mux2_1 _11631_ (.A0(_05076_),
    .A1(_05078_),
    .S(net142),
    .X(_05079_));
 sky130_fd_sc_hd__buf_6 _11632_ (.A(_05070_),
    .X(_05080_));
 sky130_fd_sc_hd__buf_6 _11633_ (.A(_05080_),
    .X(_05081_));
 sky130_fd_sc_hd__nand2_1 _11634_ (.A(_05079_),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__nand2_1 _11635_ (.A(_05073_),
    .B(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__and3_1 _11636_ (.A(_05056_),
    .B(_05069_),
    .C(_05059_),
    .X(_05084_));
 sky130_fd_sc_hd__buf_6 _11637_ (.A(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__inv_2 _11638_ (.A(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__buf_6 _11639_ (.A(_05086_),
    .X(_05087_));
 sky130_fd_sc_hd__buf_6 _11640_ (.A(_05087_),
    .X(_05089_));
 sky130_fd_sc_hd__buf_6 _11641_ (.A(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__nor2_1 _11642_ (.A(net142),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__a211o_1 _11643_ (.A1(_05083_),
    .A2(_05090_),
    .B1(net133),
    .C1(net143),
    .X(_05092_));
 sky130_fd_sc_hd__inv_2 _11644_ (.A(_05092_),
    .Y(_00002_));
 sky130_fd_sc_hd__inv_2 _11645_ (.A(net158),
    .Y(_05093_));
 sky130_fd_sc_hd__buf_6 _11646_ (.A(_05085_),
    .X(_05094_));
 sky130_fd_sc_hd__buf_6 _11647_ (.A(_05057_),
    .X(_05095_));
 sky130_fd_sc_hd__nor2_1 _11648_ (.A(net142),
    .B(net158),
    .Y(_05096_));
 sky130_fd_sc_hd__nand2_1 _11649_ (.A(net142),
    .B(net158),
    .Y(_05097_));
 sky130_fd_sc_hd__clkinvlp_2 _11650_ (.A(_05097_),
    .Y(_05099_));
 sky130_fd_sc_hd__nor2_1 _11651_ (.A(_05096_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _11652_ (.A(_05052_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__o211ai_1 _11653_ (.A1(net159),
    .A2(_05052_),
    .B1(_05095_),
    .C1(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__nor2_1 _11654_ (.A(net159),
    .B(_05062_),
    .Y(_05103_));
 sky130_fd_sc_hd__a211o_1 _11655_ (.A1(_05062_),
    .A2(_05100_),
    .B1(_05057_),
    .C1(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__nand2_1 _11656_ (.A(_05102_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__buf_6 _11657_ (.A(_05075_),
    .X(_05106_));
 sky130_fd_sc_hd__nor2_1 _11658_ (.A(_05106_),
    .B(net158),
    .Y(_05107_));
 sky130_fd_sc_hd__nor2_1 _11659_ (.A(net147),
    .B(_05100_),
    .Y(_05108_));
 sky130_fd_sc_hd__buf_6 _11660_ (.A(_05070_),
    .X(_05110_));
 sky130_fd_sc_hd__o21a_1 _11661_ (.A1(_05107_),
    .A2(_05108_),
    .B1(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a21oi_2 _11662_ (.A1(_05105_),
    .A2(_05072_),
    .B1(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__nor2_1 _11663_ (.A(_05094_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__a211o_1 _11664_ (.A1(net159),
    .A2(_05094_),
    .B1(net133),
    .C1(_05113_),
    .X(_05114_));
 sky130_fd_sc_hd__inv_2 _11665_ (.A(_05114_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_1 _11666_ (.A(_05099_),
    .B(net150),
    .Y(_05115_));
 sky130_fd_sc_hd__inv_1 _11667_ (.A(net150),
    .Y(_05116_));
 sky130_fd_sc_hd__nand2_1 _11668_ (.A(_05097_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _11669_ (.A(_05115_),
    .B(_05117_),
    .Y(_05118_));
 sky130_fd_sc_hd__buf_6 _11670_ (.A(_05061_),
    .X(_05120_));
 sky130_fd_sc_hd__clkbuf_4 _11671_ (.A(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__nor2_1 _11672_ (.A(_05118_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__a21o_1 _11673_ (.A1(_05121_),
    .A2(net150),
    .B1(_05058_),
    .X(_05123_));
 sky130_fd_sc_hd__buf_6 _11674_ (.A(_05051_),
    .X(_05124_));
 sky130_fd_sc_hd__nand3_1 _11675_ (.A(_05052_),
    .B(_05115_),
    .C(_05117_),
    .Y(_05125_));
 sky130_fd_sc_hd__o211ai_1 _11676_ (.A1(_05116_),
    .A2(_05124_),
    .B1(_05095_),
    .C1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__o21ai_1 _11677_ (.A1(_05122_),
    .A2(_05123_),
    .B1(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _11678_ (.A(_05127_),
    .B(_05072_),
    .Y(_05128_));
 sky130_fd_sc_hd__nand2_1 _11679_ (.A(_05118_),
    .B(_05106_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(net147),
    .B(_05116_),
    .Y(_05131_));
 sky130_fd_sc_hd__a21oi_1 _11681_ (.A1(_05129_),
    .A2(_05131_),
    .B1(_05071_),
    .Y(_05132_));
 sky130_fd_sc_hd__inv_2 _11682_ (.A(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand2_1 _11683_ (.A(_05128_),
    .B(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hd__nor2_1 _11684_ (.A(net150),
    .B(_05090_),
    .Y(_05135_));
 sky130_fd_sc_hd__a211o_1 _11685_ (.A1(_05134_),
    .A2(_05090_),
    .B1(net133),
    .C1(net151),
    .X(_05136_));
 sky130_fd_sc_hd__inv_2 _11686_ (.A(_05136_),
    .Y(_00024_));
 sky130_fd_sc_hd__inv_2 _11687_ (.A(net200),
    .Y(_05137_));
 sky130_fd_sc_hd__nor2_1 _11688_ (.A(_05137_),
    .B(_05115_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_1 _11689_ (.A(_05115_),
    .B(_05137_),
    .Y(_05139_));
 sky130_fd_sc_hd__or2b_1 _11690_ (.A(_05138_),
    .B_N(_05139_),
    .X(_05141_));
 sky130_fd_sc_hd__o21bai_1 _11691_ (.A1(_05106_),
    .A2(_05074_),
    .B1_N(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__o211ai_1 _11692_ (.A1(_05137_),
    .A2(_05124_),
    .B1(_05095_),
    .C1(_05142_),
    .Y(_05143_));
 sky130_fd_sc_hd__nor2_1 _11693_ (.A(_05141_),
    .B(_05120_),
    .Y(_05144_));
 sky130_fd_sc_hd__a211o_1 _11694_ (.A1(net139),
    .A2(_05120_),
    .B1(_05057_),
    .C1(_05144_),
    .X(_05145_));
 sky130_fd_sc_hd__nand2_1 _11695_ (.A(_05143_),
    .B(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__nand2_1 _11696_ (.A(_05141_),
    .B(_05078_),
    .Y(_05147_));
 sky130_fd_sc_hd__nand2_1 _11697_ (.A(net147),
    .B(_05137_),
    .Y(_05148_));
 sky130_fd_sc_hd__a21oi_1 _11698_ (.A1(_05147_),
    .A2(net148),
    .B1(_05072_),
    .Y(_05149_));
 sky130_fd_sc_hd__a21oi_2 _11699_ (.A1(_05146_),
    .A2(_05072_),
    .B1(net149),
    .Y(_05150_));
 sky130_fd_sc_hd__nor2_1 _11700_ (.A(_05094_),
    .B(_05150_),
    .Y(_05152_));
 sky130_fd_sc_hd__a211o_1 _11701_ (.A1(_05137_),
    .A2(_05094_),
    .B1(net133),
    .C1(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__inv_2 _11702_ (.A(_05153_),
    .Y(_00026_));
 sky130_fd_sc_hd__or2_1 _11703_ (.A(net154),
    .B(_05138_),
    .X(_05154_));
 sky130_fd_sc_hd__nand2_1 _11704_ (.A(_05138_),
    .B(net154),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_1 _11705_ (.A(_05154_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__clkinvlp_2 _11706_ (.A(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand3_4 _11707_ (.A(_04948_),
    .B(_05049_),
    .C(net146),
    .Y(_05158_));
 sky130_fd_sc_hd__buf_4 _11708_ (.A(_05158_),
    .X(_05159_));
 sky130_fd_sc_hd__nor2_1 _11709_ (.A(_05157_),
    .B(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__buf_6 _11710_ (.A(_05074_),
    .X(_05162_));
 sky130_fd_sc_hd__nand3_1 _11711_ (.A(_05162_),
    .B(_05078_),
    .C(_05156_),
    .Y(_05163_));
 sky130_fd_sc_hd__buf_6 _11712_ (.A(net146),
    .X(_05164_));
 sky130_fd_sc_hd__o21a_1 _11713_ (.A1(_05164_),
    .A2(net154),
    .B1(_05110_),
    .X(_05165_));
 sky130_fd_sc_hd__nand2_1 _11714_ (.A(_05163_),
    .B(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__nor2_1 _11715_ (.A(_05160_),
    .B(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__nor2_1 _11716_ (.A(_05094_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__inv_2 _11717_ (.A(net154),
    .Y(_05169_));
 sky130_fd_sc_hd__buf_6 _11718_ (.A(_05051_),
    .X(_05170_));
 sky130_fd_sc_hd__nor2_1 _11719_ (.A(_05169_),
    .B(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__buf_6 _11720_ (.A(_05051_),
    .X(_05173_));
 sky130_fd_sc_hd__nand2_1 _11721_ (.A(net102),
    .B(_05157_),
    .Y(_05174_));
 sky130_fd_sc_hd__buf_6 _11722_ (.A(_05058_),
    .X(_05175_));
 sky130_fd_sc_hd__nand2_1 _11723_ (.A(_05174_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__buf_6 _11724_ (.A(_05057_),
    .X(_05177_));
 sky130_fd_sc_hd__mux2_1 _11725_ (.A0(_05157_),
    .A1(net154),
    .S(_05120_),
    .X(_05178_));
 sky130_fd_sc_hd__o21a_1 _11726_ (.A1(_05177_),
    .A2(_05178_),
    .B1(_05072_),
    .X(_05179_));
 sky130_fd_sc_hd__o21ai_1 _11727_ (.A1(_05171_),
    .A2(_05176_),
    .B1(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand2_1 _11728_ (.A(_05168_),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__clkbuf_4 _11729_ (.A(_05086_),
    .X(_05182_));
 sky130_fd_sc_hd__nor2_1 _11730_ (.A(net154),
    .B(_05182_),
    .Y(_05184_));
 sky130_fd_sc_hd__inv_2 _11731_ (.A(net155),
    .Y(_05185_));
 sky130_fd_sc_hd__nand2_1 _11732_ (.A(_05181_),
    .B(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__or2_1 _11733_ (.A(_01277_),
    .B(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__inv_2 _11734_ (.A(_05187_),
    .Y(_00027_));
 sky130_fd_sc_hd__inv_2 _11735_ (.A(net152),
    .Y(_05188_));
 sky130_fd_sc_hd__or2_1 _11736_ (.A(_05188_),
    .B(_05155_),
    .X(_05189_));
 sky130_fd_sc_hd__nand2_1 _11737_ (.A(_05155_),
    .B(_05188_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand2_1 _11738_ (.A(_05189_),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__clkinvlp_2 _11739_ (.A(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__nor2_1 _11740_ (.A(_05192_),
    .B(_05158_),
    .Y(_05194_));
 sky130_fd_sc_hd__nand3_1 _11741_ (.A(_05074_),
    .B(_05106_),
    .C(_05191_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21a_1 _11742_ (.A1(_05075_),
    .A2(net152),
    .B1(_05080_),
    .X(_05196_));
 sky130_fd_sc_hd__nand2_1 _11743_ (.A(_05195_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__nor2_1 _11744_ (.A(_05194_),
    .B(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__nor2_1 _11745_ (.A(_05085_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__inv_2 _11746_ (.A(_05051_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand2_1 _11747_ (.A(_05200_),
    .B(net152),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_1 _11748_ (.A(_05052_),
    .B(_05192_),
    .Y(_05202_));
 sky130_fd_sc_hd__nand3_1 _11749_ (.A(_05201_),
    .B(_05095_),
    .C(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(_05192_),
    .A1(net152),
    .S(_05061_),
    .X(_05205_));
 sky130_fd_sc_hd__o21a_1 _11751_ (.A1(_05058_),
    .A2(_05205_),
    .B1(_05071_),
    .X(_05206_));
 sky130_fd_sc_hd__nand2_1 _11752_ (.A(_05203_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__nand2_1 _11753_ (.A(_05199_),
    .B(_05207_),
    .Y(_05208_));
 sky130_fd_sc_hd__nor2_1 _11754_ (.A(net152),
    .B(_05182_),
    .Y(_05209_));
 sky130_fd_sc_hd__inv_2 _11755_ (.A(net153),
    .Y(_05210_));
 sky130_fd_sc_hd__nand2_1 _11756_ (.A(_05208_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__or2_1 _11757_ (.A(_01277_),
    .B(_05211_),
    .X(_05212_));
 sky130_fd_sc_hd__inv_2 _11758_ (.A(_05212_),
    .Y(_00028_));
 sky130_fd_sc_hd__clkinvlp_2 _11759_ (.A(net144),
    .Y(_05213_));
 sky130_fd_sc_hd__or2_1 _11760_ (.A(_05213_),
    .B(_05189_),
    .X(_05215_));
 sky130_fd_sc_hd__nand2_1 _11761_ (.A(_05189_),
    .B(_05213_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_1 _11762_ (.A(_05215_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__clkinvlp_2 _11763_ (.A(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__nor2_1 _11764_ (.A(_05218_),
    .B(_05159_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand3_1 _11765_ (.A(_05162_),
    .B(_05078_),
    .C(_05217_),
    .Y(_05220_));
 sky130_fd_sc_hd__o21a_1 _11766_ (.A1(_05164_),
    .A2(net144),
    .B1(_05110_),
    .X(_05221_));
 sky130_fd_sc_hd__nand2_1 _11767_ (.A(_05220_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__nor2_1 _11768_ (.A(_05219_),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__nor2_1 _11769_ (.A(_05094_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__nor2_1 _11770_ (.A(_05213_),
    .B(_05170_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand2_1 _11771_ (.A(_05173_),
    .B(_05218_),
    .Y(_05227_));
 sky130_fd_sc_hd__nand2_1 _11772_ (.A(_05227_),
    .B(_05175_),
    .Y(_05228_));
 sky130_fd_sc_hd__mux2_1 _11773_ (.A0(_05218_),
    .A1(net144),
    .S(_05120_),
    .X(_05229_));
 sky130_fd_sc_hd__o21a_1 _11774_ (.A1(_05177_),
    .A2(_05229_),
    .B1(_05072_),
    .X(_05230_));
 sky130_fd_sc_hd__o21ai_1 _11775_ (.A1(_05226_),
    .A2(_05228_),
    .B1(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand2_1 _11776_ (.A(_05224_),
    .B(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__nor2_1 _11777_ (.A(net144),
    .B(_05182_),
    .Y(_05233_));
 sky130_fd_sc_hd__inv_2 _11778_ (.A(net145),
    .Y(_05234_));
 sky130_fd_sc_hd__nand2_1 _11779_ (.A(_05232_),
    .B(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__or2_1 _11780_ (.A(_01277_),
    .B(_05235_),
    .X(_05237_));
 sky130_fd_sc_hd__inv_2 _11781_ (.A(_05237_),
    .Y(_00029_));
 sky130_fd_sc_hd__inv_2 _11782_ (.A(net156),
    .Y(_05238_));
 sky130_fd_sc_hd__or2_2 _11783_ (.A(_05238_),
    .B(_05215_),
    .X(_05239_));
 sky130_fd_sc_hd__nand2_1 _11784_ (.A(_05215_),
    .B(_05238_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand2_1 _11785_ (.A(_05239_),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hd__clkinvlp_2 _11786_ (.A(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__nor2_1 _11787_ (.A(_05242_),
    .B(_05159_),
    .Y(_05243_));
 sky130_fd_sc_hd__nand3_1 _11788_ (.A(_05162_),
    .B(_05078_),
    .C(_05241_),
    .Y(_05244_));
 sky130_fd_sc_hd__o21a_1 _11789_ (.A1(_05164_),
    .A2(net156),
    .B1(_05110_),
    .X(_05245_));
 sky130_fd_sc_hd__nand2_1 _11790_ (.A(_05244_),
    .B(_05245_),
    .Y(_05247_));
 sky130_fd_sc_hd__nor2_1 _11791_ (.A(_05243_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__nor2_1 _11792_ (.A(_05094_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__nor2_1 _11793_ (.A(_05238_),
    .B(_05170_),
    .Y(_05250_));
 sky130_fd_sc_hd__nand2_1 _11794_ (.A(_05124_),
    .B(_05242_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_1 _11795_ (.A(_05251_),
    .B(_05175_),
    .Y(_05252_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(_05242_),
    .A1(net156),
    .S(_05061_),
    .X(_05253_));
 sky130_fd_sc_hd__o21a_1 _11797_ (.A1(_05177_),
    .A2(_05253_),
    .B1(_05072_),
    .X(_05254_));
 sky130_fd_sc_hd__o21ai_1 _11798_ (.A1(_05250_),
    .A2(_05252_),
    .B1(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__nand2_1 _11799_ (.A(_05249_),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__nor2_1 _11800_ (.A(net156),
    .B(_05182_),
    .Y(_05258_));
 sky130_fd_sc_hd__inv_2 _11801_ (.A(net157),
    .Y(_05259_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(_05256_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__or2_1 _11803_ (.A(_01277_),
    .B(_05260_),
    .X(_05261_));
 sky130_fd_sc_hd__inv_2 _11804_ (.A(_05261_),
    .Y(_00030_));
 sky130_fd_sc_hd__clkbuf_2 _11805_ (.A(net137),
    .X(_05262_));
 sky130_fd_sc_hd__inv_1 _11806_ (.A(net167),
    .Y(_05263_));
 sky130_fd_sc_hd__or2_1 _11807_ (.A(_05263_),
    .B(_05239_),
    .X(_05264_));
 sky130_fd_sc_hd__nand2_1 _11808_ (.A(_05239_),
    .B(_05263_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_1 _11809_ (.A(_05264_),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__clkinvlp_2 _11810_ (.A(_05266_),
    .Y(_05268_));
 sky130_fd_sc_hd__nor2_1 _11811_ (.A(_05268_),
    .B(_05158_),
    .Y(_05269_));
 sky130_fd_sc_hd__nand3_1 _11812_ (.A(_05074_),
    .B(_05106_),
    .C(_05266_),
    .Y(_05270_));
 sky130_fd_sc_hd__o21a_1 _11813_ (.A1(_05075_),
    .A2(net167),
    .B1(_05080_),
    .X(_05271_));
 sky130_fd_sc_hd__nand2_1 _11814_ (.A(_05270_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__o21a_1 _11815_ (.A1(_05269_),
    .A2(_05272_),
    .B1(_05087_),
    .X(_05273_));
 sky130_fd_sc_hd__nor2_1 _11816_ (.A(_05263_),
    .B(_05173_),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2_1 _11817_ (.A(_05124_),
    .B(_05268_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_1 _11818_ (.A(_05275_),
    .B(_05095_),
    .Y(_05276_));
 sky130_fd_sc_hd__mux2_1 _11819_ (.A0(_05268_),
    .A1(net167),
    .S(_05061_),
    .X(_05277_));
 sky130_fd_sc_hd__o21a_1 _11820_ (.A1(_05058_),
    .A2(_05277_),
    .B1(_05072_),
    .X(_05279_));
 sky130_fd_sc_hd__o21ai_1 _11821_ (.A1(_05274_),
    .A2(_05276_),
    .B1(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__nand2_1 _11822_ (.A(_05273_),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__nor2_1 _11823_ (.A(net167),
    .B(_05182_),
    .Y(_05282_));
 sky130_fd_sc_hd__inv_2 _11824_ (.A(net168),
    .Y(_05283_));
 sky130_fd_sc_hd__nand2_1 _11825_ (.A(_05281_),
    .B(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__or2_1 _11826_ (.A(_05262_),
    .B(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__inv_2 _11827_ (.A(_05285_),
    .Y(_00031_));
 sky130_fd_sc_hd__inv_2 _11828_ (.A(net169),
    .Y(_05286_));
 sky130_fd_sc_hd__nor2_1 _11829_ (.A(_05286_),
    .B(_05264_),
    .Y(_05287_));
 sky130_fd_sc_hd__inv_2 _11830_ (.A(_05287_),
    .Y(_05289_));
 sky130_fd_sc_hd__nand2_1 _11831_ (.A(_05264_),
    .B(_05286_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand2_1 _11832_ (.A(_05289_),
    .B(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__clkinvlp_2 _11833_ (.A(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nor2_1 _11834_ (.A(_05292_),
    .B(_05158_),
    .Y(_05293_));
 sky130_fd_sc_hd__nand3_1 _11835_ (.A(_05074_),
    .B(_05106_),
    .C(_05291_),
    .Y(_05294_));
 sky130_fd_sc_hd__o21a_1 _11836_ (.A1(_05075_),
    .A2(net169),
    .B1(_05080_),
    .X(_05295_));
 sky130_fd_sc_hd__nand2_1 _11837_ (.A(_05294_),
    .B(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__o21a_1 _11838_ (.A1(_05293_),
    .A2(_05296_),
    .B1(_05087_),
    .X(_05297_));
 sky130_fd_sc_hd__nor2_1 _11839_ (.A(_05286_),
    .B(_05173_),
    .Y(_05298_));
 sky130_fd_sc_hd__nand2_1 _11840_ (.A(_05124_),
    .B(_05292_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _11841_ (.A(_05300_),
    .B(_05095_),
    .Y(_05301_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(_05292_),
    .A1(net169),
    .S(_05061_),
    .X(_05302_));
 sky130_fd_sc_hd__o21a_1 _11843_ (.A1(_05058_),
    .A2(_05302_),
    .B1(_05072_),
    .X(_05303_));
 sky130_fd_sc_hd__o21ai_1 _11844_ (.A1(_05298_),
    .A2(_05301_),
    .B1(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__nand2_1 _11845_ (.A(_05297_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__nor2_1 _11846_ (.A(net169),
    .B(_05086_),
    .Y(_05306_));
 sky130_fd_sc_hd__inv_2 _11847_ (.A(net170),
    .Y(_05307_));
 sky130_fd_sc_hd__nand2_1 _11848_ (.A(_05305_),
    .B(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__or2_1 _11849_ (.A(_05262_),
    .B(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__inv_2 _11850_ (.A(_05309_),
    .Y(_00032_));
 sky130_fd_sc_hd__inv_1 _11851_ (.A(net171),
    .Y(_05311_));
 sky130_fd_sc_hd__nand2_1 _11852_ (.A(net167),
    .B(net169),
    .Y(_05312_));
 sky130_fd_sc_hd__or2_1 _11853_ (.A(_05312_),
    .B(_05239_),
    .X(_05313_));
 sky130_fd_sc_hd__nor2_1 _11854_ (.A(_05311_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__inv_2 _11855_ (.A(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_1 _11856_ (.A(_05313_),
    .B(_05311_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand2_1 _11857_ (.A(_05315_),
    .B(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__inv_2 _11858_ (.A(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__nor2_1 _11859_ (.A(_05318_),
    .B(_05158_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand3_1 _11860_ (.A(_05074_),
    .B(_05164_),
    .C(_05317_),
    .Y(_05321_));
 sky130_fd_sc_hd__o21a_1 _11861_ (.A1(net146),
    .A2(net171),
    .B1(_05070_),
    .X(_05322_));
 sky130_fd_sc_hd__nand2_1 _11862_ (.A(_05321_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__o21a_1 _11863_ (.A1(_05319_),
    .A2(_05323_),
    .B1(_05086_),
    .X(_05324_));
 sky130_fd_sc_hd__nand2_1 _11864_ (.A(_05052_),
    .B(_05318_),
    .Y(_05325_));
 sky130_fd_sc_hd__o211ai_1 _11865_ (.A1(_05311_),
    .A2(_05052_),
    .B1(_05177_),
    .C1(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__nand2_1 _11866_ (.A(_05318_),
    .B(_05063_),
    .Y(_05327_));
 sky130_fd_sc_hd__a21oi_1 _11867_ (.A1(_05120_),
    .A2(net171),
    .B1(_05057_),
    .Y(_05328_));
 sky130_fd_sc_hd__a21oi_1 _11868_ (.A1(_05327_),
    .A2(_05328_),
    .B1(_05110_),
    .Y(_05329_));
 sky130_fd_sc_hd__nand2_1 _11869_ (.A(_05326_),
    .B(net224),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _11870_ (.A(_05324_),
    .B(_05330_),
    .Y(_05332_));
 sky130_fd_sc_hd__nor2_1 _11871_ (.A(net171),
    .B(_05086_),
    .Y(_05333_));
 sky130_fd_sc_hd__inv_2 _11872_ (.A(net172),
    .Y(_05334_));
 sky130_fd_sc_hd__nand2_2 _11873_ (.A(_05332_),
    .B(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__or2_1 _11874_ (.A(_05262_),
    .B(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__inv_2 _11875_ (.A(_05336_),
    .Y(_00003_));
 sky130_fd_sc_hd__nor2_1 _11876_ (.A(net176),
    .B(_05314_),
    .Y(_05337_));
 sky130_fd_sc_hd__nor2_1 _11877_ (.A(_05311_),
    .B(_05289_),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _11878_ (.A(_05338_),
    .B(net176),
    .Y(_05339_));
 sky130_fd_sc_hd__inv_2 _11879_ (.A(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__nor2_1 _11880_ (.A(_05337_),
    .B(_05340_),
    .Y(_05342_));
 sky130_fd_sc_hd__nor2_1 _11881_ (.A(_05342_),
    .B(_05159_),
    .Y(_05343_));
 sky130_fd_sc_hd__clkinvlp_2 _11882_ (.A(_05342_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand3_1 _11883_ (.A(_05162_),
    .B(_05078_),
    .C(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__o21a_1 _11884_ (.A1(_05164_),
    .A2(net176),
    .B1(_05080_),
    .X(_05346_));
 sky130_fd_sc_hd__nand2_1 _11885_ (.A(_05345_),
    .B(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__nor2_1 _11886_ (.A(_05343_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__nor2_1 _11887_ (.A(_05085_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__inv_1 _11888_ (.A(net176),
    .Y(_05350_));
 sky130_fd_sc_hd__nor2_1 _11889_ (.A(_05350_),
    .B(_05173_),
    .Y(_05351_));
 sky130_fd_sc_hd__nand2_1 _11890_ (.A(_05124_),
    .B(_05342_),
    .Y(_05353_));
 sky130_fd_sc_hd__nand2_1 _11891_ (.A(_05353_),
    .B(_05095_),
    .Y(_05354_));
 sky130_fd_sc_hd__nor2_1 _11892_ (.A(_05350_),
    .B(_05062_),
    .Y(_05355_));
 sky130_fd_sc_hd__nor2_1 _11893_ (.A(_05120_),
    .B(_05344_),
    .Y(_05356_));
 sky130_fd_sc_hd__o31a_1 _11894_ (.A1(_05058_),
    .A2(_05355_),
    .A3(_05356_),
    .B1(_05071_),
    .X(_05357_));
 sky130_fd_sc_hd__o21ai_1 _11895_ (.A1(_05351_),
    .A2(_05354_),
    .B1(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand2_1 _11896_ (.A(_05349_),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__nor2_1 _11897_ (.A(net176),
    .B(_05086_),
    .Y(_05360_));
 sky130_fd_sc_hd__inv_2 _11898_ (.A(net177),
    .Y(_05361_));
 sky130_fd_sc_hd__nand2_1 _11899_ (.A(_05359_),
    .B(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__or2_1 _11900_ (.A(_05262_),
    .B(_05362_),
    .X(_05364_));
 sky130_fd_sc_hd__inv_2 _11901_ (.A(_05364_),
    .Y(_00004_));
 sky130_fd_sc_hd__inv_2 _11902_ (.A(net178),
    .Y(_05365_));
 sky130_fd_sc_hd__or3_1 _11903_ (.A(_05311_),
    .B(_05350_),
    .C(_05312_),
    .X(_05366_));
 sky130_fd_sc_hd__or2_1 _11904_ (.A(_05366_),
    .B(_05239_),
    .X(_05367_));
 sky130_fd_sc_hd__nor2_1 _11905_ (.A(_05365_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__nand2_1 _11906_ (.A(_05367_),
    .B(_05365_),
    .Y(_05369_));
 sky130_fd_sc_hd__inv_2 _11907_ (.A(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__nor2_2 _11908_ (.A(_05368_),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__nor2_1 _11909_ (.A(_05371_),
    .B(_05159_),
    .Y(_05372_));
 sky130_fd_sc_hd__clkinvlp_2 _11910_ (.A(_05371_),
    .Y(_05374_));
 sky130_fd_sc_hd__nand3_1 _11911_ (.A(_05162_),
    .B(_05106_),
    .C(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__o21a_1 _11912_ (.A1(_05164_),
    .A2(net178),
    .B1(_05080_),
    .X(_05376_));
 sky130_fd_sc_hd__nand2_1 _11913_ (.A(_05375_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__o21a_1 _11914_ (.A1(_05372_),
    .A2(_05377_),
    .B1(_05087_),
    .X(_05378_));
 sky130_fd_sc_hd__nand2_1 _11915_ (.A(_05170_),
    .B(_05371_),
    .Y(_05379_));
 sky130_fd_sc_hd__o211ai_1 _11916_ (.A1(_05365_),
    .A2(_05170_),
    .B1(_05175_),
    .C1(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_05371_),
    .B(_05063_),
    .Y(_05381_));
 sky130_fd_sc_hd__a21oi_1 _11918_ (.A1(_05121_),
    .A2(net178),
    .B1(_05177_),
    .Y(_05382_));
 sky130_fd_sc_hd__a21oi_1 _11919_ (.A1(_05381_),
    .A2(_05382_),
    .B1(_05081_),
    .Y(_05383_));
 sky130_fd_sc_hd__nand2_1 _11920_ (.A(_05380_),
    .B(_05383_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand2_1 _11921_ (.A(_05378_),
    .B(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__nor2_1 _11922_ (.A(net178),
    .B(_05182_),
    .Y(_05387_));
 sky130_fd_sc_hd__inv_2 _11923_ (.A(net179),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _11924_ (.A(_05386_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__or2_1 _11925_ (.A(_05262_),
    .B(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__inv_2 _11926_ (.A(_05390_),
    .Y(_00005_));
 sky130_fd_sc_hd__nor2_1 _11927_ (.A(_05365_),
    .B(_05339_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _11928_ (.A(_05391_),
    .B(net180),
    .Y(_05392_));
 sky130_fd_sc_hd__or2_1 _11929_ (.A(net180),
    .B(_05368_),
    .X(_05393_));
 sky130_fd_sc_hd__and2_1 _11930_ (.A(_05392_),
    .B(_05393_),
    .X(_05395_));
 sky130_fd_sc_hd__nor2_1 _11931_ (.A(_05395_),
    .B(_05158_),
    .Y(_05396_));
 sky130_fd_sc_hd__o21a_1 _11932_ (.A1(net146),
    .A2(net180),
    .B1(_05070_),
    .X(_05397_));
 sky130_fd_sc_hd__o21ai_1 _11933_ (.A1(_05395_),
    .A2(_05076_),
    .B1(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__o21a_1 _11934_ (.A1(_05396_),
    .A2(_05398_),
    .B1(_05086_),
    .X(_05399_));
 sky130_fd_sc_hd__clkinvlp_2 _11935_ (.A(net180),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_1 _11936_ (.A(_05052_),
    .B(_05395_),
    .Y(_05401_));
 sky130_fd_sc_hd__o211ai_1 _11937_ (.A1(net181),
    .A2(_05052_),
    .B1(_05177_),
    .C1(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__nand2_1 _11938_ (.A(_05395_),
    .B(_05062_),
    .Y(_05403_));
 sky130_fd_sc_hd__a21oi_1 _11939_ (.A1(_05120_),
    .A2(net180),
    .B1(_05057_),
    .Y(_05404_));
 sky130_fd_sc_hd__a21oi_1 _11940_ (.A1(_05403_),
    .A2(_05404_),
    .B1(_05110_),
    .Y(_05406_));
 sky130_fd_sc_hd__nand2_1 _11941_ (.A(_05402_),
    .B(net231),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_1 _11942_ (.A(_05399_),
    .B(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_1 _11943_ (.A(_05085_),
    .B(net181),
    .Y(_05409_));
 sky130_fd_sc_hd__nand2_1 _11944_ (.A(_05408_),
    .B(_05409_),
    .Y(_05410_));
 sky130_fd_sc_hd__or2_1 _11945_ (.A(_05262_),
    .B(_05410_),
    .X(_05411_));
 sky130_fd_sc_hd__inv_2 _11946_ (.A(_05411_),
    .Y(_00006_));
 sky130_fd_sc_hd__inv_2 _11947_ (.A(net173),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _11948_ (.A(_05392_),
    .B(net174),
    .Y(_05413_));
 sky130_fd_sc_hd__nand2_1 _11949_ (.A(net178),
    .B(net180),
    .Y(_05414_));
 sky130_fd_sc_hd__or3_1 _11950_ (.A(net174),
    .B(_05414_),
    .C(_05367_),
    .X(_05416_));
 sky130_fd_sc_hd__nand2_1 _11951_ (.A(_05413_),
    .B(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__inv_2 _11952_ (.A(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__nor2_1 _11953_ (.A(_05418_),
    .B(_05158_),
    .Y(_05419_));
 sky130_fd_sc_hd__o21a_1 _11954_ (.A1(net146),
    .A2(net173),
    .B1(_05070_),
    .X(_05420_));
 sky130_fd_sc_hd__o21ai_1 _11955_ (.A1(_05418_),
    .A2(_05076_),
    .B1(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__nor2_1 _11956_ (.A(_05419_),
    .B(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__nor2_1 _11957_ (.A(_05085_),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__nand2_1 _11958_ (.A(_05051_),
    .B(_05418_),
    .Y(_05424_));
 sky130_fd_sc_hd__o211ai_1 _11959_ (.A1(net174),
    .A2(_05051_),
    .B1(_05058_),
    .C1(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _11960_ (.A(_05418_),
    .B(_05062_),
    .Y(_05427_));
 sky130_fd_sc_hd__a21oi_1 _11961_ (.A1(_05120_),
    .A2(net173),
    .B1(_05057_),
    .Y(_05428_));
 sky130_fd_sc_hd__a21oi_1 _11962_ (.A1(_05427_),
    .A2(_05428_),
    .B1(_05110_),
    .Y(_05429_));
 sky130_fd_sc_hd__nand2_1 _11963_ (.A(_05425_),
    .B(net214),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _11964_ (.A(_05423_),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__nand2_1 _11965_ (.A(_05085_),
    .B(net174),
    .Y(_05432_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(_05431_),
    .B(net175),
    .Y(_05433_));
 sky130_fd_sc_hd__or2_1 _11967_ (.A(_05262_),
    .B(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__inv_2 _11968_ (.A(_05434_),
    .Y(_00007_));
 sky130_fd_sc_hd__inv_2 _11969_ (.A(net187),
    .Y(_05435_));
 sky130_fd_sc_hd__or3_1 _11970_ (.A(net174),
    .B(net188),
    .C(_05392_),
    .X(_05437_));
 sky130_fd_sc_hd__nand2_1 _11971_ (.A(_05416_),
    .B(net188),
    .Y(_05438_));
 sky130_fd_sc_hd__nand2_1 _11972_ (.A(_05437_),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__clkinvlp_2 _11973_ (.A(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__nor2_1 _11974_ (.A(_05440_),
    .B(_05158_),
    .Y(_05441_));
 sky130_fd_sc_hd__o21a_1 _11975_ (.A1(_05075_),
    .A2(net187),
    .B1(_05070_),
    .X(_05442_));
 sky130_fd_sc_hd__o21ai_1 _11976_ (.A1(_05440_),
    .A2(_05076_),
    .B1(net220),
    .Y(_05443_));
 sky130_fd_sc_hd__o21a_1 _11977_ (.A1(_05441_),
    .A2(_05443_),
    .B1(_05086_),
    .X(_05444_));
 sky130_fd_sc_hd__nand2_1 _11978_ (.A(_05052_),
    .B(_05440_),
    .Y(_05445_));
 sky130_fd_sc_hd__o211ai_1 _11979_ (.A1(net188),
    .A2(_05124_),
    .B1(_05095_),
    .C1(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__nor2_1 _11980_ (.A(net188),
    .B(_05062_),
    .Y(_05448_));
 sky130_fd_sc_hd__nor2_1 _11981_ (.A(_05120_),
    .B(_05439_),
    .Y(_05449_));
 sky130_fd_sc_hd__o31a_1 _11982_ (.A1(_05057_),
    .A2(_05448_),
    .A3(_05449_),
    .B1(_05071_),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_1 _11983_ (.A(_05446_),
    .B(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__nand2_1 _11984_ (.A(_05444_),
    .B(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__nand2_1 _11985_ (.A(_05094_),
    .B(net188),
    .Y(_05453_));
 sky130_fd_sc_hd__nand2_1 _11986_ (.A(_05452_),
    .B(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__or2_1 _11987_ (.A(_05262_),
    .B(_05454_),
    .X(_05455_));
 sky130_fd_sc_hd__inv_2 _11988_ (.A(_05455_),
    .Y(_00008_));
 sky130_fd_sc_hd__or4_1 _11989_ (.A(net174),
    .B(_05435_),
    .C(_05414_),
    .D(_05366_),
    .X(_05456_));
 sky130_fd_sc_hd__nor2_2 _11990_ (.A(_05239_),
    .B(_05456_),
    .Y(_05458_));
 sky130_fd_sc_hd__or2_1 _11991_ (.A(\M00r[18] ),
    .B(_05458_),
    .X(_05459_));
 sky130_fd_sc_hd__nand2_1 _11992_ (.A(_05458_),
    .B(\M00r[18] ),
    .Y(_05460_));
 sky130_fd_sc_hd__nand2_1 _11993_ (.A(_05459_),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__inv_2 _11994_ (.A(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__nor2_1 _11995_ (.A(_05462_),
    .B(_05159_),
    .Y(_05463_));
 sky130_fd_sc_hd__nand3_1 _11996_ (.A(_05162_),
    .B(_05078_),
    .C(_05461_),
    .Y(_05464_));
 sky130_fd_sc_hd__o21a_1 _11997_ (.A1(_05164_),
    .A2(\M00r[18] ),
    .B1(_05080_),
    .X(_05465_));
 sky130_fd_sc_hd__nand2_1 _11998_ (.A(_05464_),
    .B(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__nor2_1 _11999_ (.A(_05463_),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__nor2_1 _12000_ (.A(_05085_),
    .B(_05467_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_1 _12001_ (.A(_05200_),
    .B(\M00r[18] ),
    .Y(_05470_));
 sky130_fd_sc_hd__nand2_1 _12002_ (.A(net102),
    .B(_05462_),
    .Y(_05471_));
 sky130_fd_sc_hd__nand3_1 _12003_ (.A(_05470_),
    .B(_05175_),
    .C(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_1 _12004_ (.A(_05462_),
    .B(_05063_),
    .Y(_05473_));
 sky130_fd_sc_hd__a21oi_1 _12005_ (.A1(_05121_),
    .A2(\M00r[18] ),
    .B1(_05177_),
    .Y(_05474_));
 sky130_fd_sc_hd__a21oi_1 _12006_ (.A1(_05473_),
    .A2(_05474_),
    .B1(_05081_),
    .Y(_05475_));
 sky130_fd_sc_hd__nand2_1 _12007_ (.A(_05472_),
    .B(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _12008_ (.A(_05469_),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__nor2_1 _12009_ (.A(\M00r[18] ),
    .B(_05182_),
    .Y(_05478_));
 sky130_fd_sc_hd__inv_2 _12010_ (.A(_05478_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2_1 _12011_ (.A(_05477_),
    .B(net186),
    .Y(_05481_));
 sky130_fd_sc_hd__or2_1 _12012_ (.A(_05262_),
    .B(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__inv_2 _12013_ (.A(_05482_),
    .Y(_00009_));
 sky130_fd_sc_hd__inv_2 _12014_ (.A(net182),
    .Y(_05483_));
 sky130_fd_sc_hd__nand2_1 _12015_ (.A(_05460_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__nand2_1 _12016_ (.A(\M00r[18] ),
    .B(net182),
    .Y(_05485_));
 sky130_fd_sc_hd__inv_2 _12017_ (.A(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand2_1 _12018_ (.A(_05458_),
    .B(net196),
    .Y(_05487_));
 sky130_fd_sc_hd__nand2_1 _12019_ (.A(net248),
    .B(net197),
    .Y(_05488_));
 sky130_fd_sc_hd__clkinvlp_2 _12020_ (.A(net198),
    .Y(_05490_));
 sky130_fd_sc_hd__nor2_1 _12021_ (.A(_05490_),
    .B(_05158_),
    .Y(_05491_));
 sky130_fd_sc_hd__nand3_1 _12022_ (.A(_05074_),
    .B(_05106_),
    .C(net198),
    .Y(_05492_));
 sky130_fd_sc_hd__o21a_1 _12023_ (.A1(_05075_),
    .A2(net182),
    .B1(_05080_),
    .X(_05493_));
 sky130_fd_sc_hd__nand2_1 _12024_ (.A(_05492_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__o21a_1 _12025_ (.A1(_05491_),
    .A2(_05494_),
    .B1(_05087_),
    .X(_05495_));
 sky130_fd_sc_hd__nor2_1 _12026_ (.A(_05483_),
    .B(_05173_),
    .Y(_05496_));
 sky130_fd_sc_hd__nand2_1 _12027_ (.A(_05124_),
    .B(_05490_),
    .Y(_05497_));
 sky130_fd_sc_hd__nand2_1 _12028_ (.A(_05497_),
    .B(_05175_),
    .Y(_05498_));
 sky130_fd_sc_hd__nand2_1 _12029_ (.A(_05490_),
    .B(_05063_),
    .Y(_05499_));
 sky130_fd_sc_hd__a21oi_1 _12030_ (.A1(_05121_),
    .A2(net182),
    .B1(_05058_),
    .Y(_05501_));
 sky130_fd_sc_hd__a21oi_1 _12031_ (.A1(_05499_),
    .A2(_05501_),
    .B1(_05081_),
    .Y(_05502_));
 sky130_fd_sc_hd__o21ai_1 _12032_ (.A1(_05496_),
    .A2(_05498_),
    .B1(_05502_),
    .Y(_05503_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_05495_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__nor2_1 _12034_ (.A(net182),
    .B(_05182_),
    .Y(_05505_));
 sky130_fd_sc_hd__inv_2 _12035_ (.A(net183),
    .Y(_05506_));
 sky130_fd_sc_hd__nand2_1 _12036_ (.A(_05504_),
    .B(_05506_),
    .Y(_05507_));
 sky130_fd_sc_hd__or2_1 _12037_ (.A(_05262_),
    .B(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__inv_2 _12038_ (.A(_05508_),
    .Y(_00010_));
 sky130_fd_sc_hd__clkinvlp_2 _12039_ (.A(net160),
    .Y(_05509_));
 sky130_fd_sc_hd__or2_1 _12040_ (.A(_05509_),
    .B(net197),
    .X(_05511_));
 sky130_fd_sc_hd__nand2_1 _12041_ (.A(net197),
    .B(_05509_),
    .Y(_05512_));
 sky130_fd_sc_hd__nand2_1 _12042_ (.A(_05511_),
    .B(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hd__inv_2 _12043_ (.A(_05513_),
    .Y(_05514_));
 sky130_fd_sc_hd__nor2_1 _12044_ (.A(_05514_),
    .B(_05159_),
    .Y(_05515_));
 sky130_fd_sc_hd__nand3_1 _12045_ (.A(_05162_),
    .B(_05078_),
    .C(_05513_),
    .Y(_05516_));
 sky130_fd_sc_hd__o21a_1 _12046_ (.A1(_05164_),
    .A2(net160),
    .B1(_05110_),
    .X(_05517_));
 sky130_fd_sc_hd__nand2_1 _12047_ (.A(_05516_),
    .B(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__nor2_1 _12048_ (.A(_05515_),
    .B(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__nor2_1 _12049_ (.A(_05085_),
    .B(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__nand2_1 _12050_ (.A(_05200_),
    .B(net160),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_1 _12051_ (.A(net102),
    .B(_05514_),
    .Y(_05523_));
 sky130_fd_sc_hd__nand3_1 _12052_ (.A(_05522_),
    .B(_05175_),
    .C(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__nand2_1 _12053_ (.A(_05514_),
    .B(_05063_),
    .Y(_05525_));
 sky130_fd_sc_hd__a21oi_1 _12054_ (.A1(_05121_),
    .A2(net160),
    .B1(_05177_),
    .Y(_05526_));
 sky130_fd_sc_hd__a21oi_1 _12055_ (.A1(_05525_),
    .A2(_05526_),
    .B1(_05081_),
    .Y(_05527_));
 sky130_fd_sc_hd__nand2_1 _12056_ (.A(_05524_),
    .B(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _12057_ (.A(_05520_),
    .B(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__nor2_1 _12058_ (.A(net160),
    .B(_05182_),
    .Y(_05530_));
 sky130_fd_sc_hd__inv_2 _12059_ (.A(net161),
    .Y(_05531_));
 sky130_fd_sc_hd__nand2_1 _12060_ (.A(_05529_),
    .B(_05531_),
    .Y(_05533_));
 sky130_fd_sc_hd__or2_1 _12061_ (.A(net133),
    .B(_05533_),
    .X(_05534_));
 sky130_fd_sc_hd__inv_2 _12062_ (.A(_05534_),
    .Y(_00011_));
 sky130_fd_sc_hd__clkinvlp_2 _12063_ (.A(net164),
    .Y(_05535_));
 sky130_fd_sc_hd__inv_2 _12064_ (.A(\M00r[18] ),
    .Y(_05536_));
 sky130_fd_sc_hd__or3_1 _12065_ (.A(_05536_),
    .B(_05483_),
    .C(_05437_),
    .X(_05537_));
 sky130_fd_sc_hd__or3_1 _12066_ (.A(_05509_),
    .B(_05535_),
    .C(net206),
    .X(_05538_));
 sky130_fd_sc_hd__nand2_1 _12067_ (.A(_05511_),
    .B(_05535_),
    .Y(_05539_));
 sky130_fd_sc_hd__nand2_1 _12068_ (.A(net207),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__inv_2 _12069_ (.A(net208),
    .Y(_05541_));
 sky130_fd_sc_hd__nor2_1 _12070_ (.A(_05541_),
    .B(_05159_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand3_1 _12071_ (.A(_05162_),
    .B(_05106_),
    .C(net208),
    .Y(_05544_));
 sky130_fd_sc_hd__o21a_1 _12072_ (.A1(_05075_),
    .A2(net164),
    .B1(_05080_),
    .X(_05545_));
 sky130_fd_sc_hd__nand2_1 _12073_ (.A(_05544_),
    .B(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21a_1 _12074_ (.A1(_05543_),
    .A2(_05546_),
    .B1(_05087_),
    .X(_05547_));
 sky130_fd_sc_hd__nand2_1 _12075_ (.A(net102),
    .B(_05541_),
    .Y(_05548_));
 sky130_fd_sc_hd__o211ai_1 _12076_ (.A1(_05535_),
    .A2(_05170_),
    .B1(_05175_),
    .C1(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__nand2_1 _12077_ (.A(_05541_),
    .B(_05063_),
    .Y(_05550_));
 sky130_fd_sc_hd__a21oi_1 _12078_ (.A1(_05121_),
    .A2(net164),
    .B1(_05177_),
    .Y(_05551_));
 sky130_fd_sc_hd__a21oi_1 _12079_ (.A1(_05550_),
    .A2(_05551_),
    .B1(_05081_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand2_1 _12080_ (.A(_05549_),
    .B(_05552_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(_05547_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__nor2_1 _12082_ (.A(net164),
    .B(_05182_),
    .Y(_05556_));
 sky130_fd_sc_hd__inv_2 _12083_ (.A(net165),
    .Y(_05557_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(_05555_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__or2_1 _12085_ (.A(net133),
    .B(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__inv_2 _12086_ (.A(_05559_),
    .Y(_00012_));
 sky130_fd_sc_hd__and4_1 _12087_ (.A(_05458_),
    .B(net160),
    .C(net164),
    .D(net196),
    .X(_05560_));
 sky130_fd_sc_hd__or2_1 _12088_ (.A(net166),
    .B(_05560_),
    .X(_05561_));
 sky130_fd_sc_hd__nand2_1 _12089_ (.A(_05560_),
    .B(net166),
    .Y(_05562_));
 sky130_fd_sc_hd__nand2_1 _12090_ (.A(_05561_),
    .B(_05562_),
    .Y(_05564_));
 sky130_fd_sc_hd__inv_2 _12091_ (.A(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__nor2_1 _12092_ (.A(_05565_),
    .B(_05159_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand3_1 _12093_ (.A(_05162_),
    .B(_05078_),
    .C(_05564_),
    .Y(_05567_));
 sky130_fd_sc_hd__o21a_1 _12094_ (.A1(_05164_),
    .A2(net166),
    .B1(_05110_),
    .X(_05568_));
 sky130_fd_sc_hd__nand2_1 _12095_ (.A(_05567_),
    .B(_05568_),
    .Y(_05569_));
 sky130_fd_sc_hd__nor2_1 _12096_ (.A(_05566_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__nor2_1 _12097_ (.A(_05094_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__inv_2 _12098_ (.A(net166),
    .Y(_05572_));
 sky130_fd_sc_hd__nor2_1 _12099_ (.A(_05572_),
    .B(_05170_),
    .Y(_05573_));
 sky130_fd_sc_hd__nand2_1 _12100_ (.A(net102),
    .B(_05565_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand2_1 _12101_ (.A(_05575_),
    .B(_05175_),
    .Y(_05576_));
 sky130_fd_sc_hd__nand2_1 _12102_ (.A(_05565_),
    .B(_05063_),
    .Y(_05577_));
 sky130_fd_sc_hd__a21oi_1 _12103_ (.A1(_05121_),
    .A2(net166),
    .B1(_05177_),
    .Y(_05578_));
 sky130_fd_sc_hd__a21oi_1 _12104_ (.A1(_05577_),
    .A2(_05578_),
    .B1(_05081_),
    .Y(_05579_));
 sky130_fd_sc_hd__o21ai_1 _12105_ (.A1(_05573_),
    .A2(_05576_),
    .B1(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__nand2_1 _12106_ (.A(_05571_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__o21ai_1 _12107_ (.A1(net203),
    .A2(_05089_),
    .B1(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__or2_1 _12108_ (.A(net133),
    .B(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__inv_2 _12109_ (.A(_05583_),
    .Y(_00014_));
 sky130_fd_sc_hd__clkinvlp_2 _12110_ (.A(net162),
    .Y(_05585_));
 sky130_fd_sc_hd__or3_1 _12111_ (.A(_05572_),
    .B(_05585_),
    .C(_05538_),
    .X(_05586_));
 sky130_fd_sc_hd__nand2_1 _12112_ (.A(_05562_),
    .B(_05585_),
    .Y(_05587_));
 sky130_fd_sc_hd__nand2_1 _12113_ (.A(_05586_),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__clkinvlp_2 _12114_ (.A(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__nor2_1 _12115_ (.A(_05589_),
    .B(_05159_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand3_1 _12116_ (.A(_05162_),
    .B(_05078_),
    .C(_05588_),
    .Y(_05591_));
 sky130_fd_sc_hd__o21a_1 _12117_ (.A1(_05164_),
    .A2(net162),
    .B1(_05110_),
    .X(_05592_));
 sky130_fd_sc_hd__nand2_1 _12118_ (.A(_05591_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__nor2_1 _12119_ (.A(_05590_),
    .B(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__nor2_1 _12120_ (.A(_05094_),
    .B(_05594_),
    .Y(_05596_));
 sky130_fd_sc_hd__nor2_1 _12121_ (.A(_05585_),
    .B(_05170_),
    .Y(_05597_));
 sky130_fd_sc_hd__nand2_1 _12122_ (.A(_05170_),
    .B(_05589_),
    .Y(_05598_));
 sky130_fd_sc_hd__nand2_1 _12123_ (.A(_05598_),
    .B(_05175_),
    .Y(_05599_));
 sky130_fd_sc_hd__nand2_1 _12124_ (.A(_05589_),
    .B(_05063_),
    .Y(_05600_));
 sky130_fd_sc_hd__a21oi_1 _12125_ (.A1(_05121_),
    .A2(net162),
    .B1(_05095_),
    .Y(_05601_));
 sky130_fd_sc_hd__a21oi_1 _12126_ (.A1(_05600_),
    .A2(_05601_),
    .B1(_05081_),
    .Y(_05602_));
 sky130_fd_sc_hd__o21ai_1 _12127_ (.A1(_05597_),
    .A2(_05599_),
    .B1(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__nand2_1 _12128_ (.A(_05596_),
    .B(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__nor2_1 _12129_ (.A(net162),
    .B(_05087_),
    .Y(_05605_));
 sky130_fd_sc_hd__inv_2 _12130_ (.A(net163),
    .Y(_05607_));
 sky130_fd_sc_hd__nand2_1 _12131_ (.A(_05604_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__or2_1 _12132_ (.A(net133),
    .B(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__inv_2 _12133_ (.A(_05609_),
    .Y(_00015_));
 sky130_fd_sc_hd__xor2_1 _12134_ (.A(net189),
    .B(_05586_),
    .X(_05610_));
 sky130_fd_sc_hd__clkinvlp_2 _12135_ (.A(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__nor2_1 _12136_ (.A(_05611_),
    .B(_05158_),
    .Y(_05612_));
 sky130_fd_sc_hd__nand3_1 _12137_ (.A(_05074_),
    .B(_05106_),
    .C(_05610_),
    .Y(_05613_));
 sky130_fd_sc_hd__o21a_1 _12138_ (.A1(_05075_),
    .A2(net189),
    .B1(_05080_),
    .X(_05614_));
 sky130_fd_sc_hd__nand2_1 _12139_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__nor2_1 _12140_ (.A(_05612_),
    .B(_05615_),
    .Y(_05617_));
 sky130_fd_sc_hd__nor2_1 _12141_ (.A(_05085_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__inv_2 _12142_ (.A(net189),
    .Y(_05619_));
 sky130_fd_sc_hd__nor2_1 _12143_ (.A(_05619_),
    .B(_05124_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _12144_ (.A(_05124_),
    .B(_05611_),
    .Y(_05621_));
 sky130_fd_sc_hd__nand2_1 _12145_ (.A(_05621_),
    .B(_05095_),
    .Y(_05622_));
 sky130_fd_sc_hd__nand2_1 _12146_ (.A(_05611_),
    .B(_05063_),
    .Y(_05623_));
 sky130_fd_sc_hd__a21oi_1 _12147_ (.A1(_05121_),
    .A2(net189),
    .B1(_05058_),
    .Y(_05624_));
 sky130_fd_sc_hd__a21oi_1 _12148_ (.A1(_05623_),
    .A2(_05624_),
    .B1(_05081_),
    .Y(_05625_));
 sky130_fd_sc_hd__o21ai_1 _12149_ (.A1(_05620_),
    .A2(_05622_),
    .B1(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand2_1 _12150_ (.A(_05618_),
    .B(_05626_),
    .Y(_05628_));
 sky130_fd_sc_hd__nor2_1 _12151_ (.A(net189),
    .B(_05086_),
    .Y(_05629_));
 sky130_fd_sc_hd__inv_2 _12152_ (.A(net190),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_1 _12153_ (.A(_05628_),
    .B(net191),
    .Y(_05631_));
 sky130_fd_sc_hd__nand2_1 _12154_ (.A(_01277_),
    .B(net130),
    .Y(_05632_));
 sky130_fd_sc_hd__o21ai_1 _12155_ (.A1(_01277_),
    .A2(_05631_),
    .B1(net131),
    .Y(_00016_));
 sky130_fd_sc_hd__nand2_1 _12156_ (.A(_05362_),
    .B(net176),
    .Y(_05633_));
 sky130_fd_sc_hd__nand3_1 _12157_ (.A(_05359_),
    .B(_05350_),
    .C(_05089_),
    .Y(_05634_));
 sky130_fd_sc_hd__nand2_1 _12158_ (.A(_05633_),
    .B(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__nand2_1 _12159_ (.A(_05335_),
    .B(net171),
    .Y(_05636_));
 sky130_fd_sc_hd__nand2_1 _12160_ (.A(_05308_),
    .B(net169),
    .Y(_05638_));
 sky130_fd_sc_hd__nand2_1 _12161_ (.A(_05636_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__nor2_1 _12162_ (.A(_05635_),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__nand2_1 _12163_ (.A(_05631_),
    .B(net189),
    .Y(_05641_));
 sky130_fd_sc_hd__nand3_1 _12164_ (.A(_05628_),
    .B(_05619_),
    .C(_05089_),
    .Y(_05642_));
 sky130_fd_sc_hd__nand2_1 _12165_ (.A(_05641_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__nand2_1 _12166_ (.A(_05507_),
    .B(net182),
    .Y(_05644_));
 sky130_fd_sc_hd__nand3_1 _12167_ (.A(_05504_),
    .B(_05483_),
    .C(_05089_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2_1 _12168_ (.A(_05644_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__nor2_1 _12169_ (.A(_05643_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_1 _12170_ (.A(_05640_),
    .B(_05647_),
    .Y(_05649_));
 sky130_fd_sc_hd__nand2_1 _12171_ (.A(_05558_),
    .B(net164),
    .Y(_05650_));
 sky130_fd_sc_hd__buf_6 _12172_ (.A(_05087_),
    .X(_05651_));
 sky130_fd_sc_hd__nand3_1 _12173_ (.A(_05604_),
    .B(_05585_),
    .C(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_1 _12174_ (.A(_05650_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__nand2_1 _12175_ (.A(_05582_),
    .B(net166),
    .Y(_05654_));
 sky130_fd_sc_hd__nand3_1 _12176_ (.A(_05555_),
    .B(_05535_),
    .C(_05651_),
    .Y(_05655_));
 sky130_fd_sc_hd__nand2_1 _12177_ (.A(_05654_),
    .B(_05655_),
    .Y(_05656_));
 sky130_fd_sc_hd__nor2_1 _12178_ (.A(_05653_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand2_1 _12179_ (.A(_05284_),
    .B(net167),
    .Y(_05658_));
 sky130_fd_sc_hd__nand3_1 _12180_ (.A(_05386_),
    .B(_05365_),
    .C(_05089_),
    .Y(_05660_));
 sky130_fd_sc_hd__nand2_1 _12181_ (.A(_05658_),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__nand2_1 _12182_ (.A(_05389_),
    .B(net178),
    .Y(_05662_));
 sky130_fd_sc_hd__nand3_1 _12183_ (.A(_05305_),
    .B(_05286_),
    .C(_05651_),
    .Y(_05663_));
 sky130_fd_sc_hd__nand2_1 _12184_ (.A(_05662_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__nor2_1 _12185_ (.A(_05661_),
    .B(_05664_),
    .Y(_05665_));
 sky130_fd_sc_hd__nand2_1 _12186_ (.A(_05657_),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__nor2_1 _12187_ (.A(_05649_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand3_1 _12188_ (.A(_05431_),
    .B(net174),
    .C(_05089_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21ai_1 _12189_ (.A1(net171),
    .A2(_05335_),
    .B1(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__inv_2 _12190_ (.A(_05669_),
    .Y(_05671_));
 sky130_fd_sc_hd__nand3_1 _12191_ (.A(_05408_),
    .B(net181),
    .C(_05087_),
    .Y(_05672_));
 sky130_fd_sc_hd__nand2_1 _12192_ (.A(_05433_),
    .B(net213),
    .Y(_05673_));
 sky130_fd_sc_hd__nand2_1 _12193_ (.A(_05672_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__inv_2 _12194_ (.A(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_1 _12195_ (.A(_05671_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand2_1 _12196_ (.A(_05410_),
    .B(net180),
    .Y(_05677_));
 sky130_fd_sc_hd__nand3_1 _12197_ (.A(_05452_),
    .B(net188),
    .C(_05089_),
    .Y(_05678_));
 sky130_fd_sc_hd__nand2_1 _12198_ (.A(_05677_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__inv_2 _12199_ (.A(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__a21oi_1 _12200_ (.A1(_05454_),
    .A2(net219),
    .B1(_05170_),
    .Y(_05682_));
 sky130_fd_sc_hd__nand2_1 _12201_ (.A(_05680_),
    .B(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__nor2_1 _12202_ (.A(_05676_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__nand2_1 _12203_ (.A(_05667_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand3_1 _12204_ (.A(_05208_),
    .B(_05188_),
    .C(_05087_),
    .Y(_05686_));
 sky130_fd_sc_hd__inv_2 _12205_ (.A(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__nand2_1 _12206_ (.A(_05186_),
    .B(net154),
    .Y(_05688_));
 sky130_fd_sc_hd__nand2_1 _12207_ (.A(_05211_),
    .B(net152),
    .Y(_05689_));
 sky130_fd_sc_hd__nand2_1 _12208_ (.A(_05688_),
    .B(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__nor2_1 _12209_ (.A(_05687_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__nand3_1 _12210_ (.A(_05181_),
    .B(_05169_),
    .C(_05089_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand3_1 _12211_ (.A(_05232_),
    .B(_05213_),
    .C(_05089_),
    .Y(_05694_));
 sky130_fd_sc_hd__nand2_1 _12212_ (.A(_05693_),
    .B(_05694_),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_1 _12213_ (.A(_05481_),
    .B(\M00r[18] ),
    .Y(_05696_));
 sky130_fd_sc_hd__nand3_1 _12214_ (.A(_05477_),
    .B(_05536_),
    .C(_05651_),
    .Y(_05697_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(_05696_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__nor2_1 _12216_ (.A(_05695_),
    .B(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__nand2_1 _12217_ (.A(_05691_),
    .B(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__nand2_1 _12218_ (.A(_05235_),
    .B(net144),
    .Y(_05701_));
 sky130_fd_sc_hd__nand3_1 _12219_ (.A(_05256_),
    .B(_05238_),
    .C(_05651_),
    .Y(_05702_));
 sky130_fd_sc_hd__nand2_1 _12220_ (.A(_05701_),
    .B(_05702_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_1 _12221_ (.A(_05608_),
    .B(net162),
    .Y(_05705_));
 sky130_fd_sc_hd__nand3_1 _12222_ (.A(_05529_),
    .B(_05509_),
    .C(_05651_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand2_1 _12223_ (.A(_05705_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nor2_1 _12224_ (.A(_05704_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_1 _12225_ (.A(_05533_),
    .B(net160),
    .Y(_05709_));
 sky130_fd_sc_hd__nand3_1 _12226_ (.A(_05581_),
    .B(_05572_),
    .C(_05651_),
    .Y(_05710_));
 sky130_fd_sc_hd__nand2_1 _12227_ (.A(_05709_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__nand3_1 _12228_ (.A(_05281_),
    .B(_05263_),
    .C(_05651_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _12229_ (.A(_05260_),
    .B(net156),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _12230_ (.A(_05712_),
    .B(_05713_),
    .Y(_05715_));
 sky130_fd_sc_hd__nor2_1 _12231_ (.A(_05711_),
    .B(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__nand2_1 _12232_ (.A(_05708_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__nor2_1 _12233_ (.A(_05700_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__inv_2 _12234_ (.A(_05112_),
    .Y(_05719_));
 sky130_fd_sc_hd__nand3_1 _12235_ (.A(_05719_),
    .B(net216),
    .C(_05090_),
    .Y(_05720_));
 sky130_fd_sc_hd__nand3_1 _12236_ (.A(_05112_),
    .B(net159),
    .C(_05090_),
    .Y(_05721_));
 sky130_fd_sc_hd__nand2_1 _12237_ (.A(_05720_),
    .B(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__inv_2 _12238_ (.A(_05134_),
    .Y(_05723_));
 sky130_fd_sc_hd__nand3_1 _12239_ (.A(_05723_),
    .B(_05116_),
    .C(_05090_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand3_1 _12240_ (.A(_05083_),
    .B(net210),
    .C(_05090_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_1 _12241_ (.A(_05724_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__nor2_1 _12242_ (.A(_05722_),
    .B(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__nand3_1 _12243_ (.A(_05134_),
    .B(net227),
    .C(_05090_),
    .Y(_05729_));
 sky130_fd_sc_hd__nand3_1 _12244_ (.A(_05150_),
    .B(_05137_),
    .C(_05651_),
    .Y(_05730_));
 sky130_fd_sc_hd__nand2_1 _12245_ (.A(_05729_),
    .B(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__inv_2 _12246_ (.A(_05150_),
    .Y(_05732_));
 sky130_fd_sc_hd__nand3_1 _12247_ (.A(_05732_),
    .B(net200),
    .C(_05090_),
    .Y(_05733_));
 sky130_fd_sc_hd__o2111ai_1 _12248_ (.A1(_05081_),
    .A2(_05064_),
    .B1(_01298_),
    .C1(_05651_),
    .D1(_05082_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand2_1 _12249_ (.A(_05733_),
    .B(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__nor2_1 _12250_ (.A(_05731_),
    .B(_05735_),
    .Y(_05737_));
 sky130_fd_sc_hd__nand3_1 _12251_ (.A(_05718_),
    .B(_05728_),
    .C(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__nor2_1 _12252_ (.A(_05685_),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__nor2_1 _12253_ (.A(_01277_),
    .B(_05739_),
    .Y(_00000_));
 sky130_fd_sc_hd__nand2_1 _12254_ (.A(_01277_),
    .B(net124),
    .Y(_05740_));
 sky130_fd_sc_hd__inv_2 _12255_ (.A(net125),
    .Y(_00001_));
 sky130_fd_sc_hd__nand2_1 _12256_ (.A(_01277_),
    .B(net127),
    .Y(_05741_));
 sky130_fd_sc_hd__inv_2 _12257_ (.A(net128),
    .Y(_00033_));
 sky130_fd_sc_hd__clkbuf_1 _12258_ (.A(net25),
    .X(_05742_));
 sky130_fd_sc_hd__clkbuf_1 _12259_ (.A(_05742_),
    .X(inv_f_c));
 sky130_fd_sc_hd__inv_2 _12260_ (.A(net25),
    .Y(ov_f_c));
 sky130_fd_sc_hd__nand2_1 _12261_ (.A(\out_f_c[22] ),
    .B(ov_f_c),
    .Y(forward_c));
 sky130_fd_sc_hd__dfrtp_1 _12262_ (.CLK(clknet_3_7__leaf_clk),
    .D(net129),
    .RESET_B(net80),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _12263_ (.CLK(clknet_3_6__leaf_clk),
    .D(net83),
    .RESET_B(net80),
    .Q(net72));
 sky130_fd_sc_hd__conb_1 _12263__83 (.LO(net83));
 sky130_fd_sc_hd__dfrtp_1 _12264_ (.CLK(clknet_3_7__leaf_clk),
    .D(net141),
    .RESET_B(net80),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _12265_ (.CLK(clknet_3_7__leaf_clk),
    .D(net126),
    .RESET_B(net80),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _12266_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00000_),
    .RESET_B(net77),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _12267_ (.CLK(clknet_3_7__leaf_clk),
    .D(ov_f_c),
    .RESET_B(net80),
    .Q(ov_f));
 sky130_fd_sc_hd__dfrtp_1 _12268_ (.CLK(clknet_3_5__leaf_clk),
    .D(\out_f_c[22] ),
    .RESET_B(net81),
    .Q(\out_f[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12269_ (.CLK(clknet_3_7__leaf_clk),
    .D(net84),
    .RESET_B(net81),
    .Q(done0_r));
 sky130_fd_sc_hd__conb_1 _12269__84 (.HI(net84));
 sky130_fd_sc_hd__dfrtp_1 _12270_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[1] ),
    .RESET_B(net75),
    .Q(\M00r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12271_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sq.out[2] ),
    .RESET_B(net77),
    .Q(\M00r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12272_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[3] ),
    .RESET_B(net73),
    .Q(\M00r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12273_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[4] ),
    .RESET_B(net73),
    .Q(\M00r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12274_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[5] ),
    .RESET_B(net73),
    .Q(\M00r[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12275_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[6] ),
    .RESET_B(net74),
    .Q(\M00r[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12276_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[7] ),
    .RESET_B(net73),
    .Q(\M00r[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12277_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[8] ),
    .RESET_B(net73),
    .Q(\M00r[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12278_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[9] ),
    .RESET_B(net73),
    .Q(\M00r[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12279_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[10] ),
    .RESET_B(net74),
    .Q(\M00r[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12280_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[11] ),
    .RESET_B(net74),
    .Q(\M00r[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12281_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[12] ),
    .RESET_B(net73),
    .Q(\M00r[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12282_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[13] ),
    .RESET_B(net73),
    .Q(\M00r[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12283_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[14] ),
    .RESET_B(net74),
    .Q(\M00r[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12284_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[15] ),
    .RESET_B(net74),
    .Q(\M00r[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12285_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[16] ),
    .RESET_B(net75),
    .Q(\M00r[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12286_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[17] ),
    .RESET_B(net73),
    .Q(\M00r[17] ));
 sky130_fd_sc_hd__dfrtp_4 _12287_ (.CLK(clknet_3_3__leaf_clk),
    .D(\sq.out[18] ),
    .RESET_B(net77),
    .Q(\M00r[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12288_ (.CLK(clknet_3_1__leaf_clk),
    .D(\sq.out[19] ),
    .RESET_B(net75),
    .Q(\M00r[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12289_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sq.out[20] ),
    .RESET_B(net77),
    .Q(\M00r[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12290_ (.CLK(clknet_3_0__leaf_clk),
    .D(\sq.out[21] ),
    .RESET_B(net73),
    .Q(\M00r[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12291_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sq.out[22] ),
    .RESET_B(net77),
    .Q(\M00r[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12292_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sq.out[23] ),
    .RESET_B(net77),
    .Q(\M00r[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12293_ (.CLK(clknet_3_4__leaf_clk),
    .D(\sq.out[24] ),
    .RESET_B(net77),
    .Q(\M00r[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12294_ (.CLK(clknet_3_6__leaf_clk),
    .D(inv_f_c),
    .RESET_B(net80),
    .Q(inv_f));
 sky130_fd_sc_hd__dfrtp_1 _12295_ (.CLK(clknet_3_4__leaf_clk),
    .D(forward_c),
    .RESET_B(net77),
    .Q(forward));
 sky130_fd_sc_hd__dfrtp_1 _12296_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00002_),
    .RESET_B(net76),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _12297_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00013_),
    .RESET_B(net76),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _12298_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00024_),
    .RESET_B(net76),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _12299_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00026_),
    .RESET_B(net76),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _12300_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00027_),
    .RESET_B(net76),
    .Q(net65));
 sky130_fd_sc_hd__dfrtp_1 _12301_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00028_),
    .RESET_B(net76),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _12302_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00029_),
    .RESET_B(net76),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _12303_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00030_),
    .RESET_B(net76),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _12304_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00031_),
    .RESET_B(net76),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _12305_ (.CLK(clknet_3_2__leaf_clk),
    .D(_00032_),
    .RESET_B(net76),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _12306_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00003_),
    .RESET_B(net79),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _12307_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00004_),
    .RESET_B(net79),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _12308_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00005_),
    .RESET_B(net77),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _12309_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00006_),
    .RESET_B(net77),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _12310_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00007_),
    .RESET_B(net78),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _12311_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00008_),
    .RESET_B(net78),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_1 _12312_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00009_),
    .RESET_B(net78),
    .Q(net47));
 sky130_fd_sc_hd__dfrtp_1 _12313_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00010_),
    .RESET_B(net78),
    .Q(net48));
 sky130_fd_sc_hd__dfrtp_1 _12314_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00011_),
    .RESET_B(net78),
    .Q(net49));
 sky130_fd_sc_hd__dfrtp_1 _12315_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00012_),
    .RESET_B(net78),
    .Q(net50));
 sky130_fd_sc_hd__dfrtp_1 _12316_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00014_),
    .RESET_B(net81),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _12317_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00015_),
    .RESET_B(net81),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _12318_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00016_),
    .RESET_B(net81),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _12319_ (.CLK(clknet_3_6__leaf_clk),
    .D(_00017_),
    .RESET_B(net81),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _12320_ (.CLK(clknet_3_6__leaf_clk),
    .D(_00018_),
    .RESET_B(net81),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _12321_ (.CLK(clknet_3_6__leaf_clk),
    .D(_00019_),
    .RESET_B(net81),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _12322_ (.CLK(clknet_3_7__leaf_clk),
    .D(net135),
    .RESET_B(net81),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_1 _12323_ (.CLK(clknet_3_6__leaf_clk),
    .D(_00021_),
    .RESET_B(net80),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _12324_ (.CLK(clknet_3_7__leaf_clk),
    .D(_00022_),
    .RESET_B(net80),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _12325_ (.CLK(clknet_3_7__leaf_clk),
    .D(_00023_),
    .RESET_B(net80),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _12326_ (.CLK(clknet_3_7__leaf_clk),
    .D(net138),
    .RESET_B(net80),
    .Q(net63));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(net75),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(net36),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(net79),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net79),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(net36),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(net36),
    .X(net81));
 sky130_fd_sc_hd__conb_1 fp_sqr_82 (.LO(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_05480_),
    .X(net186));
 sky130_fd_sc_hd__buf_1 hold103 (.A(net218),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 hold104 (.A(_05435_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 hold105 (.A(net245),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_05629_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_05630_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net242),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_05487_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_05488_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\M00r[5] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net139),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\M00r[20] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\M00r[22] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net166),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_05537_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_05538_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_05540_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\M00r[2] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net142),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\M00r[23] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\M00r[16] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net173),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_05429_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\M00r[3] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(net158),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\M00r[7] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\M00r[17] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net187),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_05442_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\M00r[6] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\M00r[14] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\M00r[12] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_05329_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\M00r[9] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\M00r[4] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net150),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\M00r[8] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\M00r[11] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\M00r[15] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_05406_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\M00r[13] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\M00r[10] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\out_f[22] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\M00r[19] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\M00r[21] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\M00r[1] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_05486_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\M00r[24] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_05484_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net140),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(inv_f),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_05740_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_00001_),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(ov_f),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_05741_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_00033_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net236),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_05632_),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net136),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 hold49 (.A(_00751_),
    .X(net133));
 sky130_fd_sc_hd__buf_1 hold50 (.A(_00773_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_00020_),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(forward),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net132),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_00025_),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net199),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(done0_r),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net123),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_2 hold58 (.A(net209),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_05091_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_2 hold60 (.A(net228),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_05233_),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 hold62 (.A(net239),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 hold63 (.A(_05050_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_05148_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_05149_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_2 hold66 (.A(net226),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_05135_),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_2 hold68 (.A(net217),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_05209_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_2 hold70 (.A(net221),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_05184_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_2 hold72 (.A(net225),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_05258_),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_2 hold74 (.A(net215),
    .X(net158));
 sky130_fd_sc_hd__buf_1 hold75 (.A(_05093_),
    .X(net159));
 sky130_fd_sc_hd__buf_2 hold76 (.A(net201),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_05530_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 hold78 (.A(net211),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_05605_),
    .X(net163));
 sky130_fd_sc_hd__buf_2 hold80 (.A(net238),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_05556_),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 hold82 (.A(net202),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_2 hold83 (.A(net233),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_05282_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 hold85 (.A(net229),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_05306_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 hold87 (.A(net223),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_05333_),
    .X(net172));
 sky130_fd_sc_hd__buf_1 hold89 (.A(net212),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 hold90 (.A(_05412_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_05432_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_2 hold92 (.A(net232),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_05360_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 hold94 (.A(net222),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_05387_),
    .X(net179));
 sky130_fd_sc_hd__buf_2 hold96 (.A(net230),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_05400_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 hold98 (.A(net237),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_05505_),
    .X(net183));
 sky130_fd_sc_hd__buf_2 input1 (.A(in1[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(in1[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(in1[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(in1[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(in1[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(in1[21]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(in1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(in1[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(in1[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(in1[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(in1[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(in1[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(in1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(in1[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in1[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(in1[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_4 input25 (.A(in1[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(in1[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(in1[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(in1[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(in1[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(in1[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(in1[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(in1[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(in1[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(round_m[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(round_m[1]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_8 input35 (.A(round_m[2]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 input36 (.A(rst),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(in1[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(in1[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(in1[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(in1[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(in1[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(in1[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(done));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(inexact));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(inv));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(out[0]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(out[10]));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .X(out[11]));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(out[12]));
 sky130_fd_sc_hd__buf_2 output44 (.A(net44),
    .X(out[13]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(out[14]));
 sky130_fd_sc_hd__clkbuf_4 output46 (.A(net46),
    .X(out[15]));
 sky130_fd_sc_hd__clkbuf_4 output47 (.A(net47),
    .X(out[16]));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net48),
    .X(out[17]));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net49),
    .X(out[18]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(out[19]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(out[20]));
 sky130_fd_sc_hd__clkbuf_4 output53 (.A(net53),
    .X(out[21]));
 sky130_fd_sc_hd__clkbuf_4 output54 (.A(net54),
    .X(out[22]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(out[23]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(out[24]));
 sky130_fd_sc_hd__clkbuf_4 output57 (.A(net57),
    .X(out[25]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(out[26]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(out[27]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(out[28]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(out[29]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(out[2]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(out[30]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(out[3]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(out[4]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(out[5]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(out[6]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(out[7]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(out[8]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(out[9]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(ov));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(un));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer1 (.A(_03738_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 rebuffer15 (.A(_04956_),
    .X(net99));
 sky130_fd_sc_hd__buf_1 rebuffer16 (.A(_02829_),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 rebuffer19 (.A(_05820_),
    .X(net103));
 sky130_fd_sc_hd__buf_2 rebuffer2 (.A(_05989_),
    .X(net117));
 sky130_fd_sc_hd__buf_1 rebuffer24 (.A(_01639_),
    .X(net108));
 sky130_fd_sc_hd__buf_1 rebuffer25 (.A(net108),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 rebuffer26 (.A(net109),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 rebuffer28 (.A(_00446_),
    .X(net112));
 sky130_fd_sc_hd__buf_6 rebuffer29 (.A(_00446_),
    .X(net113));
 sky130_fd_sc_hd__buf_1 rebuffer3 (.A(_05989_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 rebuffer4 (.A(net87),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(_02357_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 rebuffer8 (.A(_02139_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 rebuffer9 (.A(net92),
    .X(net93));
 sky130_fd_sc_hd__buf_6 split1 (.A(_03090_),
    .X(net85));
 sky130_fd_sc_hd__buf_4 split10 (.A(_03771_),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 split11 (.A(_03834_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 split12 (.A(_05820_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 split13 (.A(_03437_),
    .X(net97));
 sky130_fd_sc_hd__dlymetal6s2s_1 split14 (.A(_01359_),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 split15 (.A(_00295_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 split17 (.A(_04531_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 split18 (.A(_05173_),
    .X(net102));
 sky130_fd_sc_hd__buf_2 split2 (.A(_03436_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 split20 (.A(_00841_),
    .X(net104));
 sky130_fd_sc_hd__buf_2 split21 (.A(_02107_),
    .X(net105));
 sky130_fd_sc_hd__buf_4 split22 (.A(_00088_),
    .X(net106));
 sky130_fd_sc_hd__buf_2 split23 (.A(_02324_),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 split27 (.A(_02873_),
    .X(net111));
 sky130_fd_sc_hd__buf_4 split3 (.A(_01110_),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 split30 (.A(_02414_),
    .X(net114));
 sky130_fd_sc_hd__buf_4 split31 (.A(_05822_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 split5 (.A(_05985_),
    .X(net89));
 sky130_fd_sc_hd__buf_6 split6 (.A(_00569_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 split7 (.A(_05999_),
    .X(net91));
 sky130_fd_sc_hd__buf_6 split8 (.A(_00592_),
    .X(net120));
 sky130_fd_sc_hd__buf_2 split9 (.A(_04204_),
    .X(net121));
 assign out[31] = net82;
endmodule

