// This is the unpowered netlist.
module fp_mul (act,
    clk,
    done,
    inexact,
    inv,
    ov,
    rst,
    un,
    in1,
    in2,
    out,
    round_m);
 input act;
 input clk;
 output done;
 output inexact;
 output inv;
 output ov;
 input rst;
 output un;
 input [31:0] in1;
 input [31:0] in2;
 output [31:0] out;
 input [2:0] round_m;

 wire \M000[0] ;
 wire \M000[10] ;
 wire \M000[11] ;
 wire \M000[12] ;
 wire \M000[13] ;
 wire \M000[14] ;
 wire \M000[15] ;
 wire \M000[16] ;
 wire \M000[17] ;
 wire \M000[18] ;
 wire \M000[19] ;
 wire \M000[1] ;
 wire \M000[20] ;
 wire \M000[21] ;
 wire \M000[22] ;
 wire \M000[23] ;
 wire \M000[24] ;
 wire \M000[25] ;
 wire \M000[26] ;
 wire \M000[27] ;
 wire \M000[28] ;
 wire \M000[29] ;
 wire \M000[2] ;
 wire \M000[30] ;
 wire \M000[31] ;
 wire \M000[32] ;
 wire \M000[33] ;
 wire \M000[34] ;
 wire \M000[35] ;
 wire \M000[36] ;
 wire \M000[37] ;
 wire \M000[38] ;
 wire \M000[39] ;
 wire \M000[3] ;
 wire \M000[40] ;
 wire \M000[41] ;
 wire \M000[42] ;
 wire \M000[43] ;
 wire \M000[44] ;
 wire \M000[45] ;
 wire \M000[46] ;
 wire \M000[47] ;
 wire \M000[4] ;
 wire \M000[5] ;
 wire \M000[6] ;
 wire \M000[7] ;
 wire \M000[8] ;
 wire \M000[9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire done0_reg;
 wire forward;
 wire forward_c;
 wire inv_f;
 wire inv_f_c;
 wire \m1.out[0] ;
 wire \m1.out[10] ;
 wire \m1.out[11] ;
 wire \m1.out[12] ;
 wire \m1.out[13] ;
 wire \m1.out[14] ;
 wire \m1.out[15] ;
 wire \m1.out[16] ;
 wire \m1.out[17] ;
 wire \m1.out[18] ;
 wire \m1.out[19] ;
 wire \m1.out[1] ;
 wire \m1.out[20] ;
 wire \m1.out[21] ;
 wire \m1.out[22] ;
 wire \m1.out[23] ;
 wire \m1.out[24] ;
 wire \m1.out[25] ;
 wire \m1.out[26] ;
 wire \m1.out[27] ;
 wire \m1.out[28] ;
 wire \m1.out[29] ;
 wire \m1.out[2] ;
 wire \m1.out[30] ;
 wire \m1.out[31] ;
 wire \m1.out[32] ;
 wire \m1.out[33] ;
 wire \m1.out[34] ;
 wire \m1.out[35] ;
 wire \m1.out[36] ;
 wire \m1.out[37] ;
 wire \m1.out[38] ;
 wire \m1.out[39] ;
 wire \m1.out[3] ;
 wire \m1.out[40] ;
 wire \m1.out[41] ;
 wire \m1.out[42] ;
 wire \m1.out[43] ;
 wire \m1.out[44] ;
 wire \m1.out[45] ;
 wire \m1.out[46] ;
 wire \m1.out[47] ;
 wire \m1.out[4] ;
 wire \m1.out[5] ;
 wire \m1.out[6] ;
 wire \m1.out[7] ;
 wire \m1.out[8] ;
 wire \m1.out[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \out_f[23] ;
 wire \out_f[31] ;
 wire \out_f_c[23] ;
 wire \out_f_c[31] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA__06475__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__C (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__A2 (.DIODE(_01292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__B1 (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__C (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__S (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__C (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__A1 (.DIODE(\M000[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__B1 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__B1 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__S (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A3 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__A (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__B (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__B (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__B (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06797__B (.DIODE(_04803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06798__A (.DIODE(_04803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__A (.DIODE(_04519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__A (.DIODE(_04650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__A (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__B (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__A1 (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06823__S (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__A (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__A (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__B (.DIODE(_05437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06857__A (.DIODE(_05437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__B1 (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__B (.DIODE(_05306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__B (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__B (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__A1 (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__B (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__B1 (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__B (.DIODE(_06146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__S (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__B (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__B1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__A (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__A (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__B (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__C (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__D (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A (.DIODE(_06185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__A (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__B (.DIODE(_06189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__C (.DIODE(_06190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__A (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__B (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__C (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__D (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__A (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__A (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__A (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__A (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__C (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__D (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__A (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__A (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__C (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__D (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__A (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__A (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__B (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__C (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__D (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__B (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__C (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__D (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__A (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__B (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A (.DIODE(_06249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__B (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A_N (.DIODE(_06244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07047__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__B (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__C (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__D (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07056__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__B (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__C (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__D (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__A (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__B (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__C (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__D (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__B (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__C (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__D (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__C (.DIODE(_06294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A1 (.DIODE(_06180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A4 (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__A (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__C_N (.DIODE(_06249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07084__D (.DIODE(_06244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__D (.DIODE(_06294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__A (.DIODE(_06190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__B (.DIODE(_06180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__B (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__D (.DIODE(_06294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A (.DIODE(_06180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__D (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A (.DIODE(_06180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__D (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__A (.DIODE(_06317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__A (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__A (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__B (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__A (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__B (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__D (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A1 (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A2 (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B1 (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B2 (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__B (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__A (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__B (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__C (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__D (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A1 (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__A2 (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__B1 (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__B2 (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__B (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__C (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__D (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A1 (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A2 (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B1 (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B2 (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__A (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__B (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__C (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__D (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A1 (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A2 (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B1 (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B2 (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__B (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__B (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A2 (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__B (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__B (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A2 (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__B (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A1 (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A2 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__B (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A1 (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A2 (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__B (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__C (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__B (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A (.DIODE(_00069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A1 (.DIODE(_00069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__B (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07515__A (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A (.DIODE(_00069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A1 (.DIODE(_00069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__B (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A1 (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A2 (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__B1 (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__B2 (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__A (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__B (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__B (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__B (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__B (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__B (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07783__B (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__B (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__B (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__B (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A1 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__B (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__B (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__B (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__B (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__B (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__A (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08161__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08161__B (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__B (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08269__A (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08269__B (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A (.DIODE(_06268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A (.DIODE(_06275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A (.DIODE(_06260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__A (.DIODE(_06272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__B (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__B (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__B (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__C (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__D (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A1 (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A2 (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__B1 (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__B2 (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B (.DIODE(_01268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A (.DIODE(_01268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__B (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__B (.DIODE(_01294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A (.DIODE(_01294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__B (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08506__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__C (.DIODE(_01294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__B (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__B (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A (.DIODE(_01346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08552__C (.DIODE(_01346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08557__A (.DIODE(_01354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A (.DIODE(_01354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__B (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B (.DIODE(_01396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A (.DIODE(_01396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__B (.DIODE(_01396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__B (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__B (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__C (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08618__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A1 (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A2 (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A (.DIODE(_01294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__B (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08674__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__A (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08684__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__A (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__A (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__B (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__C (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__A (.DIODE(_01543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A (.DIODE(_01543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__B (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08754__B (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__A (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__B (.DIODE(_01354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08776__A (.DIODE(_01354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__A (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08790__B (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__B (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A1 (.DIODE(_01268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__B (.DIODE(_01543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A (.DIODE(_01543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__A (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__B (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__B (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__A (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__B (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__A2 (.DIODE(_01531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__B (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09016__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__B (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__C (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__D (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A1 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A2 (.DIODE(_06209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__B1 (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__B2 (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09024__B (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A (.DIODE(_01580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09075__A (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__B (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09079__B (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09097__B (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09107__C (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__A (.DIODE(_01955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__A (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__B (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__B (.DIODE(_06229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09208__B (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09210__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B (.DIODE(_06210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__A1 (.DIODE(_01268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__B (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__B (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__B (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__B (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09379__C (.DIODE(_02250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__B (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__B (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__B (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09412__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09440__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09442__B (.DIODE(_06201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__B (.DIODE(_06213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__B (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__C (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__B (.DIODE(_06204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__B (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__A (.DIODE(_06270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__B (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__B (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__B (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09576__B (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__C (.DIODE(_02490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__B (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__B (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__B (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__B (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09636__B (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__B (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09692__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__B (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__B (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__B (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__C (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__D (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A2 (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B2 (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A (.DIODE(_06327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__B (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09788__B (.DIODE(_06329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__A (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__B (.DIODE(_06271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__C (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__B (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__B (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__B (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__A (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__C (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__A (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__B (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__B (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__B (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__C (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A1 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A2 (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__B (.DIODE(_06208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B (.DIODE(_06195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A1 (.DIODE(_01268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__B (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A (.DIODE(_06269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__B (.DIODE(_06276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__C (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10063__B (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10065__B (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__A (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__B (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__B (.DIODE(_03054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__C (.DIODE(_03054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10178__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__B (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__B (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__A (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__B (.DIODE(_06205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__C (.DIODE(_06214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A2 (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__B1 (.DIODE(_06206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__A (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__B (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__A (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__A (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__C (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__B (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__A (.DIODE(_00299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__B (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__B (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10368__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10368__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__B (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__B (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__C (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__B (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__B (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__A (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__B (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__C (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__A2 (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B (.DIODE(_06211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__B (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__C (.DIODE(_06215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__B (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__B (.DIODE(_06262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__C (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__B (.DIODE(_06227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__A (.DIODE(_03371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__B (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__B (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A1 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__A2 (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__B (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__B (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__A (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10752__A (.DIODE(_06259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10752__B (.DIODE(_06261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10752__C (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10753__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A (.DIODE(_06263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__B (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10794__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__B (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__B (.DIODE(_06219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__B (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__B (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__C (.DIODE(_00176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__A (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__A1 (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__A2 (.DIODE(_06196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__B1 (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__A2 (.DIODE(_06212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__A (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__B (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10976__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__A (.DIODE(_00175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__B (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__C (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__B (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__A (.DIODE(_06289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__B (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__B (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__B (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__A (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__B (.DIODE(_00921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__B (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__B (.DIODE(_00780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__A (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__B (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__A (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11114__A (.DIODE(_06387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__A (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A1 (.DIODE(_04200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A2 (.DIODE(_02969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__B1_N (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A (.DIODE(_04209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__B (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__B (.DIODE(_00069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__B (.DIODE(_06266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__C (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__A (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A (.DIODE(_00439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__B (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A (.DIODE(_06286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__B (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__B (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__B (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__B (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__B (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__A (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__B (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__B (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__B (.DIODE(_06220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A_N (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__B (.DIODE(_04294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__B (.DIODE(_06199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__C (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A (.DIODE(_00270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A1 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__B (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__C (.DIODE(_06202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11324__A_N (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__C (.DIODE(_04340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__A2 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__A1 (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__A2 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__B1 (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A (.DIODE(_06264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__B (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__C (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__B (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__B (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__A (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__A (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__B (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__A (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11436__B (.DIODE(_06230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__B (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__C (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11438__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__A (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A1 (.DIODE(_04495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__B (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__B (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__A (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__B (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__C (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A1 (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A2 (.DIODE(_06226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__B1 (.DIODE(_06200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A1 (.DIODE(_04206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__B (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__B (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A (.DIODE(_00561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__B (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__A1 (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__A2 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__B1 (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B (.DIODE(_06290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__C (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__A (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__B (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__B (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__A (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__B (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11634__A (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11634__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__B (.DIODE(_00926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__B (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__A (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__B (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__B (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__C (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__A (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A1 (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__A (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__C (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11701__B (.DIODE(_04783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__A (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11711__B (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__A (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__B (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__C (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__D (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__A1 (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__A2 (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__B1 (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__B2 (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__B (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A2 (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B1 (.DIODE(_06288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__B (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__C (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__D (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A1 (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A2 (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B1 (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__B2 (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__A (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__A (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__B (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__B (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__C (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__D (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__A1 (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__A2 (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__B1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__B2 (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__A (.DIODE(_04740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__A_N (.DIODE(_04790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__B (.DIODE(_04790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__C (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__B (.DIODE(_04926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__A_N (.DIODE(_04926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__B (.DIODE(_04783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__A (.DIODE(_04783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A1 (.DIODE(_04204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A (.DIODE(_04200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__B (.DIODE(_04945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__B (.DIODE(_01268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__B (.DIODE(_04950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A (.DIODE(_04950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__B (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A2 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__B1 (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__A (.DIODE(_06282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11878__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__A (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__B (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__C (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__D (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__A1 (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__A2 (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__B1 (.DIODE(_06284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__B2 (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11893__A (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11893__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__B (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__B (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__A (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__B (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__A (.DIODE(_04495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__A1 (.DIODE(_04495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__A (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__C_N (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A2 (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__B1 (.DIODE(_06231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A2 (.DIODE(_06225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__A1 (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__B (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A1 (.DIODE(_06280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A2 (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__B1 (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__B (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__C (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__D (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A1 (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A2 (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__B1 (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__B2 (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__B (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__B (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__C (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__D (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__B (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__B (.DIODE(_06228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__A1 (.DIODE(_04950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__A (.DIODE(_06278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__B (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__A1 (.DIODE(_00701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__A2 (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__B1 (.DIODE(_00849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__B (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__B (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A1 (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__B (.DIODE(_00918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__B (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__B (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__A (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__B (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__C (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__D (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__B (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__C (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__D (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__A1 (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__A2 (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__B1 (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__B2 (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__A (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__B (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__B (.DIODE(_06177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__B (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__A (.DIODE(_06283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A1 (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A2 (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__B1 (.DIODE(_06279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A2 (.DIODE(_06236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A3 (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__C (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__D (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__A1 (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__A2 (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B2 (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__A (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__B (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__C (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__D (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__C_N (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A2 (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__B1 (.DIODE(_06218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A2 (.DIODE(_06221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__A (.DIODE(_04950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A1 (.DIODE(_01831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A2 (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__B1 (.DIODE(_01158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A (.DIODE(_01211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__B (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__A (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12346__B (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__A (.DIODE(_06242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12348__B (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12362__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__C (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__D (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__B2 (.DIODE(_01280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__A (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12425__B (.DIODE(_02180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A (.DIODE(_01422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__A1 (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__B1 (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__A (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__B (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__B (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__C (.DIODE(_06175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__D (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A1 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A2 (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__B1 (.DIODE(_06243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__B2 (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__A2 (.DIODE(_06240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__A3 (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__C (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__D (.DIODE(_06173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A1 (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A2 (.DIODE(_06171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__B1 (.DIODE(_06298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__B2 (.DIODE(_01278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__A (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__B (.DIODE(_06222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__B (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__A_N (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__A (.DIODE(_06237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__B (.DIODE(_06185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__B (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__C (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__D (.DIODE(_06187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__A1 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__A2 (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__B1 (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__B2 (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__B (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__C (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A2 (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__B1 (.DIODE(_06174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__A (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__B (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__A (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__C (.DIODE(_05748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__A1 (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__A2 (.DIODE(_01692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__B1 (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__B2 (.DIODE(_01921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A (.DIODE(_06234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__A (.DIODE(_04495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12595__B (.DIODE(_06185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A1 (.DIODE(_04495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A (.DIODE(_06172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12647__A (.DIODE(_04950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__A (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__B (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__C (.DIODE(_05748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A1 (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A2 (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__B1 (.DIODE(_03905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__B2 (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__A (.DIODE(_06239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__12671__A (.DIODE(_06241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__B (.DIODE(_06185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__A (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__B (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__C (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A1 (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A2 (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__B1 (.DIODE(_06176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__A (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__B (.DIODE(_06183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A1 (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A1 (.DIODE(_04853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12767__B (.DIODE(_02423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A (.DIODE(_06248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12769__A (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A1 (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A1 (.DIODE(_04495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A (.DIODE(_06299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__B (.DIODE(_06184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__B (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__B (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A2 (.DIODE(_01922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A (.DIODE(_06250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A2 (.DIODE(_06247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A3 (.DIODE(_02181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A2 (.DIODE(_01446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12900__A2 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12901__A1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A2 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__A2 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A1 (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12907__A2 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12908__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A (.DIODE(_01336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12919__A (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12921__A (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__S (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__S (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__A (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12951__S (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A (.DIODE(_04378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__S (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__B1 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__S (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12966__B1 (.DIODE(_03072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12967__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12970__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__RESET_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12972__RESET_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__RESET_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__RESET_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__RESET_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__RESET_B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13001__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__RESET_B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__RESET_B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13030__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__CLK (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__D (.DIODE(\m1.out[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__D (.DIODE(\m1.out[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13033__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__D (.DIODE(\m1.out[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13034__RESET_B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__D (.DIODE(\m1.out[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13037__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13039__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13040__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__CLK (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13050__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__RESET_B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__13052__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13052__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__CLK (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__D (.DIODE(inv_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__D (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__CLK (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold160_A (.DIODE(\M000[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold39_A (.DIODE(_01292_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_998 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_900 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_814 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1010 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06458_ (.A(net164),
    .Y(_01117_));
 sky130_fd_sc_hd__buf_2 _06459_ (.A(net165),
    .X(_01128_));
 sky130_fd_sc_hd__inv_2 _06460_ (.A(net182),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _06461_ (.A(_01128_),
    .B(net183),
    .Y(_01150_));
 sky130_fd_sc_hd__o21ai_1 _06462_ (.A1(net231),
    .A2(_01128_),
    .B1(net184),
    .Y(_01161_));
 sky130_fd_sc_hd__inv_2 _06463_ (.A(net138),
    .Y(_01172_));
 sky130_fd_sc_hd__nand2_1 _06464_ (.A(net139),
    .B(net164),
    .Y(_01183_));
 sky130_fd_sc_hd__o21ai_1 _06465_ (.A1(net164),
    .A2(net179),
    .B1(net140),
    .Y(_01194_));
 sky130_fd_sc_hd__inv_2 _06466_ (.A(net141),
    .Y(_01205_));
 sky130_fd_sc_hd__or4_1 _06467_ (.A(\M000[17] ),
    .B(\M000[16] ),
    .C(\M000[19] ),
    .D(\M000[18] ),
    .X(_01216_));
 sky130_fd_sc_hd__or3_1 _06468_ (.A(net155),
    .B(\M000[20] ),
    .C(_01216_),
    .X(_01227_));
 sky130_fd_sc_hd__or4_1 _06469_ (.A(\M000[9] ),
    .B(\M000[8] ),
    .C(\M000[11] ),
    .D(\M000[10] ),
    .X(_01238_));
 sky130_fd_sc_hd__or4_1 _06470_ (.A(\M000[1] ),
    .B(\M000[0] ),
    .C(\M000[3] ),
    .D(\M000[2] ),
    .X(_01249_));
 sky130_fd_sc_hd__or4_1 _06471_ (.A(\M000[5] ),
    .B(\M000[4] ),
    .C(\M000[7] ),
    .D(\M000[6] ),
    .X(_01260_));
 sky130_fd_sc_hd__or4_1 _06472_ (.A(\M000[13] ),
    .B(\M000[12] ),
    .C(\M000[15] ),
    .D(\M000[14] ),
    .X(_01271_));
 sky130_fd_sc_hd__or4_2 _06473_ (.A(_01238_),
    .B(_01249_),
    .C(_01260_),
    .D(_01271_),
    .X(_01281_));
 sky130_fd_sc_hd__or2_4 _06474_ (.A(net156),
    .B(_01281_),
    .X(_01292_));
 sky130_fd_sc_hd__inv_2 _06475_ (.A(net67),
    .Y(_01303_));
 sky130_fd_sc_hd__inv_2 _06476_ (.A(net66),
    .Y(_01314_));
 sky130_fd_sc_hd__and3_1 _06477_ (.A(_01303_),
    .B(_01314_),
    .C(net65),
    .X(_01325_));
 sky130_fd_sc_hd__clkbuf_4 _06478_ (.A(_01325_),
    .X(_01336_));
 sky130_fd_sc_hd__clkbuf_4 _06479_ (.A(net164),
    .X(_01347_));
 sky130_fd_sc_hd__clkbuf_4 _06480_ (.A(_01347_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _06481_ (.A0(net132),
    .A1(net179),
    .S(_01358_),
    .X(_01369_));
 sky130_fd_sc_hd__o211a_1 _06482_ (.A1(net142),
    .A2(_01292_),
    .B1(_01336_),
    .C1(net133),
    .X(_01380_));
 sky130_fd_sc_hd__inv_2 _06483_ (.A(net143),
    .Y(_01391_));
 sky130_fd_sc_hd__nor2_1 _06484_ (.A(net133),
    .B(net157),
    .Y(_01402_));
 sky130_fd_sc_hd__and3_1 _06485_ (.A(_01303_),
    .B(net66),
    .C(net65),
    .X(_01413_));
 sky130_fd_sc_hd__inv_2 _06486_ (.A(net65),
    .Y(_01424_));
 sky130_fd_sc_hd__and3_1 _06487_ (.A(_01303_),
    .B(_01424_),
    .C(net66),
    .X(_01435_));
 sky130_fd_sc_hd__xnor2_4 _06488_ (.A(net25),
    .B(net57),
    .Y(_01446_));
 sky130_fd_sc_hd__mux2_1 _06489_ (.A0(_01413_),
    .A1(_01435_),
    .S(_01446_),
    .X(_01457_));
 sky130_fd_sc_hd__clkbuf_4 _06490_ (.A(_01457_),
    .X(_01468_));
 sky130_fd_sc_hd__nand2_2 _06491_ (.A(net158),
    .B(_01468_),
    .Y(_01478_));
 sky130_fd_sc_hd__and3_1 _06492_ (.A(_01314_),
    .B(_01424_),
    .C(net67),
    .X(_01489_));
 sky130_fd_sc_hd__inv_2 _06493_ (.A(_01489_),
    .Y(_01500_));
 sky130_fd_sc_hd__inv_2 _06494_ (.A(net133),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_4 _06495_ (.A(_01500_),
    .B(_01511_),
    .Y(_01522_));
 sky130_fd_sc_hd__nor2_2 _06496_ (.A(_01522_),
    .B(_01468_),
    .Y(_01533_));
 sky130_fd_sc_hd__inv_2 _06497_ (.A(_01533_),
    .Y(_01544_));
 sky130_fd_sc_hd__nand2_2 _06498_ (.A(_01478_),
    .B(_01544_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _06499_ (.A(net144),
    .B(_01555_),
    .Y(_01566_));
 sky130_fd_sc_hd__inv_2 _06500_ (.A(net145),
    .Y(_01577_));
 sky130_fd_sc_hd__buf_1 _06501_ (.A(net129),
    .X(_01588_));
 sky130_fd_sc_hd__inv_2 _06502_ (.A(net189),
    .Y(_01599_));
 sky130_fd_sc_hd__nand2_1 _06503_ (.A(_01128_),
    .B(net190),
    .Y(_01610_));
 sky130_fd_sc_hd__o21ai_1 _06504_ (.A1(net272),
    .A2(_01128_),
    .B1(net191),
    .Y(_01621_));
 sky130_fd_sc_hd__inv_2 _06505_ (.A(net202),
    .Y(_01632_));
 sky130_fd_sc_hd__mux2_1 _06506_ (.A0(net203),
    .A1(net190),
    .S(net164),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _06507_ (.A0(net139),
    .A1(net203),
    .S(net164),
    .X(_01654_));
 sky130_fd_sc_hd__or2_1 _06508_ (.A(net141),
    .B(net204),
    .X(_01665_));
 sky130_fd_sc_hd__or2_1 _06509_ (.A(_01643_),
    .B(_01665_),
    .X(_01676_));
 sky130_fd_sc_hd__nor2_1 _06510_ (.A(net192),
    .B(_01676_),
    .Y(_01686_));
 sky130_fd_sc_hd__or2_1 _06511_ (.A(net263),
    .B(net165),
    .X(_01697_));
 sky130_fd_sc_hd__o21a_1 _06512_ (.A1(_01347_),
    .A2(net283),
    .B1(_01697_),
    .X(_01708_));
 sky130_fd_sc_hd__inv_2 _06513_ (.A(net284),
    .Y(_01719_));
 sky130_fd_sc_hd__mux2_1 _06514_ (.A0(net272),
    .A1(net283),
    .S(_01347_),
    .X(_01730_));
 sky130_fd_sc_hd__inv_2 _06515_ (.A(net273),
    .Y(_01741_));
 sky130_fd_sc_hd__nor2_1 _06516_ (.A(_01719_),
    .B(_01741_),
    .Y(_01752_));
 sky130_fd_sc_hd__mux2_1 _06517_ (.A0(net237),
    .A1(\M000[31] ),
    .S(_01347_),
    .X(_01763_));
 sky130_fd_sc_hd__inv_2 _06518_ (.A(net238),
    .Y(_01774_));
 sky130_fd_sc_hd__mux2_1 _06519_ (.A0(net263),
    .A1(net237),
    .S(_01347_),
    .X(_01785_));
 sky130_fd_sc_hd__inv_2 _06520_ (.A(net264),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _06521_ (.A(net239),
    .B(_01796_),
    .Y(_01807_));
 sky130_fd_sc_hd__and3_1 _06522_ (.A(_01686_),
    .B(_01752_),
    .C(_01807_),
    .X(_01818_));
 sky130_fd_sc_hd__inv_2 _06523_ (.A(net278),
    .Y(_01829_));
 sky130_fd_sc_hd__mux2_2 _06524_ (.A0(net279),
    .A1(net183),
    .S(_01347_),
    .X(_01840_));
 sky130_fd_sc_hd__inv_2 _06525_ (.A(_01840_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _06526_ (.A(_01818_),
    .B(_01851_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_1 _06527_ (.A(_01862_),
    .B(net185),
    .Y(_01873_));
 sky130_fd_sc_hd__or2_1 _06528_ (.A(net185),
    .B(_01862_),
    .X(_01884_));
 sky130_fd_sc_hd__a21oi_1 _06529_ (.A1(_01873_),
    .A2(_01884_),
    .B1(net146),
    .Y(_01895_));
 sky130_fd_sc_hd__a211oi_1 _06530_ (.A1(net185),
    .A2(net146),
    .B1(net130),
    .C1(_01895_),
    .Y(_00033_));
 sky130_fd_sc_hd__mux2_1 _06531_ (.A0(net231),
    .A1(net225),
    .S(_01347_),
    .X(_01915_));
 sky130_fd_sc_hd__inv_2 _06532_ (.A(net232),
    .Y(_01926_));
 sky130_fd_sc_hd__nor2_1 _06533_ (.A(net185),
    .B(_01840_),
    .Y(_01937_));
 sky130_fd_sc_hd__nand2_1 _06534_ (.A(_01818_),
    .B(_01937_),
    .Y(_01948_));
 sky130_fd_sc_hd__or2_1 _06535_ (.A(_01926_),
    .B(_01948_),
    .X(_01959_));
 sky130_fd_sc_hd__nand2_1 _06536_ (.A(_01948_),
    .B(_01926_),
    .Y(_01970_));
 sky130_fd_sc_hd__nand2_1 _06537_ (.A(_01959_),
    .B(_01970_),
    .Y(_01981_));
 sky130_fd_sc_hd__buf_2 _06538_ (.A(_01522_),
    .X(_01992_));
 sky130_fd_sc_hd__and2_1 _06539_ (.A(_01981_),
    .B(_01992_),
    .X(_02003_));
 sky130_fd_sc_hd__inv_2 _06540_ (.A(_01468_),
    .Y(_02014_));
 sky130_fd_sc_hd__nor2_2 _06541_ (.A(_02014_),
    .B(net158),
    .Y(_02025_));
 sky130_fd_sc_hd__buf_2 _06542_ (.A(_02025_),
    .X(_02036_));
 sky130_fd_sc_hd__and2_1 _06543_ (.A(_02036_),
    .B(_01981_),
    .X(_02047_));
 sky130_fd_sc_hd__buf_2 _06544_ (.A(_01478_),
    .X(_02058_));
 sky130_fd_sc_hd__clkbuf_4 _06545_ (.A(_01544_),
    .X(_02069_));
 sky130_fd_sc_hd__a21oi_1 _06546_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net232),
    .Y(_02080_));
 sky130_fd_sc_hd__or3_1 _06547_ (.A(_02003_),
    .B(_02047_),
    .C(_02080_),
    .X(_02091_));
 sky130_fd_sc_hd__inv_2 _06548_ (.A(_01336_),
    .Y(_02102_));
 sky130_fd_sc_hd__clkbuf_4 _06549_ (.A(_02102_),
    .X(_02113_));
 sky130_fd_sc_hd__clkbuf_4 _06550_ (.A(_02113_),
    .X(_02124_));
 sky130_fd_sc_hd__clkbuf_4 _06551_ (.A(net188),
    .X(_02135_));
 sky130_fd_sc_hd__clkbuf_4 _06552_ (.A(_02113_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_4 _06553_ (.A(net133),
    .X(_02157_));
 sky130_fd_sc_hd__clkbuf_4 _06554_ (.A(_02157_),
    .X(_02167_));
 sky130_fd_sc_hd__buf_2 _06555_ (.A(_02157_),
    .X(_02178_));
 sky130_fd_sc_hd__nor2_1 _06556_ (.A(_02178_),
    .B(net232),
    .Y(_02189_));
 sky130_fd_sc_hd__a21oi_1 _06557_ (.A1(_01981_),
    .A2(_02167_),
    .B1(_02189_),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_1 _06558_ (.A(_02146_),
    .B(net233),
    .Y(_02211_));
 sky130_fd_sc_hd__a211o_1 _06559_ (.A1(_02091_),
    .A2(_02124_),
    .B1(_02135_),
    .C1(net234),
    .X(_02222_));
 sky130_fd_sc_hd__inv_2 _06560_ (.A(net235),
    .Y(_00003_));
 sky130_fd_sc_hd__or2_1 _06561_ (.A(net258),
    .B(net165),
    .X(_02243_));
 sky130_fd_sc_hd__o21a_1 _06562_ (.A1(_01358_),
    .A2(net225),
    .B1(_02243_),
    .X(_02254_));
 sky130_fd_sc_hd__a21oi_1 _06563_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net226),
    .Y(_02265_));
 sky130_fd_sc_hd__inv_2 _06564_ (.A(net226),
    .Y(_02276_));
 sky130_fd_sc_hd__and2_1 _06565_ (.A(_01959_),
    .B(_02276_),
    .X(_02287_));
 sky130_fd_sc_hd__nand2_1 _06566_ (.A(_01686_),
    .B(_01752_),
    .Y(_02298_));
 sky130_fd_sc_hd__or2_1 _06567_ (.A(_01796_),
    .B(_02298_),
    .X(_02309_));
 sky130_fd_sc_hd__or2_1 _06568_ (.A(net239),
    .B(_02309_),
    .X(_02320_));
 sky130_fd_sc_hd__or2_1 _06569_ (.A(_01840_),
    .B(_02320_),
    .X(_02331_));
 sky130_fd_sc_hd__or3_1 _06570_ (.A(net185),
    .B(_01926_),
    .C(net280),
    .X(_02342_));
 sky130_fd_sc_hd__nor2_1 _06571_ (.A(_02276_),
    .B(_02342_),
    .Y(_02353_));
 sky130_fd_sc_hd__or2_1 _06572_ (.A(_02287_),
    .B(_02353_),
    .X(_02364_));
 sky130_fd_sc_hd__and2_1 _06573_ (.A(_02364_),
    .B(_01992_),
    .X(_02375_));
 sky130_fd_sc_hd__and2_1 _06574_ (.A(_02364_),
    .B(_02036_),
    .X(_02386_));
 sky130_fd_sc_hd__or3_1 _06575_ (.A(_02265_),
    .B(_02375_),
    .C(_02386_),
    .X(_02397_));
 sky130_fd_sc_hd__nor2_1 _06576_ (.A(net226),
    .B(_02178_),
    .Y(_02408_));
 sky130_fd_sc_hd__a21oi_1 _06577_ (.A1(_02364_),
    .A2(_02167_),
    .B1(net227),
    .Y(_02418_));
 sky130_fd_sc_hd__nor2_1 _06578_ (.A(_02146_),
    .B(net228),
    .Y(_02429_));
 sky130_fd_sc_hd__a211o_1 _06579_ (.A1(_02397_),
    .A2(_02124_),
    .B1(_02135_),
    .C1(net229),
    .X(_02440_));
 sky130_fd_sc_hd__inv_2 _06580_ (.A(net230),
    .Y(_00004_));
 sky130_fd_sc_hd__mux2_1 _06581_ (.A0(net258),
    .A1(net207),
    .S(_01347_),
    .X(_02461_));
 sky130_fd_sc_hd__inv_2 _06582_ (.A(net259),
    .Y(_02472_));
 sky130_fd_sc_hd__and3_1 _06583_ (.A(_01937_),
    .B(net232),
    .C(net226),
    .X(_02483_));
 sky130_fd_sc_hd__nand2_1 _06584_ (.A(_01818_),
    .B(_02483_),
    .Y(_02494_));
 sky130_fd_sc_hd__or2_1 _06585_ (.A(_02472_),
    .B(_02494_),
    .X(_02505_));
 sky130_fd_sc_hd__nand2_1 _06586_ (.A(_02494_),
    .B(_02472_),
    .Y(_02516_));
 sky130_fd_sc_hd__nand2_1 _06587_ (.A(_02505_),
    .B(_02516_),
    .Y(_02527_));
 sky130_fd_sc_hd__and2_1 _06588_ (.A(_02527_),
    .B(_01522_),
    .X(_02538_));
 sky130_fd_sc_hd__and2_1 _06589_ (.A(_02025_),
    .B(_02527_),
    .X(_02549_));
 sky130_fd_sc_hd__a21oi_1 _06590_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net259),
    .Y(_02560_));
 sky130_fd_sc_hd__or3_1 _06591_ (.A(_02538_),
    .B(_02549_),
    .C(_02560_),
    .X(_02571_));
 sky130_fd_sc_hd__nor2_1 _06592_ (.A(_02178_),
    .B(net259),
    .Y(_02582_));
 sky130_fd_sc_hd__a21oi_1 _06593_ (.A1(_02527_),
    .A2(_02167_),
    .B1(_02582_),
    .Y(_02593_));
 sky130_fd_sc_hd__nor2_1 _06594_ (.A(_02146_),
    .B(net260),
    .Y(_02604_));
 sky130_fd_sc_hd__a211o_1 _06595_ (.A1(_02571_),
    .A2(_02124_),
    .B1(_02135_),
    .C1(net261),
    .X(_02615_));
 sky130_fd_sc_hd__inv_2 _06596_ (.A(net262),
    .Y(_00005_));
 sky130_fd_sc_hd__or2_1 _06597_ (.A(net248),
    .B(net165),
    .X(_02636_));
 sky130_fd_sc_hd__o21a_1 _06598_ (.A1(_01347_),
    .A2(net207),
    .B1(_02636_),
    .X(_02647_));
 sky130_fd_sc_hd__a21oi_1 _06599_ (.A1(_01478_),
    .A2(_02069_),
    .B1(net208),
    .Y(_02658_));
 sky130_fd_sc_hd__inv_2 _06600_ (.A(net208),
    .Y(_02669_));
 sky130_fd_sc_hd__and2_1 _06601_ (.A(_02505_),
    .B(_02669_),
    .X(_02680_));
 sky130_fd_sc_hd__nand2_1 _06602_ (.A(_02353_),
    .B(net259),
    .Y(_02690_));
 sky130_fd_sc_hd__nor2_1 _06603_ (.A(_02669_),
    .B(_02690_),
    .Y(_02701_));
 sky130_fd_sc_hd__or2_1 _06604_ (.A(_02680_),
    .B(_02701_),
    .X(_02712_));
 sky130_fd_sc_hd__and2_1 _06605_ (.A(_02712_),
    .B(_01992_),
    .X(_02723_));
 sky130_fd_sc_hd__and2_1 _06606_ (.A(_02712_),
    .B(_02036_),
    .X(_02734_));
 sky130_fd_sc_hd__or3_1 _06607_ (.A(_02658_),
    .B(_02723_),
    .C(_02734_),
    .X(_02745_));
 sky130_fd_sc_hd__nor2_1 _06608_ (.A(net208),
    .B(_02178_),
    .Y(_02756_));
 sky130_fd_sc_hd__a21oi_1 _06609_ (.A1(_02712_),
    .A2(_02167_),
    .B1(net209),
    .Y(_02767_));
 sky130_fd_sc_hd__nor2_1 _06610_ (.A(_02146_),
    .B(net210),
    .Y(_02778_));
 sky130_fd_sc_hd__a211o_1 _06611_ (.A1(_02745_),
    .A2(_02124_),
    .B1(_02135_),
    .C1(net211),
    .X(_02789_));
 sky130_fd_sc_hd__inv_2 _06612_ (.A(net212),
    .Y(_00006_));
 sky130_fd_sc_hd__mux2_1 _06613_ (.A0(net248),
    .A1(net268),
    .S(_01358_),
    .X(_02810_));
 sky130_fd_sc_hd__a21oi_1 _06614_ (.A1(_01478_),
    .A2(_02069_),
    .B1(net249),
    .Y(_02821_));
 sky130_fd_sc_hd__inv_2 _06615_ (.A(net249),
    .Y(_02832_));
 sky130_fd_sc_hd__or3_1 _06616_ (.A(_02472_),
    .B(_02669_),
    .C(_02494_),
    .X(_02843_));
 sky130_fd_sc_hd__or2_1 _06617_ (.A(_02832_),
    .B(_02843_),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _06618_ (.A(_02843_),
    .B(_02832_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _06619_ (.A(_02854_),
    .B(_02865_),
    .Y(_02876_));
 sky130_fd_sc_hd__and2_1 _06620_ (.A(_02876_),
    .B(_01992_),
    .X(_02887_));
 sky130_fd_sc_hd__and2_1 _06621_ (.A(_02876_),
    .B(_02036_),
    .X(_02898_));
 sky130_fd_sc_hd__or3_1 _06622_ (.A(_02821_),
    .B(_02887_),
    .C(_02898_),
    .X(_02909_));
 sky130_fd_sc_hd__nor2_1 _06623_ (.A(_02157_),
    .B(net249),
    .Y(_02920_));
 sky130_fd_sc_hd__a21oi_1 _06624_ (.A1(_02876_),
    .A2(_02167_),
    .B1(net250),
    .Y(_02931_));
 sky130_fd_sc_hd__nor2_1 _06625_ (.A(_02146_),
    .B(net251),
    .Y(_02942_));
 sky130_fd_sc_hd__a211o_1 _06626_ (.A1(_02909_),
    .A2(_02124_),
    .B1(_02135_),
    .C1(net252),
    .X(_02953_));
 sky130_fd_sc_hd__inv_2 _06627_ (.A(net253),
    .Y(_00007_));
 sky130_fd_sc_hd__or2_1 _06628_ (.A(net255),
    .B(_01128_),
    .X(_02973_));
 sky130_fd_sc_hd__o21a_1 _06629_ (.A1(_01358_),
    .A2(net268),
    .B1(_02973_),
    .X(_02984_));
 sky130_fd_sc_hd__inv_2 _06630_ (.A(net269),
    .Y(_02995_));
 sky130_fd_sc_hd__and2_1 _06631_ (.A(_02854_),
    .B(_02995_),
    .X(_03006_));
 sky130_fd_sc_hd__nand2_1 _06632_ (.A(_02701_),
    .B(net249),
    .Y(_03017_));
 sky130_fd_sc_hd__nor2_1 _06633_ (.A(_02995_),
    .B(_03017_),
    .Y(_03028_));
 sky130_fd_sc_hd__or2_1 _06634_ (.A(_03006_),
    .B(_03028_),
    .X(_03039_));
 sky130_fd_sc_hd__nor2_1 _06635_ (.A(net269),
    .B(_02167_),
    .Y(_03050_));
 sky130_fd_sc_hd__a21oi_1 _06636_ (.A1(net281),
    .A2(_02167_),
    .B1(_03050_),
    .Y(_03061_));
 sky130_fd_sc_hd__inv_2 _06637_ (.A(net130),
    .Y(_03072_));
 sky130_fd_sc_hd__a21oi_1 _06638_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net269),
    .Y(_03083_));
 sky130_fd_sc_hd__and2_1 _06639_ (.A(net281),
    .B(_01992_),
    .X(_03094_));
 sky130_fd_sc_hd__and2_1 _06640_ (.A(net281),
    .B(_02036_),
    .X(_03105_));
 sky130_fd_sc_hd__o31ai_1 _06641_ (.A1(_03083_),
    .A2(_03094_),
    .A3(_03105_),
    .B1(_02124_),
    .Y(_03116_));
 sky130_fd_sc_hd__o211ai_1 _06642_ (.A1(_02124_),
    .A2(net282),
    .B1(_03072_),
    .C1(_03116_),
    .Y(_03127_));
 sky130_fd_sc_hd__inv_2 _06643_ (.A(_03127_),
    .Y(_00008_));
 sky130_fd_sc_hd__mux2_1 _06644_ (.A0(net255),
    .A1(net219),
    .S(_01347_),
    .X(_03148_));
 sky130_fd_sc_hd__nor2_1 _06645_ (.A(_02669_),
    .B(_02472_),
    .Y(_03159_));
 sky130_fd_sc_hd__and4_1 _06646_ (.A(_02483_),
    .B(net249),
    .C(_03159_),
    .D(net269),
    .X(_03170_));
 sky130_fd_sc_hd__and2_1 _06647_ (.A(_01818_),
    .B(net270),
    .X(_03181_));
 sky130_fd_sc_hd__or2_1 _06648_ (.A(net256),
    .B(net271),
    .X(_03192_));
 sky130_fd_sc_hd__nand2_1 _06649_ (.A(net271),
    .B(net256),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2_1 _06650_ (.A(_03192_),
    .B(_03203_),
    .Y(_03214_));
 sky130_fd_sc_hd__and2_1 _06651_ (.A(_03214_),
    .B(_01522_),
    .X(_03225_));
 sky130_fd_sc_hd__and2_1 _06652_ (.A(_02025_),
    .B(_03214_),
    .X(_03235_));
 sky130_fd_sc_hd__a21oi_1 _06653_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net256),
    .Y(_03246_));
 sky130_fd_sc_hd__or3_1 _06654_ (.A(_03225_),
    .B(_03235_),
    .C(_03246_),
    .X(_03257_));
 sky130_fd_sc_hd__nor2_1 _06655_ (.A(_02157_),
    .B(net256),
    .Y(_03268_));
 sky130_fd_sc_hd__a21oi_1 _06656_ (.A1(_03214_),
    .A2(_02167_),
    .B1(_03268_),
    .Y(_03279_));
 sky130_fd_sc_hd__nor2_1 _06657_ (.A(_02113_),
    .B(_03279_),
    .Y(_03290_));
 sky130_fd_sc_hd__a211o_1 _06658_ (.A1(_03257_),
    .A2(_02124_),
    .B1(_02135_),
    .C1(_03290_),
    .X(_03301_));
 sky130_fd_sc_hd__inv_2 _06659_ (.A(_03301_),
    .Y(_00009_));
 sky130_fd_sc_hd__or2_1 _06660_ (.A(net195),
    .B(_01128_),
    .X(_03322_));
 sky130_fd_sc_hd__o21a_1 _06661_ (.A1(_01358_),
    .A2(net219),
    .B1(_03322_),
    .X(_03333_));
 sky130_fd_sc_hd__a21oi_1 _06662_ (.A1(_01478_),
    .A2(_01544_),
    .B1(net220),
    .Y(_03344_));
 sky130_fd_sc_hd__inv_2 _06663_ (.A(net220),
    .Y(_03355_));
 sky130_fd_sc_hd__and2_1 _06664_ (.A(_03203_),
    .B(_03355_),
    .X(_03366_));
 sky130_fd_sc_hd__nand2_1 _06665_ (.A(_03028_),
    .B(_03148_),
    .Y(_03377_));
 sky130_fd_sc_hd__nor2_1 _06666_ (.A(_03355_),
    .B(_03377_),
    .Y(_03388_));
 sky130_fd_sc_hd__or2_1 _06667_ (.A(_03366_),
    .B(_03388_),
    .X(_03399_));
 sky130_fd_sc_hd__and2_1 _06668_ (.A(_03399_),
    .B(_01992_),
    .X(_03410_));
 sky130_fd_sc_hd__and2_1 _06669_ (.A(_03399_),
    .B(_02036_),
    .X(_03421_));
 sky130_fd_sc_hd__or3_1 _06670_ (.A(_03344_),
    .B(_03410_),
    .C(_03421_),
    .X(_03432_));
 sky130_fd_sc_hd__nor2_1 _06671_ (.A(net220),
    .B(_02178_),
    .Y(_03443_));
 sky130_fd_sc_hd__a21oi_1 _06672_ (.A1(_03399_),
    .A2(_02178_),
    .B1(_03443_),
    .Y(_03454_));
 sky130_fd_sc_hd__nor2_1 _06673_ (.A(_02113_),
    .B(net221),
    .Y(_03465_));
 sky130_fd_sc_hd__a211o_1 _06674_ (.A1(_03432_),
    .A2(_02146_),
    .B1(_02135_),
    .C1(net222),
    .X(_03476_));
 sky130_fd_sc_hd__inv_2 _06675_ (.A(net223),
    .Y(_00010_));
 sky130_fd_sc_hd__mux2_1 _06676_ (.A0(net195),
    .A1(net242),
    .S(_01358_),
    .X(_03496_));
 sky130_fd_sc_hd__inv_2 _06677_ (.A(net196),
    .Y(_03507_));
 sky130_fd_sc_hd__and2_1 _06678_ (.A(net256),
    .B(net220),
    .X(_03518_));
 sky130_fd_sc_hd__nand2_1 _06679_ (.A(_03181_),
    .B(_03518_),
    .Y(_03529_));
 sky130_fd_sc_hd__or2_1 _06680_ (.A(_03507_),
    .B(net257),
    .X(_03540_));
 sky130_fd_sc_hd__nand2_1 _06681_ (.A(net257),
    .B(_03507_),
    .Y(_03551_));
 sky130_fd_sc_hd__nand2_1 _06682_ (.A(_03540_),
    .B(_03551_),
    .Y(_03562_));
 sky130_fd_sc_hd__and2_1 _06683_ (.A(_03562_),
    .B(_01522_),
    .X(_03573_));
 sky130_fd_sc_hd__and2_1 _06684_ (.A(_02025_),
    .B(_03562_),
    .X(_03584_));
 sky130_fd_sc_hd__a21oi_1 _06685_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net196),
    .Y(_03595_));
 sky130_fd_sc_hd__or3_1 _06686_ (.A(_03573_),
    .B(_03584_),
    .C(_03595_),
    .X(_03606_));
 sky130_fd_sc_hd__nor2_1 _06687_ (.A(_02157_),
    .B(net196),
    .Y(_03617_));
 sky130_fd_sc_hd__a21oi_1 _06688_ (.A1(_03562_),
    .A2(_02178_),
    .B1(_03617_),
    .Y(_03628_));
 sky130_fd_sc_hd__nor2_1 _06689_ (.A(_02113_),
    .B(_03628_),
    .Y(_03639_));
 sky130_fd_sc_hd__a211o_1 _06690_ (.A1(_03606_),
    .A2(_02146_),
    .B1(_02135_),
    .C1(_03639_),
    .X(_03650_));
 sky130_fd_sc_hd__inv_2 _06691_ (.A(_03650_),
    .Y(_00011_));
 sky130_fd_sc_hd__or2_1 _06692_ (.A(net168),
    .B(_01128_),
    .X(_03671_));
 sky130_fd_sc_hd__o21a_1 _06693_ (.A1(_01358_),
    .A2(net242),
    .B1(_03671_),
    .X(_03682_));
 sky130_fd_sc_hd__a21oi_1 _06694_ (.A1(_01478_),
    .A2(_01544_),
    .B1(net243),
    .Y(_03693_));
 sky130_fd_sc_hd__inv_2 _06695_ (.A(net243),
    .Y(_03704_));
 sky130_fd_sc_hd__nand2_1 _06696_ (.A(_03388_),
    .B(net196),
    .Y(_03715_));
 sky130_fd_sc_hd__nor2_1 _06697_ (.A(_03704_),
    .B(_03715_),
    .Y(_03726_));
 sky130_fd_sc_hd__inv_2 _06698_ (.A(_03726_),
    .Y(_03736_));
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(_03540_),
    .B(_03704_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand2_1 _06700_ (.A(_03736_),
    .B(_03747_),
    .Y(_03758_));
 sky130_fd_sc_hd__and2_1 _06701_ (.A(_03758_),
    .B(_01992_),
    .X(_03769_));
 sky130_fd_sc_hd__and2_1 _06702_ (.A(_03758_),
    .B(_02036_),
    .X(_03780_));
 sky130_fd_sc_hd__or3_1 _06703_ (.A(_03693_),
    .B(_03769_),
    .C(_03780_),
    .X(_03791_));
 sky130_fd_sc_hd__nor2_1 _06704_ (.A(net243),
    .B(_02178_),
    .Y(_03802_));
 sky130_fd_sc_hd__a21oi_1 _06705_ (.A1(_03758_),
    .A2(_02178_),
    .B1(_03802_),
    .Y(_03813_));
 sky130_fd_sc_hd__nor2_1 _06706_ (.A(_02113_),
    .B(net244),
    .Y(_03824_));
 sky130_fd_sc_hd__a211o_1 _06707_ (.A1(_03791_),
    .A2(_02146_),
    .B1(net130),
    .C1(net245),
    .X(_03835_));
 sky130_fd_sc_hd__inv_2 _06708_ (.A(net246),
    .Y(_00012_));
 sky130_fd_sc_hd__mux2_1 _06709_ (.A0(net168),
    .A1(\M000[44] ),
    .S(_01358_),
    .X(_03856_));
 sky130_fd_sc_hd__inv_2 _06710_ (.A(net169),
    .Y(_03867_));
 sky130_fd_sc_hd__and3_1 _06711_ (.A(_03518_),
    .B(net196),
    .C(_03682_),
    .X(_03878_));
 sky130_fd_sc_hd__nand2_1 _06712_ (.A(_03181_),
    .B(net197),
    .Y(_03889_));
 sky130_fd_sc_hd__or2_1 _06713_ (.A(net170),
    .B(net198),
    .X(_03900_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(net198),
    .B(net170),
    .Y(_03911_));
 sky130_fd_sc_hd__nand2_1 _06715_ (.A(_03900_),
    .B(_03911_),
    .Y(_03922_));
 sky130_fd_sc_hd__and2_1 _06716_ (.A(_03922_),
    .B(_01522_),
    .X(_03933_));
 sky130_fd_sc_hd__and2_1 _06717_ (.A(_02025_),
    .B(_03922_),
    .X(_03944_));
 sky130_fd_sc_hd__a21oi_1 _06718_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net169),
    .Y(_03955_));
 sky130_fd_sc_hd__or3_1 _06719_ (.A(_03933_),
    .B(_03944_),
    .C(_03955_),
    .X(_03966_));
 sky130_fd_sc_hd__nor2_1 _06720_ (.A(_02157_),
    .B(net169),
    .Y(_03976_));
 sky130_fd_sc_hd__a21oi_1 _06721_ (.A1(_03922_),
    .A2(_02178_),
    .B1(_03976_),
    .Y(_03987_));
 sky130_fd_sc_hd__nor2_1 _06722_ (.A(_02113_),
    .B(net199),
    .Y(_03998_));
 sky130_fd_sc_hd__a211o_1 _06723_ (.A1(_03966_),
    .A2(_02146_),
    .B1(net130),
    .C1(net200),
    .X(_04009_));
 sky130_fd_sc_hd__inv_2 _06724_ (.A(net201),
    .Y(_00014_));
 sky130_fd_sc_hd__inv_2 _06725_ (.A(\M000[45] ),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_1 _06726_ (.A(_04030_),
    .B(_01358_),
    .Y(_04041_));
 sky130_fd_sc_hd__o21a_1 _06727_ (.A1(_01358_),
    .A2(net214),
    .B1(_04041_),
    .X(_04052_));
 sky130_fd_sc_hd__xor2_1 _06728_ (.A(net215),
    .B(_03900_),
    .X(_04063_));
 sky130_fd_sc_hd__nor2_1 _06729_ (.A(net215),
    .B(_02167_),
    .Y(_04074_));
 sky130_fd_sc_hd__a21oi_1 _06730_ (.A1(_04063_),
    .A2(_02167_),
    .B1(net216),
    .Y(_04085_));
 sky130_fd_sc_hd__or2_1 _06731_ (.A(net215),
    .B(_02058_),
    .X(_04096_));
 sky130_fd_sc_hd__nand2_1 _06732_ (.A(_04063_),
    .B(_01992_),
    .Y(_04107_));
 sky130_fd_sc_hd__nand2_1 _06733_ (.A(_04063_),
    .B(_02036_),
    .Y(_04118_));
 sky130_fd_sc_hd__inv_2 _06734_ (.A(net215),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_1 _06735_ (.A(_01533_),
    .B(_04129_),
    .Y(_04140_));
 sky130_fd_sc_hd__clkbuf_4 _06736_ (.A(_01336_),
    .X(_04151_));
 sky130_fd_sc_hd__a41o_1 _06737_ (.A1(_04096_),
    .A2(_04107_),
    .A3(_04118_),
    .A4(_04140_),
    .B1(_04151_),
    .X(_04162_));
 sky130_fd_sc_hd__o211ai_1 _06738_ (.A1(_02124_),
    .A2(net217),
    .B1(_03072_),
    .C1(_04162_),
    .Y(_04173_));
 sky130_fd_sc_hd__inv_2 _06739_ (.A(net218),
    .Y(_00015_));
 sky130_fd_sc_hd__nand2_1 _06740_ (.A(_01128_),
    .B(_04030_),
    .Y(_04194_));
 sky130_fd_sc_hd__o21a_1 _06741_ (.A1(_01128_),
    .A2(net149),
    .B1(_04194_),
    .X(_04205_));
 sky130_fd_sc_hd__inv_2 _06742_ (.A(net150),
    .Y(_04215_));
 sky130_fd_sc_hd__or3_1 _06743_ (.A(_03867_),
    .B(_04129_),
    .C(net198),
    .X(_04226_));
 sky130_fd_sc_hd__or2_1 _06744_ (.A(_04215_),
    .B(_04226_),
    .X(_04237_));
 sky130_fd_sc_hd__nand2_1 _06745_ (.A(_04226_),
    .B(_04215_),
    .Y(_04248_));
 sky130_fd_sc_hd__nand2_1 _06746_ (.A(_04237_),
    .B(_04248_),
    .Y(_04259_));
 sky130_fd_sc_hd__a21oi_1 _06747_ (.A1(_02058_),
    .A2(_02069_),
    .B1(net150),
    .Y(_04270_));
 sky130_fd_sc_hd__a21oi_1 _06748_ (.A1(_04259_),
    .A2(_02036_),
    .B1(net151),
    .Y(_04281_));
 sky130_fd_sc_hd__nand2_1 _06749_ (.A(_04259_),
    .B(_01992_),
    .Y(_04292_));
 sky130_fd_sc_hd__a21o_1 _06750_ (.A1(net152),
    .A2(_04292_),
    .B1(_04151_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_4 _06751_ (.A(_01511_),
    .X(_04314_));
 sky130_fd_sc_hd__mux2_1 _06752_ (.A0(_04259_),
    .A1(_04215_),
    .S(_04314_),
    .X(_04325_));
 sky130_fd_sc_hd__nand2_1 _06753_ (.A(_04325_),
    .B(_04151_),
    .Y(_04336_));
 sky130_fd_sc_hd__nand2_1 _06754_ (.A(net120),
    .B(_01588_),
    .Y(_04347_));
 sky130_fd_sc_hd__inv_2 _06755_ (.A(net121),
    .Y(_00001_));
 sky130_fd_sc_hd__a31o_1 _06756_ (.A1(net153),
    .A2(_04336_),
    .A3(_03072_),
    .B1(net122),
    .X(_00016_));
 sky130_fd_sc_hd__clkbuf_4 _06757_ (.A(net130),
    .X(_04378_));
 sky130_fd_sc_hd__nor2_1 _06758_ (.A(_04378_),
    .B(net158),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_1 _06759_ (.A(net16),
    .B(net48),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2_1 _06760_ (.A(net16),
    .B(net48),
    .Y(_04410_));
 sky130_fd_sc_hd__nor2b_4 _06761_ (.A(_04399_),
    .B_N(_04410_),
    .Y(_04420_));
 sky130_fd_sc_hd__or2_1 _06762_ (.A(net165),
    .B(_04420_),
    .X(_04431_));
 sky130_fd_sc_hd__inv_2 _06763_ (.A(net17),
    .Y(_04442_));
 sky130_fd_sc_hd__inv_2 _06764_ (.A(net49),
    .Y(_04453_));
 sky130_fd_sc_hd__nand2_1 _06765_ (.A(_04442_),
    .B(_04453_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2_1 _06766_ (.A(net17),
    .B(net49),
    .Y(_04475_));
 sky130_fd_sc_hd__nand2_1 _06767_ (.A(_04464_),
    .B(_04475_),
    .Y(_04486_));
 sky130_fd_sc_hd__or2_1 _06768_ (.A(_04399_),
    .B(_04486_),
    .X(_04497_));
 sky130_fd_sc_hd__nand2_1 _06769_ (.A(_04486_),
    .B(_04399_),
    .Y(_04508_));
 sky130_fd_sc_hd__nand2_4 _06770_ (.A(_04497_),
    .B(_04508_),
    .Y(_04519_));
 sky130_fd_sc_hd__or2_1 _06771_ (.A(_04431_),
    .B(_04519_),
    .X(_04530_));
 sky130_fd_sc_hd__inv_2 _06772_ (.A(net18),
    .Y(_04541_));
 sky130_fd_sc_hd__inv_2 _06773_ (.A(net50),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(_04541_),
    .B(_04552_),
    .Y(_04563_));
 sky130_fd_sc_hd__nand2_1 _06775_ (.A(net18),
    .B(net50),
    .Y(_04574_));
 sky130_fd_sc_hd__nand2_1 _06776_ (.A(_04563_),
    .B(_04574_),
    .Y(_04585_));
 sky130_fd_sc_hd__or2_1 _06777_ (.A(_04475_),
    .B(_04585_),
    .X(_04596_));
 sky130_fd_sc_hd__nand2_1 _06778_ (.A(_04585_),
    .B(_04475_),
    .Y(_04607_));
 sky130_fd_sc_hd__nand2_1 _06779_ (.A(_04596_),
    .B(_04607_),
    .Y(_04617_));
 sky130_fd_sc_hd__or2_1 _06780_ (.A(_04497_),
    .B(_04617_),
    .X(_04628_));
 sky130_fd_sc_hd__nand2_1 _06781_ (.A(_04617_),
    .B(_04497_),
    .Y(_04639_));
 sky130_fd_sc_hd__nand2_4 _06782_ (.A(_04628_),
    .B(_04639_),
    .Y(_04650_));
 sky130_fd_sc_hd__or2_1 _06783_ (.A(_04530_),
    .B(_04650_),
    .X(_04661_));
 sky130_fd_sc_hd__inv_2 _06784_ (.A(net19),
    .Y(_04672_));
 sky130_fd_sc_hd__inv_2 _06785_ (.A(net51),
    .Y(_04683_));
 sky130_fd_sc_hd__nand2_1 _06786_ (.A(_04672_),
    .B(_04683_),
    .Y(_04694_));
 sky130_fd_sc_hd__nand2_1 _06787_ (.A(net19),
    .B(net51),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_1 _06788_ (.A(_04694_),
    .B(_04705_),
    .Y(_04716_));
 sky130_fd_sc_hd__or2_1 _06789_ (.A(_04574_),
    .B(_04716_),
    .X(_04727_));
 sky130_fd_sc_hd__nand2_1 _06790_ (.A(_04716_),
    .B(_04574_),
    .Y(_04738_));
 sky130_fd_sc_hd__nand2_1 _06791_ (.A(_04727_),
    .B(_04738_),
    .Y(_04749_));
 sky130_fd_sc_hd__inv_2 _06792_ (.A(_04749_),
    .Y(_04760_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(_04628_),
    .B(_04596_),
    .Y(_04771_));
 sky130_fd_sc_hd__or2_1 _06794_ (.A(_04760_),
    .B(_04771_),
    .X(_04782_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(_04771_),
    .B(_04760_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand2_4 _06796_ (.A(_04782_),
    .B(_04792_),
    .Y(_04803_));
 sky130_fd_sc_hd__or2_1 _06797_ (.A(_04661_),
    .B(_04803_),
    .X(_04814_));
 sky130_fd_sc_hd__nand2_1 _06798_ (.A(_04803_),
    .B(_04661_),
    .Y(_04825_));
 sky130_fd_sc_hd__nand2_1 _06799_ (.A(_04814_),
    .B(_04825_),
    .Y(_04836_));
 sky130_fd_sc_hd__nand2_1 _06800_ (.A(_04519_),
    .B(_04431_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand2_2 _06801_ (.A(_04530_),
    .B(_04847_),
    .Y(_04858_));
 sky130_fd_sc_hd__nand2_1 _06802_ (.A(_04650_),
    .B(_04530_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_2 _06803_ (.A(_04661_),
    .B(_04869_),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _06804_ (.A(_04858_),
    .B(_04880_),
    .Y(_04891_));
 sky130_fd_sc_hd__inv_2 _06805_ (.A(_04891_),
    .Y(_04902_));
 sky130_fd_sc_hd__nor2_1 _06806_ (.A(_04129_),
    .B(_03867_),
    .Y(_04913_));
 sky130_fd_sc_hd__nand2_1 _06807_ (.A(_04420_),
    .B(_01128_),
    .Y(_04924_));
 sky130_fd_sc_hd__nand2_2 _06808_ (.A(_04431_),
    .B(_04924_),
    .Y(_04935_));
 sky130_fd_sc_hd__inv_2 _06809_ (.A(_04935_),
    .Y(_04946_));
 sky130_fd_sc_hd__and4_1 _06810_ (.A(_03878_),
    .B(net150),
    .C(net171),
    .D(_04946_),
    .X(_04956_));
 sky130_fd_sc_hd__nand2_1 _06811_ (.A(_03181_),
    .B(net172),
    .Y(_04967_));
 sky130_fd_sc_hd__or2_1 _06812_ (.A(_04902_),
    .B(net173),
    .X(_04978_));
 sky130_fd_sc_hd__or2_1 _06813_ (.A(_04836_),
    .B(_04978_),
    .X(_04989_));
 sky130_fd_sc_hd__nand2_1 _06814_ (.A(_04978_),
    .B(_04836_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _06815_ (.A(_04989_),
    .B(_05000_),
    .Y(_05011_));
 sky130_fd_sc_hd__inv_2 _06816_ (.A(_04836_),
    .Y(_05022_));
 sky130_fd_sc_hd__nand2_1 _06817_ (.A(_05022_),
    .B(_04314_),
    .Y(_05033_));
 sky130_fd_sc_hd__o21ai_1 _06818_ (.A1(_04314_),
    .A2(_05011_),
    .B1(_05033_),
    .Y(_05044_));
 sky130_fd_sc_hd__mux2_1 _06819_ (.A0(_05044_),
    .A1(_05022_),
    .S(_01500_),
    .X(_05055_));
 sky130_fd_sc_hd__nand2_1 _06820_ (.A(_01402_),
    .B(_05022_),
    .Y(_05066_));
 sky130_fd_sc_hd__o21ai_1 _06821_ (.A1(net158),
    .A2(_05011_),
    .B1(_05066_),
    .Y(_05077_));
 sky130_fd_sc_hd__mux2_1 _06822_ (.A0(_05055_),
    .A1(_05077_),
    .S(_01468_),
    .X(_05088_));
 sky130_fd_sc_hd__mux2_1 _06823_ (.A0(_05088_),
    .A1(net174),
    .S(_01336_),
    .X(_05098_));
 sky130_fd_sc_hd__nand2_1 _06824_ (.A(net20),
    .B(net52),
    .Y(_05109_));
 sky130_fd_sc_hd__or2_1 _06825_ (.A(net21),
    .B(net53),
    .X(_05120_));
 sky130_fd_sc_hd__nand2_1 _06826_ (.A(net21),
    .B(net53),
    .Y(_05131_));
 sky130_fd_sc_hd__nand2_1 _06827_ (.A(_05120_),
    .B(_05131_),
    .Y(_05142_));
 sky130_fd_sc_hd__or2_1 _06828_ (.A(_05109_),
    .B(_05142_),
    .X(_05153_));
 sky130_fd_sc_hd__nand2_1 _06829_ (.A(_05142_),
    .B(_05109_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_2 _06830_ (.A(_05153_),
    .B(_05164_),
    .Y(_05175_));
 sky130_fd_sc_hd__nand2_1 _06831_ (.A(_04792_),
    .B(_04727_),
    .Y(_05186_));
 sky130_fd_sc_hd__inv_2 _06832_ (.A(net20),
    .Y(_05197_));
 sky130_fd_sc_hd__inv_2 _06833_ (.A(net52),
    .Y(_05208_));
 sky130_fd_sc_hd__nand2_1 _06834_ (.A(_05197_),
    .B(_05208_),
    .Y(_05219_));
 sky130_fd_sc_hd__nand2_1 _06835_ (.A(_05219_),
    .B(_05109_),
    .Y(_05230_));
 sky130_fd_sc_hd__or2_1 _06836_ (.A(_04705_),
    .B(_05230_),
    .X(_05240_));
 sky130_fd_sc_hd__nand2_1 _06837_ (.A(_05230_),
    .B(_04705_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_05240_),
    .B(_05251_),
    .Y(_05262_));
 sky130_fd_sc_hd__inv_2 _06839_ (.A(_05262_),
    .Y(_05273_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(_05186_),
    .B(_05273_),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2_2 _06841_ (.A(_05284_),
    .B(_05240_),
    .Y(_05295_));
 sky130_fd_sc_hd__xor2_4 _06842_ (.A(_05175_),
    .B(_05295_),
    .X(_05306_));
 sky130_fd_sc_hd__or2_1 _06843_ (.A(_05273_),
    .B(_05186_),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_4 _06844_ (.A(_05317_),
    .B(_05284_),
    .Y(_05328_));
 sky130_fd_sc_hd__or2_1 _06845_ (.A(_05328_),
    .B(_04814_),
    .X(_05339_));
 sky130_fd_sc_hd__or2_1 _06846_ (.A(_05306_),
    .B(_05339_),
    .X(_05350_));
 sky130_fd_sc_hd__or2_1 _06847_ (.A(net22),
    .B(net54),
    .X(_05360_));
 sky130_fd_sc_hd__nand2_2 _06848_ (.A(net22),
    .B(net54),
    .Y(_05371_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(_05360_),
    .B(_05371_),
    .Y(_05382_));
 sky130_fd_sc_hd__or2_1 _06850_ (.A(_05131_),
    .B(_05382_),
    .X(_05393_));
 sky130_fd_sc_hd__nand2_1 _06851_ (.A(_05382_),
    .B(_05131_),
    .Y(_05404_));
 sky130_fd_sc_hd__nand2_2 _06852_ (.A(_05393_),
    .B(_05404_),
    .Y(_05415_));
 sky130_fd_sc_hd__a21bo_2 _06853_ (.A1(_05295_),
    .A2(_05164_),
    .B1_N(_05153_),
    .X(_05426_));
 sky130_fd_sc_hd__xor2_4 _06854_ (.A(_05415_),
    .B(_05426_),
    .X(_05437_));
 sky130_fd_sc_hd__nor2_1 _06855_ (.A(_05350_),
    .B(_05437_),
    .Y(_05448_));
 sky130_fd_sc_hd__inv_2 _06856_ (.A(_05448_),
    .Y(_05459_));
 sky130_fd_sc_hd__nand2_1 _06857_ (.A(_05437_),
    .B(_05350_),
    .Y(_05470_));
 sky130_fd_sc_hd__nand2_2 _06858_ (.A(_05459_),
    .B(_05470_),
    .Y(_05480_));
 sky130_fd_sc_hd__o21ai_1 _06859_ (.A1(_01522_),
    .A2(_05480_),
    .B1(_02014_),
    .Y(_05491_));
 sky130_fd_sc_hd__inv_2 _06860_ (.A(_02025_),
    .Y(_05502_));
 sky130_fd_sc_hd__a21o_1 _06861_ (.A1(_05491_),
    .A2(_05502_),
    .B1(_01336_),
    .X(_05513_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(_05339_),
    .B(_05306_),
    .Y(_05524_));
 sky130_fd_sc_hd__nand2_2 _06863_ (.A(_05350_),
    .B(_05524_),
    .Y(_05535_));
 sky130_fd_sc_hd__nand2_1 _06864_ (.A(_04814_),
    .B(_05328_),
    .Y(_05546_));
 sky130_fd_sc_hd__nand2_1 _06865_ (.A(_05339_),
    .B(_05546_),
    .Y(_05557_));
 sky130_fd_sc_hd__or4_1 _06866_ (.A(_04836_),
    .B(_04902_),
    .C(net173),
    .D(_05557_),
    .X(_05568_));
 sky130_fd_sc_hd__or2_1 _06867_ (.A(_05535_),
    .B(_05568_),
    .X(_05578_));
 sky130_fd_sc_hd__or2_1 _06868_ (.A(_05480_),
    .B(_05578_),
    .X(_05589_));
 sky130_fd_sc_hd__nand2_1 _06869_ (.A(_05578_),
    .B(_05480_),
    .Y(_05600_));
 sky130_fd_sc_hd__inv_2 _06870_ (.A(_01435_),
    .Y(_05611_));
 sky130_fd_sc_hd__and3_1 _06871_ (.A(_01303_),
    .B(_01314_),
    .C(_01424_),
    .X(_05622_));
 sky130_fd_sc_hd__inv_2 _06872_ (.A(_05622_),
    .Y(_05633_));
 sky130_fd_sc_hd__nand2_1 _06873_ (.A(_01413_),
    .B(_01446_),
    .Y(_05644_));
 sky130_fd_sc_hd__o211a_2 _06874_ (.A1(_01446_),
    .A2(_05611_),
    .B1(_05633_),
    .C1(_05644_),
    .X(_05655_));
 sky130_fd_sc_hd__inv_2 _06875_ (.A(_05655_),
    .Y(_05665_));
 sky130_fd_sc_hd__a221o_1 _06876_ (.A1(net144),
    .A2(_05513_),
    .B1(_05589_),
    .B2(_05600_),
    .C1(_05665_),
    .X(_05676_));
 sky130_fd_sc_hd__a21bo_1 _06877_ (.A1(net146),
    .A2(_05480_),
    .B1_N(_05676_),
    .X(_05687_));
 sky130_fd_sc_hd__inv_2 _06878_ (.A(_05557_),
    .Y(_05698_));
 sky130_fd_sc_hd__or2_1 _06879_ (.A(_05557_),
    .B(_04989_),
    .X(_05709_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(_04989_),
    .B(_05557_),
    .Y(_05720_));
 sky130_fd_sc_hd__and3_1 _06881_ (.A(_05709_),
    .B(net133),
    .C(_05720_),
    .X(_05731_));
 sky130_fd_sc_hd__a21o_1 _06882_ (.A1(_01511_),
    .A2(_05698_),
    .B1(net134),
    .X(_05742_));
 sky130_fd_sc_hd__mux2_1 _06883_ (.A0(net135),
    .A1(_05698_),
    .S(_01500_),
    .X(_05752_));
 sky130_fd_sc_hd__inv_2 _06884_ (.A(net158),
    .Y(_05763_));
 sky130_fd_sc_hd__and3_1 _06885_ (.A(_05709_),
    .B(_05763_),
    .C(_05720_),
    .X(_05774_));
 sky130_fd_sc_hd__a21o_1 _06886_ (.A1(_01402_),
    .A2(_05698_),
    .B1(_05774_),
    .X(_05785_));
 sky130_fd_sc_hd__mux2_1 _06887_ (.A0(_05752_),
    .A1(_05785_),
    .S(_01468_),
    .X(_05796_));
 sky130_fd_sc_hd__and2_1 _06888_ (.A(net135),
    .B(_01336_),
    .X(_05807_));
 sky130_fd_sc_hd__a21oi_1 _06889_ (.A1(_05796_),
    .A2(_02113_),
    .B1(_05807_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _06890_ (.A(net147),
    .B(net136),
    .Y(_05828_));
 sky130_fd_sc_hd__inv_2 _06891_ (.A(_05535_),
    .Y(_05839_));
 sky130_fd_sc_hd__o21ai_1 _06892_ (.A1(_01522_),
    .A2(_05535_),
    .B1(_02014_),
    .Y(_05850_));
 sky130_fd_sc_hd__inv_2 _06893_ (.A(_05850_),
    .Y(_05861_));
 sky130_fd_sc_hd__o21ai_1 _06894_ (.A1(_02025_),
    .A2(_05861_),
    .B1(_02102_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand2_1 _06895_ (.A(_05568_),
    .B(_05535_),
    .Y(_05882_));
 sky130_fd_sc_hd__a221o_1 _06896_ (.A1(net144),
    .A2(_05872_),
    .B1(_05578_),
    .B2(_05882_),
    .C1(_05665_),
    .X(_05893_));
 sky130_fd_sc_hd__o21ai_2 _06897_ (.A1(net145),
    .A2(_05839_),
    .B1(_05893_),
    .Y(_05904_));
 sky130_fd_sc_hd__inv_2 _06898_ (.A(_05904_),
    .Y(_05915_));
 sky130_fd_sc_hd__inv_2 _06899_ (.A(_04880_),
    .Y(_05926_));
 sky130_fd_sc_hd__or2_1 _06900_ (.A(_04858_),
    .B(net173),
    .X(_05937_));
 sky130_fd_sc_hd__xor2_1 _06901_ (.A(_04880_),
    .B(_05937_),
    .X(_05947_));
 sky130_fd_sc_hd__mux2_1 _06902_ (.A0(_05926_),
    .A1(_05947_),
    .S(net145),
    .X(_05958_));
 sky130_fd_sc_hd__or2_1 _06903_ (.A(_04935_),
    .B(_04237_),
    .X(_05969_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(_04237_),
    .B(_04935_),
    .Y(_05980_));
 sky130_fd_sc_hd__nor2_1 _06905_ (.A(_02157_),
    .B(_04935_),
    .Y(_05990_));
 sky130_fd_sc_hd__a31o_1 _06906_ (.A1(_05969_),
    .A2(_02157_),
    .A3(_05980_),
    .B1(_05990_),
    .X(_06001_));
 sky130_fd_sc_hd__mux2_1 _06907_ (.A0(_06001_),
    .A1(_04946_),
    .S(_01500_),
    .X(_06012_));
 sky130_fd_sc_hd__nand2_1 _06908_ (.A(_06012_),
    .B(_02014_),
    .Y(_06023_));
 sky130_fd_sc_hd__nor2_1 _06909_ (.A(_04935_),
    .B(_05763_),
    .Y(_06033_));
 sky130_fd_sc_hd__a31o_1 _06910_ (.A1(_05969_),
    .A2(_05763_),
    .A3(_05980_),
    .B1(_06033_),
    .X(_06044_));
 sky130_fd_sc_hd__nand2_1 _06911_ (.A(net159),
    .B(_01468_),
    .Y(_06054_));
 sky130_fd_sc_hd__a21o_1 _06912_ (.A1(_06023_),
    .A2(net160),
    .B1(_01336_),
    .X(_06065_));
 sky130_fd_sc_hd__inv_2 _06913_ (.A(_04858_),
    .Y(_06075_));
 sky130_fd_sc_hd__nand2_1 _06914_ (.A(net173),
    .B(_04858_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_1 _06915_ (.A1(_01522_),
    .A2(_04858_),
    .B1(_02014_),
    .Y(_06086_));
 sky130_fd_sc_hd__inv_2 _06916_ (.A(_06086_),
    .Y(_06096_));
 sky130_fd_sc_hd__o21ai_1 _06917_ (.A1(_06096_),
    .A2(_02025_),
    .B1(_02113_),
    .Y(_06105_));
 sky130_fd_sc_hd__a221o_1 _06918_ (.A1(_05937_),
    .A2(_06083_),
    .B1(net144),
    .B2(_06105_),
    .C1(_05665_),
    .X(_06115_));
 sky130_fd_sc_hd__o21ai_1 _06919_ (.A1(net145),
    .A2(_06075_),
    .B1(_06115_),
    .Y(_06124_));
 sky130_fd_sc_hd__nand2_1 _06920_ (.A(_06001_),
    .B(_01336_),
    .Y(_06134_));
 sky130_fd_sc_hd__nand3_1 _06921_ (.A(net161),
    .B(_06124_),
    .C(_06134_),
    .Y(_06140_));
 sky130_fd_sc_hd__nor3_1 _06922_ (.A(_05915_),
    .B(net166),
    .C(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__nor3b_1 _06923_ (.A(net175),
    .B(_05828_),
    .C_N(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__xnor2_2 _06924_ (.A(net24),
    .B(net56),
    .Y(_06143_));
 sky130_fd_sc_hd__xor2_4 _06925_ (.A(_05371_),
    .B(_06143_),
    .X(_06144_));
 sky130_fd_sc_hd__a21bo_1 _06926_ (.A1(_05426_),
    .A2(_05404_),
    .B1_N(_05393_),
    .X(_06145_));
 sky130_fd_sc_hd__xor2_4 _06927_ (.A(_06144_),
    .B(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__xor2_2 _06928_ (.A(_05459_),
    .B(_06146_),
    .X(_06147_));
 sky130_fd_sc_hd__or3_1 _06929_ (.A(_05480_),
    .B(_05535_),
    .C(_05568_),
    .X(_06148_));
 sky130_fd_sc_hd__xor2_1 _06930_ (.A(_06147_),
    .B(_06148_),
    .X(_06149_));
 sky130_fd_sc_hd__inv_2 _06931_ (.A(_06147_),
    .Y(_06150_));
 sky130_fd_sc_hd__mux2_1 _06932_ (.A0(_06149_),
    .A1(_06150_),
    .S(_04314_),
    .X(_06151_));
 sky130_fd_sc_hd__nor2_1 _06933_ (.A(_01489_),
    .B(_06147_),
    .Y(_06152_));
 sky130_fd_sc_hd__a21oi_1 _06934_ (.A1(_06151_),
    .A2(_01489_),
    .B1(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__mux2_1 _06935_ (.A0(_06149_),
    .A1(_06150_),
    .S(net158),
    .X(_06154_));
 sky130_fd_sc_hd__nand2_1 _06936_ (.A(_06154_),
    .B(_01468_),
    .Y(_06155_));
 sky130_fd_sc_hd__o21ai_1 _06937_ (.A1(_01468_),
    .A2(_06153_),
    .B1(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__nand2_1 _06938_ (.A(_06151_),
    .B(_01336_),
    .Y(_06157_));
 sky130_fd_sc_hd__a21boi_2 _06939_ (.A1(_06156_),
    .A2(_02113_),
    .B1_N(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__inv_2 _06940_ (.A(_06158_),
    .Y(_06159_));
 sky130_fd_sc_hd__nand2_1 _06941_ (.A(_06142_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__or4_1 _06942_ (.A(_05926_),
    .B(_04946_),
    .C(_06075_),
    .D(_05022_),
    .X(_06161_));
 sky130_fd_sc_hd__or3_1 _06943_ (.A(_05839_),
    .B(_05698_),
    .C(_06161_),
    .X(_06162_));
 sky130_fd_sc_hd__or3b_1 _06944_ (.A(_06147_),
    .B(_06162_),
    .C_N(_05480_),
    .X(_06163_));
 sky130_fd_sc_hd__a21oi_1 _06945_ (.A1(_06160_),
    .A2(_06163_),
    .B1(_04378_),
    .Y(_00035_));
 sky130_fd_sc_hd__or2_1 _06946_ (.A(net136),
    .B(net147),
    .X(_06164_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(net161),
    .B(_06134_),
    .Y(_06165_));
 sky130_fd_sc_hd__nand3b_1 _06948_ (.A_N(_06124_),
    .B(net162),
    .C(net166),
    .Y(_06166_));
 sky130_fd_sc_hd__nor3b_1 _06949_ (.A(_05904_),
    .B(_06166_),
    .C_N(_05098_),
    .Y(_06167_));
 sky130_fd_sc_hd__nand3b_1 _06950_ (.A_N(_06164_),
    .B(_06167_),
    .C(_06158_),
    .Y(_06168_));
 sky130_fd_sc_hd__or4_1 _06951_ (.A(_04836_),
    .B(_04935_),
    .C(_04902_),
    .D(_05557_),
    .X(_06169_));
 sky130_fd_sc_hd__or4_1 _06952_ (.A(_05480_),
    .B(_05535_),
    .C(_06169_),
    .D(_06150_),
    .X(_06170_));
 sky130_fd_sc_hd__a21oi_1 _06953_ (.A1(_06168_),
    .A2(_06170_),
    .B1(_04378_),
    .Y(_00034_));
 sky130_fd_sc_hd__buf_6 _06954_ (.A(net41),
    .X(_06171_));
 sky130_fd_sc_hd__buf_4 _06955_ (.A(_06171_),
    .X(_06172_));
 sky130_fd_sc_hd__buf_6 _06956_ (.A(net40),
    .X(_06173_));
 sky130_fd_sc_hd__buf_4 _06957_ (.A(_06173_),
    .X(_06174_));
 sky130_fd_sc_hd__buf_6 _06958_ (.A(net43),
    .X(_06175_));
 sky130_fd_sc_hd__buf_4 _06959_ (.A(_06175_),
    .X(_06176_));
 sky130_fd_sc_hd__buf_6 _06960_ (.A(net42),
    .X(_06177_));
 sky130_fd_sc_hd__buf_6 _06961_ (.A(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__buf_6 _06962_ (.A(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__or4_4 _06963_ (.A(_06172_),
    .B(_06174_),
    .C(_06176_),
    .D(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__inv_2 _06964_ (.A(net48),
    .Y(_06181_));
 sky130_fd_sc_hd__inv_2 _06965_ (.A(net56),
    .Y(_06182_));
 sky130_fd_sc_hd__buf_6 _06966_ (.A(net47),
    .X(_06183_));
 sky130_fd_sc_hd__buf_6 _06967_ (.A(_06183_),
    .X(_06184_));
 sky130_fd_sc_hd__inv_2 _06968_ (.A(net46),
    .Y(_06185_));
 sky130_fd_sc_hd__buf_2 _06969_ (.A(_06185_),
    .X(_06186_));
 sky130_fd_sc_hd__buf_6 _06970_ (.A(net45),
    .X(_06187_));
 sky130_fd_sc_hd__inv_2 _06971_ (.A(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__nand2_2 _06972_ (.A(_06186_),
    .B(_06188_),
    .Y(_06189_));
 sky130_fd_sc_hd__or2_2 _06973_ (.A(_06184_),
    .B(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__or3_1 _06974_ (.A(_06181_),
    .B(_06182_),
    .C(_06190_),
    .X(_06191_));
 sky130_fd_sc_hd__nand2_1 _06975_ (.A(net53),
    .B(net54),
    .Y(_06192_));
 sky130_fd_sc_hd__or4_1 _06976_ (.A(_04453_),
    .B(_04552_),
    .C(_04683_),
    .D(_05208_),
    .X(_06193_));
 sky130_fd_sc_hd__or3_1 _06977_ (.A(net57),
    .B(_06192_),
    .C(_06193_),
    .X(_06194_));
 sky130_fd_sc_hd__buf_6 _06978_ (.A(net60),
    .X(_06195_));
 sky130_fd_sc_hd__buf_6 _06979_ (.A(_06195_),
    .X(_06196_));
 sky130_fd_sc_hd__buf_6 _06980_ (.A(net59),
    .X(_06197_));
 sky130_fd_sc_hd__buf_4 _06981_ (.A(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__clkbuf_8 _06982_ (.A(net62),
    .X(_06199_));
 sky130_fd_sc_hd__buf_6 _06983_ (.A(_06199_),
    .X(_06200_));
 sky130_fd_sc_hd__buf_6 _06984_ (.A(net61),
    .X(_06201_));
 sky130_fd_sc_hd__buf_6 _06985_ (.A(_06201_),
    .X(_06202_));
 sky130_fd_sc_hd__or4_1 _06986_ (.A(_06196_),
    .B(_06198_),
    .C(_06200_),
    .D(_06202_),
    .X(_06203_));
 sky130_fd_sc_hd__buf_4 _06987_ (.A(net44),
    .X(_06204_));
 sky130_fd_sc_hd__buf_4 _06988_ (.A(_06204_),
    .X(_06205_));
 sky130_fd_sc_hd__buf_4 _06989_ (.A(_06205_),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_4 _06990_ (.A(net33),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_4 _06991_ (.A(_06207_),
    .X(_06208_));
 sky130_fd_sc_hd__clkbuf_4 _06992_ (.A(_06208_),
    .X(_06209_));
 sky130_fd_sc_hd__buf_6 _06993_ (.A(net58),
    .X(_06210_));
 sky130_fd_sc_hd__buf_6 _06994_ (.A(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__buf_6 _06995_ (.A(_06211_),
    .X(_06212_));
 sky130_fd_sc_hd__buf_6 _06996_ (.A(net55),
    .X(_06213_));
 sky130_fd_sc_hd__buf_6 _06997_ (.A(_06213_),
    .X(_06214_));
 sky130_fd_sc_hd__buf_6 _06998_ (.A(_06214_),
    .X(_06215_));
 sky130_fd_sc_hd__or4_1 _06999_ (.A(_06206_),
    .B(_06209_),
    .C(_06212_),
    .D(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__buf_6 _07000_ (.A(net37),
    .X(_06217_));
 sky130_fd_sc_hd__buf_4 _07001_ (.A(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__buf_6 _07002_ (.A(net36),
    .X(_06219_));
 sky130_fd_sc_hd__buf_6 _07003_ (.A(_06219_),
    .X(_06220_));
 sky130_fd_sc_hd__buf_6 _07004_ (.A(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__buf_4 _07005_ (.A(net39),
    .X(_06222_));
 sky130_fd_sc_hd__buf_4 _07006_ (.A(net38),
    .X(_06223_));
 sky130_fd_sc_hd__or4_1 _07007_ (.A(_06218_),
    .B(_06221_),
    .C(_06222_),
    .D(_06223_),
    .X(_06224_));
 sky130_fd_sc_hd__buf_4 _07008_ (.A(net64),
    .X(_06225_));
 sky130_fd_sc_hd__buf_4 _07009_ (.A(net63),
    .X(_06226_));
 sky130_fd_sc_hd__buf_6 _07010_ (.A(net35),
    .X(_06227_));
 sky130_fd_sc_hd__buf_4 _07011_ (.A(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__buf_6 _07012_ (.A(net34),
    .X(_06229_));
 sky130_fd_sc_hd__buf_6 _07013_ (.A(_06229_),
    .X(_06230_));
 sky130_fd_sc_hd__buf_6 _07014_ (.A(_06230_),
    .X(_06231_));
 sky130_fd_sc_hd__or4_1 _07015_ (.A(_06225_),
    .B(_06226_),
    .C(_06228_),
    .D(_06231_),
    .X(_06232_));
 sky130_fd_sc_hd__or4_4 _07016_ (.A(_06203_),
    .B(_06216_),
    .C(_06224_),
    .D(_06232_),
    .X(_06233_));
 sky130_fd_sc_hd__buf_8 _07017_ (.A(net9),
    .X(_06234_));
 sky130_fd_sc_hd__buf_6 _07018_ (.A(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__buf_6 _07019_ (.A(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__buf_6 _07020_ (.A(net8),
    .X(_06237_));
 sky130_fd_sc_hd__buf_4 _07021_ (.A(_06237_),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_8 _07022_ (.A(net11),
    .X(_06239_));
 sky130_fd_sc_hd__buf_4 _07023_ (.A(_06239_),
    .X(_06240_));
 sky130_fd_sc_hd__clkbuf_8 _07024_ (.A(net10),
    .X(_06241_));
 sky130_fd_sc_hd__buf_6 _07025_ (.A(_06241_),
    .X(_06242_));
 sky130_fd_sc_hd__buf_6 _07026_ (.A(_06242_),
    .X(_06243_));
 sky130_fd_sc_hd__or4_4 _07027_ (.A(_06236_),
    .B(_06238_),
    .C(_06240_),
    .D(_06243_),
    .X(_06244_));
 sky130_fd_sc_hd__buf_4 _07028_ (.A(net14),
    .X(_06245_));
 sky130_fd_sc_hd__buf_6 _07029_ (.A(_06245_),
    .X(_06246_));
 sky130_fd_sc_hd__buf_4 _07030_ (.A(_06246_),
    .X(_06247_));
 sky130_fd_sc_hd__buf_4 _07031_ (.A(net13),
    .X(_06248_));
 sky130_fd_sc_hd__nor2_2 _07032_ (.A(_06247_),
    .B(_06248_),
    .Y(_06249_));
 sky130_fd_sc_hd__clkinv_4 _07033_ (.A(net15),
    .Y(_06250_));
 sky130_fd_sc_hd__and2_1 _07034_ (.A(_06249_),
    .B(_06250_),
    .X(_06251_));
 sky130_fd_sc_hd__and3b_1 _07035_ (.A_N(_06244_),
    .B(net16),
    .C(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__inv_2 _07036_ (.A(_06252_),
    .Y(_06253_));
 sky130_fd_sc_hd__nand2_1 _07037_ (.A(net22),
    .B(net21),
    .Y(_06254_));
 sky130_fd_sc_hd__or4_1 _07038_ (.A(_04541_),
    .B(_04442_),
    .C(_05197_),
    .D(_04672_),
    .X(_06255_));
 sky130_fd_sc_hd__or3b_1 _07039_ (.A(_06254_),
    .B(_06255_),
    .C_N(net24),
    .X(_06256_));
 sky130_fd_sc_hd__or2_1 _07040_ (.A(net25),
    .B(_06256_),
    .X(_06257_));
 sky130_fd_sc_hd__buf_6 _07041_ (.A(net28),
    .X(_06258_));
 sky130_fd_sc_hd__buf_4 _07042_ (.A(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__buf_6 _07043_ (.A(net27),
    .X(_06260_));
 sky130_fd_sc_hd__buf_6 _07044_ (.A(_06260_),
    .X(_06261_));
 sky130_fd_sc_hd__buf_6 _07045_ (.A(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__buf_6 _07046_ (.A(net30),
    .X(_06263_));
 sky130_fd_sc_hd__buf_4 _07047_ (.A(_06263_),
    .X(_06264_));
 sky130_fd_sc_hd__buf_6 _07048_ (.A(net29),
    .X(_06265_));
 sky130_fd_sc_hd__buf_6 _07049_ (.A(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__or4_1 _07050_ (.A(_06259_),
    .B(_06262_),
    .C(_06264_),
    .D(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__buf_6 _07051_ (.A(net12),
    .X(_06268_));
 sky130_fd_sc_hd__buf_6 _07052_ (.A(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__buf_6 _07053_ (.A(net1),
    .X(_06270_));
 sky130_fd_sc_hd__buf_6 _07054_ (.A(_06270_),
    .X(_06271_));
 sky130_fd_sc_hd__buf_6 _07055_ (.A(net26),
    .X(_06272_));
 sky130_fd_sc_hd__buf_6 _07056_ (.A(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__buf_6 _07057_ (.A(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__buf_6 _07058_ (.A(net23),
    .X(_06275_));
 sky130_fd_sc_hd__buf_6 _07059_ (.A(_06275_),
    .X(_06276_));
 sky130_fd_sc_hd__or4_1 _07060_ (.A(_06269_),
    .B(_06271_),
    .C(_06274_),
    .D(_06276_),
    .X(_06277_));
 sky130_fd_sc_hd__clkbuf_8 _07061_ (.A(net5),
    .X(_06278_));
 sky130_fd_sc_hd__buf_4 _07062_ (.A(_06278_),
    .X(_06279_));
 sky130_fd_sc_hd__buf_4 _07063_ (.A(net4),
    .X(_06280_));
 sky130_fd_sc_hd__buf_8 _07064_ (.A(net7),
    .X(_06281_));
 sky130_fd_sc_hd__buf_4 _07065_ (.A(_06281_),
    .X(_06282_));
 sky130_fd_sc_hd__buf_6 _07066_ (.A(net6),
    .X(_06283_));
 sky130_fd_sc_hd__buf_4 _07067_ (.A(_06283_),
    .X(_06284_));
 sky130_fd_sc_hd__or4_1 _07068_ (.A(_06279_),
    .B(_06280_),
    .C(_06282_),
    .D(_06284_),
    .X(_06285_));
 sky130_fd_sc_hd__clkbuf_8 _07069_ (.A(net32),
    .X(_06286_));
 sky130_fd_sc_hd__buf_6 _07070_ (.A(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__buf_6 _07071_ (.A(_06287_),
    .X(_06288_));
 sky130_fd_sc_hd__buf_4 _07072_ (.A(net31),
    .X(_06289_));
 sky130_fd_sc_hd__buf_4 _07073_ (.A(_06289_),
    .X(_06290_));
 sky130_fd_sc_hd__buf_4 _07074_ (.A(net3),
    .X(_06291_));
 sky130_fd_sc_hd__buf_4 _07075_ (.A(net2),
    .X(_06292_));
 sky130_fd_sc_hd__or4_1 _07076_ (.A(_06288_),
    .B(_06290_),
    .C(_06291_),
    .D(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__or4_4 _07077_ (.A(_06267_),
    .B(_06277_),
    .C(_06285_),
    .D(_06293_),
    .X(_06294_));
 sky130_fd_sc_hd__or3_2 _07078_ (.A(_06253_),
    .B(_06257_),
    .C(_06294_),
    .X(_06295_));
 sky130_fd_sc_hd__o41a_1 _07079_ (.A1(_06180_),
    .A2(_06191_),
    .A3(_06194_),
    .A4(_06233_),
    .B1(_06295_),
    .X(_06296_));
 sky130_fd_sc_hd__or4_1 _07080_ (.A(net18),
    .B(net17),
    .C(net20),
    .D(net19),
    .X(_06297_));
 sky130_fd_sc_hd__buf_4 _07081_ (.A(net15),
    .X(_06298_));
 sky130_fd_sc_hd__clkbuf_8 _07082_ (.A(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__or3b_1 _07083_ (.A(_06299_),
    .B(net16),
    .C_N(_06249_),
    .X(_06300_));
 sky130_fd_sc_hd__or4_1 _07084_ (.A(net22),
    .B(net21),
    .C(net24),
    .D(_06244_),
    .X(_06301_));
 sky130_fd_sc_hd__or4_1 _07085_ (.A(_06297_),
    .B(_06300_),
    .C(_06301_),
    .D(_06294_),
    .X(_06302_));
 sky130_fd_sc_hd__or4_1 _07086_ (.A(net52),
    .B(net53),
    .C(net54),
    .D(net56),
    .X(_06303_));
 sky130_fd_sc_hd__or4_1 _07087_ (.A(net48),
    .B(net49),
    .C(net50),
    .D(net51),
    .X(_06304_));
 sky130_fd_sc_hd__or4_1 _07088_ (.A(_06190_),
    .B(_06180_),
    .C(_06303_),
    .D(_06304_),
    .X(_06305_));
 sky130_fd_sc_hd__nor2_1 _07089_ (.A(_06305_),
    .B(_06233_),
    .Y(_06306_));
 sky130_fd_sc_hd__inv_2 _07090_ (.A(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__and2_1 _07091_ (.A(_06302_),
    .B(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__inv_2 _07092_ (.A(_06308_),
    .Y(_06309_));
 sky130_fd_sc_hd__inv_2 _07093_ (.A(net25),
    .Y(_06310_));
 sky130_fd_sc_hd__or4_1 _07094_ (.A(_06310_),
    .B(_06253_),
    .C(_06256_),
    .D(_06294_),
    .X(_06311_));
 sky130_fd_sc_hd__a21o_1 _07095_ (.A1(_06311_),
    .A2(_06295_),
    .B1(_06307_),
    .X(_06312_));
 sky130_fd_sc_hd__o21ai_4 _07096_ (.A1(_06296_),
    .A2(_06309_),
    .B1(_06312_),
    .Y(inv_f_c));
 sky130_fd_sc_hd__nand2_4 _07097_ (.A(_06312_),
    .B(_06309_),
    .Y(\out_f_c[23] ));
 sky130_fd_sc_hd__inv_2 _07098_ (.A(net57),
    .Y(_06313_));
 sky130_fd_sc_hd__or3_1 _07099_ (.A(_06313_),
    .B(_06192_),
    .C(_06193_),
    .X(_06314_));
 sky130_fd_sc_hd__or4_2 _07100_ (.A(_06180_),
    .B(_06191_),
    .C(_06314_),
    .D(_06233_),
    .X(_06315_));
 sky130_fd_sc_hd__or4_1 _07101_ (.A(_06180_),
    .B(_06191_),
    .C(_06194_),
    .D(_06233_),
    .X(_06316_));
 sky130_fd_sc_hd__o2111ai_4 _07102_ (.A1(_06310_),
    .A2(_06315_),
    .B1(_06316_),
    .C1(_06295_),
    .D1(_06308_),
    .Y(_06317_));
 sky130_fd_sc_hd__inv_2 _07103_ (.A(_06317_),
    .Y(\out_f_c[31] ));
 sky130_fd_sc_hd__nand2_1 _07104_ (.A(_06271_),
    .B(_06209_),
    .Y(_06318_));
 sky130_fd_sc_hd__inv_2 _07105_ (.A(_06318_),
    .Y(\m1.out[0] ));
 sky130_fd_sc_hd__nand2_1 _07106_ (.A(_06315_),
    .B(_06311_),
    .Y(_06319_));
 sky130_fd_sc_hd__or3b_4 _07107_ (.A(_06319_),
    .B(_06309_),
    .C_N(_06296_),
    .X(_06320_));
 sky130_fd_sc_hd__clkbuf_1 _07108_ (.A(_06320_),
    .X(forward_c));
 sky130_fd_sc_hd__nand2_1 _07109_ (.A(_06269_),
    .B(_06209_),
    .Y(_06321_));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(_06271_),
    .B(_06206_),
    .Y(_06322_));
 sky130_fd_sc_hd__nor2_1 _07111_ (.A(_06321_),
    .B(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2_1 _07112_ (.A(_06321_),
    .B(_06322_),
    .Y(_06324_));
 sky130_fd_sc_hd__and2b_1 _07113_ (.A_N(_06323_),
    .B(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__clkbuf_1 _07114_ (.A(_06325_),
    .X(\m1.out[1] ));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(_06276_),
    .B(_06209_),
    .Y(_06326_));
 sky130_fd_sc_hd__buf_6 _07116_ (.A(_06268_),
    .X(_06327_));
 sky130_fd_sc_hd__inv_4 _07117_ (.A(_06327_),
    .Y(_06328_));
 sky130_fd_sc_hd__inv_2 _07118_ (.A(net1),
    .Y(_06329_));
 sky130_fd_sc_hd__inv_2 _07119_ (.A(_06204_),
    .Y(_06330_));
 sky130_fd_sc_hd__inv_2 _07120_ (.A(_06214_),
    .Y(_06331_));
 sky130_fd_sc_hd__or4_1 _07121_ (.A(_06328_),
    .B(_06329_),
    .C(_06330_),
    .D(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__a22o_1 _07122_ (.A1(_06269_),
    .A2(_06206_),
    .B1(_06271_),
    .B2(_06215_),
    .X(_06333_));
 sky130_fd_sc_hd__nand2_1 _07123_ (.A(_06332_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__xnor2_1 _07124_ (.A(_06326_),
    .B(_06334_),
    .Y(_06335_));
 sky130_fd_sc_hd__inv_2 _07125_ (.A(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__or2_1 _07126_ (.A(_06323_),
    .B(_06336_),
    .X(_06337_));
 sky130_fd_sc_hd__nand2_1 _07127_ (.A(_06336_),
    .B(_06323_),
    .Y(_06338_));
 sky130_fd_sc_hd__and2_1 _07128_ (.A(_06337_),
    .B(_06338_),
    .X(_06339_));
 sky130_fd_sc_hd__clkbuf_1 _07129_ (.A(_06339_),
    .X(\m1.out[2] ));
 sky130_fd_sc_hd__nand2_1 _07130_ (.A(_06274_),
    .B(_06209_),
    .Y(_06340_));
 sky130_fd_sc_hd__inv_2 _07131_ (.A(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand2_1 _07132_ (.A(_06276_),
    .B(_06206_),
    .Y(_06342_));
 sky130_fd_sc_hd__inv_2 _07133_ (.A(_06342_),
    .Y(_06343_));
 sky130_fd_sc_hd__and4_1 _07134_ (.A(_06269_),
    .B(_06271_),
    .C(_06212_),
    .D(_06215_),
    .X(_06344_));
 sky130_fd_sc_hd__a22o_1 _07135_ (.A1(_06269_),
    .A2(_06215_),
    .B1(_06271_),
    .B2(_06212_),
    .X(_06345_));
 sky130_fd_sc_hd__or2b_1 _07136_ (.A(_06344_),
    .B_N(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__xor2_2 _07137_ (.A(_06343_),
    .B(_06346_),
    .X(_06347_));
 sky130_fd_sc_hd__o21a_1 _07138_ (.A1(_06326_),
    .A2(_06334_),
    .B1(_06332_),
    .X(_06348_));
 sky130_fd_sc_hd__xnor2_1 _07139_ (.A(_06347_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__xor2_1 _07140_ (.A(_06341_),
    .B(_06349_),
    .X(_06350_));
 sky130_fd_sc_hd__or2_1 _07141_ (.A(_06338_),
    .B(_06350_),
    .X(_06351_));
 sky130_fd_sc_hd__nand2_1 _07142_ (.A(_06350_),
    .B(_06338_),
    .Y(_06352_));
 sky130_fd_sc_hd__and2_1 _07143_ (.A(_06351_),
    .B(_06352_),
    .X(_06353_));
 sky130_fd_sc_hd__clkbuf_1 _07144_ (.A(_06353_),
    .X(\m1.out[3] ));
 sky130_fd_sc_hd__and4_1 _07145_ (.A(_06274_),
    .B(_06262_),
    .C(_06206_),
    .D(_06208_),
    .X(_06354_));
 sky130_fd_sc_hd__inv_2 _07146_ (.A(_06354_),
    .Y(_06355_));
 sky130_fd_sc_hd__a22o_1 _07147_ (.A1(_06274_),
    .A2(_06206_),
    .B1(_06262_),
    .B2(_06209_),
    .X(_06356_));
 sky130_fd_sc_hd__and2_1 _07148_ (.A(_06355_),
    .B(_06356_),
    .X(_06357_));
 sky130_fd_sc_hd__a21oi_1 _07149_ (.A1(_06345_),
    .A2(_06343_),
    .B1(_06344_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand2_1 _07150_ (.A(_06276_),
    .B(_06215_),
    .Y(_06359_));
 sky130_fd_sc_hd__and4_1 _07151_ (.A(_06269_),
    .B(_06271_),
    .C(_06212_),
    .D(_06198_),
    .X(_06360_));
 sky130_fd_sc_hd__a22o_1 _07152_ (.A1(_06269_),
    .A2(_06212_),
    .B1(_06271_),
    .B2(_06198_),
    .X(_06361_));
 sky130_fd_sc_hd__nor2b_1 _07153_ (.A(_06360_),
    .B_N(_06361_),
    .Y(_06362_));
 sky130_fd_sc_hd__xor2_1 _07154_ (.A(_06359_),
    .B(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__nor2_1 _07155_ (.A(_06358_),
    .B(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__nand2_1 _07156_ (.A(_06363_),
    .B(_06358_),
    .Y(_06365_));
 sky130_fd_sc_hd__nand2b_1 _07157_ (.A_N(_06364_),
    .B(_06365_),
    .Y(_06366_));
 sky130_fd_sc_hd__xor2_1 _07158_ (.A(_06357_),
    .B(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nand2_1 _07159_ (.A(_06348_),
    .B(_06347_),
    .Y(_06368_));
 sky130_fd_sc_hd__nor2_1 _07160_ (.A(_06347_),
    .B(_06348_),
    .Y(_06369_));
 sky130_fd_sc_hd__a21oi_1 _07161_ (.A1(_06368_),
    .A2(_06341_),
    .B1(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_1 _07162_ (.A(_06367_),
    .B(_06370_),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2_1 _07163_ (.A(_06370_),
    .B(_06367_),
    .Y(_06372_));
 sky130_fd_sc_hd__nand2b_1 _07164_ (.A_N(_06371_),
    .B(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__nor2_1 _07165_ (.A(_06373_),
    .B(_06351_),
    .Y(_06374_));
 sky130_fd_sc_hd__and2_1 _07166_ (.A(_06351_),
    .B(_06373_),
    .X(_06375_));
 sky130_fd_sc_hd__nor2_1 _07167_ (.A(_06374_),
    .B(_06375_),
    .Y(\m1.out[4] ));
 sky130_fd_sc_hd__a21oi_1 _07168_ (.A1(_06365_),
    .A2(_06357_),
    .B1(_06364_),
    .Y(_06376_));
 sky130_fd_sc_hd__nand2_1 _07169_ (.A(_06259_),
    .B(_06208_),
    .Y(_06377_));
 sky130_fd_sc_hd__inv_2 _07170_ (.A(_06273_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_1 _07171_ (.A(_06262_),
    .B(_06205_),
    .Y(_06379_));
 sky130_fd_sc_hd__or3_1 _07172_ (.A(_06378_),
    .B(_06331_),
    .C(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__o21ai_1 _07173_ (.A1(_06378_),
    .A2(_06331_),
    .B1(_06379_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _07174_ (.A(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__xnor2_1 _07175_ (.A(_06377_),
    .B(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__inv_2 _07176_ (.A(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__inv_2 _07177_ (.A(_06359_),
    .Y(_06385_));
 sky130_fd_sc_hd__a21oi_1 _07178_ (.A1(_06361_),
    .A2(_06385_),
    .B1(_06360_),
    .Y(_06386_));
 sky130_fd_sc_hd__inv_2 _07179_ (.A(_06195_),
    .Y(_06387_));
 sky130_fd_sc_hd__nand2_1 _07180_ (.A(_06327_),
    .B(_06198_),
    .Y(_06388_));
 sky130_fd_sc_hd__nor3_1 _07181_ (.A(_06329_),
    .B(_06387_),
    .C(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__o21ai_2 _07182_ (.A1(_06329_),
    .A2(_06387_),
    .B1(_06388_),
    .Y(_06390_));
 sky130_fd_sc_hd__inv_2 _07183_ (.A(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__buf_4 _07184_ (.A(_06275_),
    .X(_06392_));
 sky130_fd_sc_hd__nand2_1 _07185_ (.A(_06392_),
    .B(_06211_),
    .Y(_06393_));
 sky130_fd_sc_hd__o21ai_1 _07186_ (.A1(_06389_),
    .A2(_06391_),
    .B1(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__inv_2 _07187_ (.A(_06393_),
    .Y(_06395_));
 sky130_fd_sc_hd__nand3b_1 _07188_ (.A_N(_06389_),
    .B(_06395_),
    .C(_06390_),
    .Y(_06396_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(_06394_),
    .B(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__or2_1 _07190_ (.A(_06386_),
    .B(_06397_),
    .X(_06398_));
 sky130_fd_sc_hd__nand2_1 _07191_ (.A(_06397_),
    .B(_06386_),
    .Y(_06399_));
 sky130_fd_sc_hd__nand2_1 _07192_ (.A(_06398_),
    .B(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__xor2_1 _07193_ (.A(_06384_),
    .B(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__nor2_1 _07194_ (.A(_06376_),
    .B(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand2_1 _07195_ (.A(_06401_),
    .B(_06376_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2b_1 _07196_ (.A_N(_06402_),
    .B(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__nand2b_1 _07197_ (.A_N(_06404_),
    .B(_06354_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_1 _07198_ (.A(_06404_),
    .B(_06355_),
    .Y(_06406_));
 sky130_fd_sc_hd__a21o_1 _07199_ (.A1(_06405_),
    .A2(_06406_),
    .B1(_06371_),
    .X(_06407_));
 sky130_fd_sc_hd__nand3_2 _07200_ (.A(_06405_),
    .B(_06371_),
    .C(_06406_),
    .Y(_06408_));
 sky130_fd_sc_hd__a21oi_1 _07201_ (.A1(_06407_),
    .A2(_06408_),
    .B1(_06374_),
    .Y(_06409_));
 sky130_fd_sc_hd__nand3_1 _07202_ (.A(_06374_),
    .B(_06408_),
    .C(_06407_),
    .Y(_06410_));
 sky130_fd_sc_hd__and2b_1 _07203_ (.A_N(_06409_),
    .B(_06410_),
    .X(_06411_));
 sky130_fd_sc_hd__clkbuf_1 _07204_ (.A(_06411_),
    .X(\m1.out[5] ));
 sky130_fd_sc_hd__a21oi_1 _07205_ (.A1(_06403_),
    .A2(_06354_),
    .B1(_06402_),
    .Y(_06412_));
 sky130_fd_sc_hd__inv_2 _07206_ (.A(net61),
    .Y(_06413_));
 sky130_fd_sc_hd__nand2_1 _07207_ (.A(_06268_),
    .B(_06195_),
    .Y(_06414_));
 sky130_fd_sc_hd__nor3_1 _07208_ (.A(_06329_),
    .B(_06413_),
    .C(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__o21ai_2 _07209_ (.A1(_06329_),
    .A2(_06413_),
    .B1(_06414_),
    .Y(_06416_));
 sky130_fd_sc_hd__inv_2 _07210_ (.A(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__nand2_1 _07211_ (.A(_06275_),
    .B(_06197_),
    .Y(_06418_));
 sky130_fd_sc_hd__o21ai_1 _07212_ (.A1(_06415_),
    .A2(_06417_),
    .B1(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__inv_2 _07213_ (.A(_06418_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand3b_1 _07214_ (.A_N(_06415_),
    .B(_06420_),
    .C(_06416_),
    .Y(_06421_));
 sky130_fd_sc_hd__nand2_1 _07215_ (.A(_06419_),
    .B(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__a21oi_1 _07216_ (.A1(_06390_),
    .A2(_06395_),
    .B1(_06389_),
    .Y(_06423_));
 sky130_fd_sc_hd__nand2_1 _07217_ (.A(_06422_),
    .B(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand3b_1 _07218_ (.A_N(_06423_),
    .B(_06419_),
    .C(_06421_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _07219_ (.A(_06424_),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__nand2_1 _07220_ (.A(_06261_),
    .B(_06213_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand2_1 _07221_ (.A(_06273_),
    .B(_06210_),
    .Y(_06428_));
 sky130_fd_sc_hd__xor2_1 _07222_ (.A(_06427_),
    .B(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__a21o_1 _07223_ (.A1(_06259_),
    .A2(_06205_),
    .B1(_06429_),
    .X(_06430_));
 sky130_fd_sc_hd__nand3_1 _07224_ (.A(_06429_),
    .B(_06259_),
    .C(_06205_),
    .Y(_06431_));
 sky130_fd_sc_hd__nand2_1 _07225_ (.A(_06430_),
    .B(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__inv_2 _07226_ (.A(_06432_),
    .Y(_06433_));
 sky130_fd_sc_hd__nand2b_1 _07227_ (.A_N(_06426_),
    .B(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__nand2_1 _07228_ (.A(_06426_),
    .B(_06432_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_1 _07229_ (.A(_06434_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__a21boi_1 _07230_ (.A1(_06384_),
    .A2(_06399_),
    .B1_N(_06398_),
    .Y(_06437_));
 sky130_fd_sc_hd__nor2_1 _07231_ (.A(_06436_),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__nand2_1 _07232_ (.A(_06437_),
    .B(_06436_),
    .Y(_06439_));
 sky130_fd_sc_hd__inv_2 _07233_ (.A(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_1 _07234_ (.A(_06266_),
    .B(_06209_),
    .Y(_06441_));
 sky130_fd_sc_hd__o21a_1 _07235_ (.A1(_06377_),
    .A2(_06382_),
    .B1(_06380_),
    .X(_06442_));
 sky130_fd_sc_hd__nor2_1 _07236_ (.A(_06441_),
    .B(_06442_),
    .Y(_06443_));
 sky130_fd_sc_hd__inv_2 _07237_ (.A(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__nand2_1 _07238_ (.A(_06442_),
    .B(_06441_),
    .Y(_06445_));
 sky130_fd_sc_hd__and2_1 _07239_ (.A(_06444_),
    .B(_06445_),
    .X(_06446_));
 sky130_fd_sc_hd__o21bai_1 _07240_ (.A1(_06438_),
    .A2(_06440_),
    .B1_N(_06446_),
    .Y(_06447_));
 sky130_fd_sc_hd__nand3b_1 _07241_ (.A_N(_06438_),
    .B(_06446_),
    .C(_06439_),
    .Y(_06448_));
 sky130_fd_sc_hd__nand2_1 _07242_ (.A(_06447_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__nor2_1 _07243_ (.A(_06412_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__inv_2 _07244_ (.A(_06450_),
    .Y(_06451_));
 sky130_fd_sc_hd__nand2_1 _07245_ (.A(_06449_),
    .B(_06412_),
    .Y(_06452_));
 sky130_fd_sc_hd__nand2_1 _07246_ (.A(_06451_),
    .B(_06452_),
    .Y(_06453_));
 sky130_fd_sc_hd__nor2_1 _07247_ (.A(_06408_),
    .B(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__nand2_1 _07248_ (.A(_06453_),
    .B(_06408_),
    .Y(_06455_));
 sky130_fd_sc_hd__nand2b_1 _07249_ (.A_N(_06454_),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__nor2_1 _07250_ (.A(_06410_),
    .B(_06456_),
    .Y(_00036_));
 sky130_fd_sc_hd__and2_1 _07251_ (.A(_06456_),
    .B(_06410_),
    .X(_00037_));
 sky130_fd_sc_hd__nor2_1 _07252_ (.A(_00036_),
    .B(_00037_),
    .Y(\m1.out[6] ));
 sky130_fd_sc_hd__a21oi_1 _07253_ (.A1(_06439_),
    .A2(_06446_),
    .B1(_06438_),
    .Y(_00038_));
 sky130_fd_sc_hd__inv_2 _07254_ (.A(_00038_),
    .Y(_00039_));
 sky130_fd_sc_hd__nand2_1 _07255_ (.A(_06434_),
    .B(_06425_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _07256_ (.A(_06275_),
    .B(net60),
    .Y(_00041_));
 sky130_fd_sc_hd__nand2_1 _07257_ (.A(net12),
    .B(net61),
    .Y(_00042_));
 sky130_fd_sc_hd__nand2_1 _07258_ (.A(net1),
    .B(net62),
    .Y(_00043_));
 sky130_fd_sc_hd__nor2_1 _07259_ (.A(_00042_),
    .B(_00043_),
    .Y(_00044_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(_00042_),
    .B(_00043_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand2b_1 _07261_ (.A_N(_00044_),
    .B(_00045_),
    .Y(_00046_));
 sky130_fd_sc_hd__or2_1 _07262_ (.A(_00041_),
    .B(_00046_),
    .X(_00047_));
 sky130_fd_sc_hd__nand2_1 _07263_ (.A(_00046_),
    .B(_00041_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2_1 _07264_ (.A(_00047_),
    .B(_00048_),
    .Y(_00049_));
 sky130_fd_sc_hd__a21oi_1 _07265_ (.A1(_06416_),
    .A2(_06420_),
    .B1(_06415_),
    .Y(_00050_));
 sky130_fd_sc_hd__nand2_1 _07266_ (.A(_00049_),
    .B(_00050_),
    .Y(_00051_));
 sky130_fd_sc_hd__nand3b_1 _07267_ (.A_N(_00050_),
    .B(_00047_),
    .C(_00048_),
    .Y(_00052_));
 sky130_fd_sc_hd__nand2_1 _07268_ (.A(_00051_),
    .B(_00052_),
    .Y(_00053_));
 sky130_fd_sc_hd__nand2_1 _07269_ (.A(_06258_),
    .B(_06213_),
    .Y(_00054_));
 sky130_fd_sc_hd__inv_2 _07270_ (.A(_00054_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand2_1 _07271_ (.A(_06260_),
    .B(net58),
    .Y(_00056_));
 sky130_fd_sc_hd__nand2_1 _07272_ (.A(_06272_),
    .B(_06197_),
    .Y(_00057_));
 sky130_fd_sc_hd__nor2_1 _07273_ (.A(_00056_),
    .B(_00057_),
    .Y(_00058_));
 sky130_fd_sc_hd__nand2_1 _07274_ (.A(_00056_),
    .B(_00057_),
    .Y(_00059_));
 sky130_fd_sc_hd__or2b_1 _07275_ (.A(_00058_),
    .B_N(_00059_),
    .X(_00060_));
 sky130_fd_sc_hd__xor2_2 _07276_ (.A(_00055_),
    .B(_00060_),
    .X(_00061_));
 sky130_fd_sc_hd__nand2_1 _07277_ (.A(_00053_),
    .B(_00061_),
    .Y(_00062_));
 sky130_fd_sc_hd__or2_1 _07278_ (.A(_00061_),
    .B(_00053_),
    .X(_00063_));
 sky130_fd_sc_hd__nand3_2 _07279_ (.A(_00040_),
    .B(_00062_),
    .C(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__nand2_1 _07280_ (.A(_00063_),
    .B(_00062_),
    .Y(_00065_));
 sky130_fd_sc_hd__o21a_1 _07281_ (.A1(_06432_),
    .A2(_06426_),
    .B1(_06425_),
    .X(_00066_));
 sky130_fd_sc_hd__nand2_1 _07282_ (.A(_00065_),
    .B(_00066_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_1 _07283_ (.A(_00064_),
    .B(_00067_),
    .Y(_00068_));
 sky130_fd_sc_hd__clkinv_4 _07284_ (.A(_06265_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_1 _07285_ (.A(_06264_),
    .B(_06207_),
    .Y(_00070_));
 sky130_fd_sc_hd__nor3_1 _07286_ (.A(_00069_),
    .B(_06330_),
    .C(_00070_),
    .Y(_00071_));
 sky130_fd_sc_hd__inv_2 _07287_ (.A(_00071_),
    .Y(_00072_));
 sky130_fd_sc_hd__o21ai_1 _07288_ (.A1(_00069_),
    .A2(_06330_),
    .B1(_00070_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_1 _07289_ (.A(_00072_),
    .B(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__o21a_1 _07290_ (.A1(_06427_),
    .A2(_06428_),
    .B1(_06431_),
    .X(_00075_));
 sky130_fd_sc_hd__nor2_1 _07291_ (.A(_00074_),
    .B(_00075_),
    .Y(_00076_));
 sky130_fd_sc_hd__inv_2 _07292_ (.A(_00076_),
    .Y(_00077_));
 sky130_fd_sc_hd__nand2_1 _07293_ (.A(_00075_),
    .B(_00074_),
    .Y(_00078_));
 sky130_fd_sc_hd__nand2_1 _07294_ (.A(_00077_),
    .B(_00078_),
    .Y(_00079_));
 sky130_fd_sc_hd__nand2_1 _07295_ (.A(_00068_),
    .B(_00079_),
    .Y(_00080_));
 sky130_fd_sc_hd__inv_2 _07296_ (.A(_00079_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand3_2 _07297_ (.A(_00064_),
    .B(_00067_),
    .C(_00081_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand3_2 _07298_ (.A(_00039_),
    .B(_00080_),
    .C(_00082_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_1 _07299_ (.A(_00080_),
    .B(_00082_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _07300_ (.A(_00084_),
    .B(_00038_),
    .Y(_00085_));
 sky130_fd_sc_hd__nand2_1 _07301_ (.A(_00083_),
    .B(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_1 _07302_ (.A(_00086_),
    .B(_06444_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand3_1 _07303_ (.A(_00083_),
    .B(_00085_),
    .C(_06443_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_1 _07304_ (.A(_00087_),
    .B(_00088_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_1 _07305_ (.A(_00089_),
    .B(_06451_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand3_2 _07306_ (.A(_00087_),
    .B(_00088_),
    .C(_06450_),
    .Y(_00091_));
 sky130_fd_sc_hd__a21o_1 _07307_ (.A1(_00090_),
    .A2(_00091_),
    .B1(_06454_),
    .X(_00092_));
 sky130_fd_sc_hd__nand3_2 _07308_ (.A(_00090_),
    .B(_06454_),
    .C(_00091_),
    .Y(_00093_));
 sky130_fd_sc_hd__a21o_1 _07309_ (.A1(_00092_),
    .A2(_00093_),
    .B1(_00036_),
    .X(_00094_));
 sky130_fd_sc_hd__nand3_1 _07310_ (.A(_00036_),
    .B(_00093_),
    .C(_00092_),
    .Y(_00095_));
 sky130_fd_sc_hd__and2_1 _07311_ (.A(_00094_),
    .B(_00095_),
    .X(_00096_));
 sky130_fd_sc_hd__clkbuf_1 _07312_ (.A(_00096_),
    .X(\m1.out[7] ));
 sky130_fd_sc_hd__inv_2 _07313_ (.A(_00061_),
    .Y(_00097_));
 sky130_fd_sc_hd__a21boi_1 _07314_ (.A1(_00097_),
    .A2(_00051_),
    .B1_N(_00052_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_1 _07315_ (.A(_06268_),
    .B(net62),
    .Y(_00099_));
 sky130_fd_sc_hd__nand2_1 _07316_ (.A(net1),
    .B(net63),
    .Y(_00100_));
 sky130_fd_sc_hd__nor2_1 _07317_ (.A(_00099_),
    .B(_00100_),
    .Y(_00101_));
 sky130_fd_sc_hd__nand2_1 _07318_ (.A(_00099_),
    .B(_00100_),
    .Y(_00102_));
 sky130_fd_sc_hd__or2b_1 _07319_ (.A(_00101_),
    .B_N(_00102_),
    .X(_00103_));
 sky130_fd_sc_hd__nand2_1 _07320_ (.A(_06275_),
    .B(net61),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_1 _07321_ (.A(_00103_),
    .B(_00104_),
    .Y(_00105_));
 sky130_fd_sc_hd__inv_2 _07322_ (.A(_00104_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand3b_1 _07323_ (.A_N(_00101_),
    .B(_00102_),
    .C(_00106_),
    .Y(_00107_));
 sky130_fd_sc_hd__nand2_1 _07324_ (.A(_00105_),
    .B(_00107_),
    .Y(_00108_));
 sky130_fd_sc_hd__inv_2 _07325_ (.A(_00041_),
    .Y(_00109_));
 sky130_fd_sc_hd__a21oi_1 _07326_ (.A1(_00045_),
    .A2(_00109_),
    .B1(_00044_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_1 _07327_ (.A(_00108_),
    .B(_00110_),
    .Y(_00111_));
 sky130_fd_sc_hd__nand3b_1 _07328_ (.A_N(_00110_),
    .B(_00105_),
    .C(_00107_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _07329_ (.A(_06258_),
    .B(_06210_),
    .Y(_00113_));
 sky130_fd_sc_hd__inv_2 _07330_ (.A(_00113_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_1 _07331_ (.A(_06260_),
    .B(_06197_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_1 _07332_ (.A(_06272_),
    .B(net60),
    .Y(_00116_));
 sky130_fd_sc_hd__or2_1 _07333_ (.A(_00115_),
    .B(_00116_),
    .X(_00117_));
 sky130_fd_sc_hd__nand2_1 _07334_ (.A(_00115_),
    .B(_00116_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_1 _07335_ (.A(_00117_),
    .B(_00118_),
    .Y(_00119_));
 sky130_fd_sc_hd__xor2_1 _07336_ (.A(_00114_),
    .B(_00119_),
    .X(_00120_));
 sky130_fd_sc_hd__inv_2 _07337_ (.A(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__a21o_1 _07338_ (.A1(_00111_),
    .A2(_00112_),
    .B1(_00121_),
    .X(_00122_));
 sky130_fd_sc_hd__nand3_1 _07339_ (.A(_00121_),
    .B(_00111_),
    .C(_00112_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _07340_ (.A(_00122_),
    .B(_00123_),
    .Y(_00124_));
 sky130_fd_sc_hd__nor2_1 _07341_ (.A(_00098_),
    .B(_00124_),
    .Y(_00125_));
 sky130_fd_sc_hd__inv_2 _07342_ (.A(_00125_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(_00124_),
    .B(_00098_),
    .Y(_00127_));
 sky130_fd_sc_hd__nand2_1 _07344_ (.A(_00126_),
    .B(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__nand2_1 _07345_ (.A(_06263_),
    .B(net44),
    .Y(_00129_));
 sky130_fd_sc_hd__nand2_1 _07346_ (.A(net29),
    .B(_06213_),
    .Y(_00130_));
 sky130_fd_sc_hd__nor2_1 _07347_ (.A(_00129_),
    .B(_00130_),
    .Y(_00131_));
 sky130_fd_sc_hd__inv_2 _07348_ (.A(_00131_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _07349_ (.A(_00129_),
    .B(_00130_),
    .Y(_00133_));
 sky130_fd_sc_hd__nand2_1 _07350_ (.A(_06289_),
    .B(net33),
    .Y(_00134_));
 sky130_fd_sc_hd__inv_2 _07351_ (.A(_00134_),
    .Y(_00135_));
 sky130_fd_sc_hd__a21o_1 _07352_ (.A1(_00132_),
    .A2(_00133_),
    .B1(_00135_),
    .X(_00136_));
 sky130_fd_sc_hd__nand3_1 _07353_ (.A(_00132_),
    .B(_00133_),
    .C(_00135_),
    .Y(_00137_));
 sky130_fd_sc_hd__nand2_1 _07354_ (.A(_00136_),
    .B(_00137_),
    .Y(_00138_));
 sky130_fd_sc_hd__a21oi_1 _07355_ (.A1(_00059_),
    .A2(_00055_),
    .B1(_00058_),
    .Y(_00139_));
 sky130_fd_sc_hd__nand2_1 _07356_ (.A(_00138_),
    .B(_00139_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand3b_1 _07357_ (.A_N(_00139_),
    .B(_00136_),
    .C(_00137_),
    .Y(_00141_));
 sky130_fd_sc_hd__nand2_1 _07358_ (.A(_00140_),
    .B(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__or2_1 _07359_ (.A(_00072_),
    .B(_00142_),
    .X(_00143_));
 sky130_fd_sc_hd__nand2_1 _07360_ (.A(_00142_),
    .B(_00072_),
    .Y(_00144_));
 sky130_fd_sc_hd__nand2_1 _07361_ (.A(_00143_),
    .B(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__nand2_1 _07362_ (.A(_00128_),
    .B(_00145_),
    .Y(_00146_));
 sky130_fd_sc_hd__inv_2 _07363_ (.A(_00145_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand3_1 _07364_ (.A(_00126_),
    .B(_00127_),
    .C(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__nand2_1 _07365_ (.A(_00146_),
    .B(_00148_),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_2 _07366_ (.A(_00149_),
    .Y(_00150_));
 sky130_fd_sc_hd__nand2_1 _07367_ (.A(_00082_),
    .B(_00064_),
    .Y(_00151_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(_00150_),
    .B(_00151_),
    .Y(_00152_));
 sky130_fd_sc_hd__a21boi_1 _07369_ (.A1(_00081_),
    .A2(_00067_),
    .B1_N(_00064_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand2_1 _07370_ (.A(_00153_),
    .B(_00149_),
    .Y(_00154_));
 sky130_fd_sc_hd__nand3_1 _07371_ (.A(_00152_),
    .B(_00154_),
    .C(_00076_),
    .Y(_00155_));
 sky130_fd_sc_hd__nand2_1 _07372_ (.A(_00155_),
    .B(_00152_),
    .Y(_00156_));
 sky130_fd_sc_hd__a21oi_1 _07373_ (.A1(_00147_),
    .A2(_00127_),
    .B1(_00125_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand2_1 _07374_ (.A(_00123_),
    .B(_00112_),
    .Y(_00158_));
 sky130_fd_sc_hd__inv_2 _07375_ (.A(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__a21oi_1 _07376_ (.A1(_00102_),
    .A2(_00106_),
    .B1(_00101_),
    .Y(_00160_));
 sky130_fd_sc_hd__nand2_1 _07377_ (.A(_06268_),
    .B(net63),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _07378_ (.A(net1),
    .B(net64),
    .Y(_00162_));
 sky130_fd_sc_hd__nor2_1 _07379_ (.A(_00161_),
    .B(_00162_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _07380_ (.A(_00161_),
    .B(_00162_),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _07381_ (.A(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _07382_ (.A(_06275_),
    .B(_06199_),
    .Y(_00166_));
 sky130_fd_sc_hd__o21ai_1 _07383_ (.A1(_00163_),
    .A2(_00165_),
    .B1(_00166_),
    .Y(_00167_));
 sky130_fd_sc_hd__inv_2 _07384_ (.A(_00166_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand3b_1 _07385_ (.A_N(_00163_),
    .B(_00168_),
    .C(_00164_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand2_1 _07386_ (.A(_00167_),
    .B(_00169_),
    .Y(_00170_));
 sky130_fd_sc_hd__nor2_1 _07387_ (.A(_00160_),
    .B(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _07388_ (.A(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _07389_ (.A(_00170_),
    .B(_00160_),
    .Y(_00173_));
 sky130_fd_sc_hd__nand2_1 _07390_ (.A(_00172_),
    .B(_00173_),
    .Y(_00174_));
 sky130_fd_sc_hd__buf_6 _07391_ (.A(_06258_),
    .X(_00175_));
 sky130_fd_sc_hd__buf_4 _07392_ (.A(_06197_),
    .X(_00176_));
 sky130_fd_sc_hd__nand2_1 _07393_ (.A(_00175_),
    .B(_00176_),
    .Y(_00177_));
 sky130_fd_sc_hd__nand2_1 _07394_ (.A(_06260_),
    .B(net60),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _07395_ (.A(_06272_),
    .B(net61),
    .Y(_00179_));
 sky130_fd_sc_hd__or2_1 _07396_ (.A(_00178_),
    .B(_00179_),
    .X(_00180_));
 sky130_fd_sc_hd__nand2_1 _07397_ (.A(_00178_),
    .B(_00179_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _07398_ (.A(_00180_),
    .B(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__or2_1 _07399_ (.A(_00177_),
    .B(_00182_),
    .X(_00183_));
 sky130_fd_sc_hd__nand2_1 _07400_ (.A(_00182_),
    .B(_00177_),
    .Y(_00184_));
 sky130_fd_sc_hd__nand2_1 _07401_ (.A(_00183_),
    .B(_00184_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_1 _07402_ (.A(_00174_),
    .B(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__inv_2 _07403_ (.A(_00185_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand3_1 _07404_ (.A(_00187_),
    .B(_00172_),
    .C(_00173_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _07405_ (.A(_00186_),
    .B(_00188_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _07406_ (.A(_00159_),
    .B(_00189_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand3_1 _07407_ (.A(_00158_),
    .B(_00186_),
    .C(_00188_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _07408_ (.A(_00190_),
    .B(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__buf_6 _07409_ (.A(_06289_),
    .X(_00193_));
 sky130_fd_sc_hd__nand2_1 _07410_ (.A(_00193_),
    .B(_06204_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _07411_ (.A(_06263_),
    .B(_06213_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _07412_ (.A(net29),
    .B(net58),
    .Y(_00196_));
 sky130_fd_sc_hd__or2_1 _07413_ (.A(_00195_),
    .B(_00196_),
    .X(_00197_));
 sky130_fd_sc_hd__nand2_1 _07414_ (.A(_00195_),
    .B(_00196_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _07415_ (.A(_00197_),
    .B(_00198_),
    .Y(_00199_));
 sky130_fd_sc_hd__or2_1 _07416_ (.A(_00194_),
    .B(_00199_),
    .X(_00200_));
 sky130_fd_sc_hd__nand2_1 _07417_ (.A(_00199_),
    .B(_00194_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _07418_ (.A(_00200_),
    .B(_00201_),
    .Y(_00202_));
 sky130_fd_sc_hd__a21boi_2 _07419_ (.A1(_00114_),
    .A2(_00118_),
    .B1_N(_00117_),
    .Y(_00203_));
 sky130_fd_sc_hd__inv_2 _07420_ (.A(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _07421_ (.A(_00202_),
    .B(_00204_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand3_1 _07422_ (.A(_00200_),
    .B(_00201_),
    .C(_00203_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _07423_ (.A(_00205_),
    .B(_00206_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_1 _07424_ (.A(_00137_),
    .B(_00132_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _07425_ (.A(_00207_),
    .B(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand3b_1 _07426_ (.A_N(_00208_),
    .B(_00205_),
    .C(_00206_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _07427_ (.A(_00209_),
    .B(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _07428_ (.A(_00192_),
    .B(_00211_),
    .Y(_00212_));
 sky130_fd_sc_hd__inv_2 _07429_ (.A(_00211_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand3_1 _07430_ (.A(_00213_),
    .B(_00190_),
    .C(_00191_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _07431_ (.A(_00212_),
    .B(_00214_),
    .Y(_00215_));
 sky130_fd_sc_hd__nor2_1 _07432_ (.A(_00157_),
    .B(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__inv_2 _07433_ (.A(_00216_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _07434_ (.A(_00215_),
    .B(_00157_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _07435_ (.A(_06288_),
    .B(_06209_),
    .Y(_00219_));
 sky130_fd_sc_hd__and2_1 _07436_ (.A(_00143_),
    .B(_00141_),
    .X(_00220_));
 sky130_fd_sc_hd__nor2_1 _07437_ (.A(_00219_),
    .B(_00220_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _07438_ (.A(_00220_),
    .B(_00219_),
    .Y(_00222_));
 sky130_fd_sc_hd__nor2b_1 _07439_ (.A(_00221_),
    .B_N(_00222_),
    .Y(_00223_));
 sky130_fd_sc_hd__a21o_1 _07440_ (.A1(_00217_),
    .A2(_00218_),
    .B1(_00223_),
    .X(_00224_));
 sky130_fd_sc_hd__nand3_1 _07441_ (.A(_00217_),
    .B(_00218_),
    .C(_00223_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand3_2 _07442_ (.A(_00156_),
    .B(_00224_),
    .C(_00225_),
    .Y(_00226_));
 sky130_fd_sc_hd__inv_2 _07443_ (.A(_00156_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _07444_ (.A(_00224_),
    .B(_00225_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _07445_ (.A(_00227_),
    .B(_00228_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _07446_ (.A(_00226_),
    .B(_00229_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _07447_ (.A(_00088_),
    .B(_00083_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _07448_ (.A(_00152_),
    .B(_00154_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _07449_ (.A(_00232_),
    .B(_00077_),
    .Y(_00233_));
 sky130_fd_sc_hd__nand3_1 _07450_ (.A(_00231_),
    .B(_00233_),
    .C(_00155_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _07451_ (.A(_00230_),
    .B(_00234_),
    .Y(_00235_));
 sky130_fd_sc_hd__a21boi_1 _07452_ (.A1(_06443_),
    .A2(_00085_),
    .B1_N(_00083_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _07453_ (.A(_00233_),
    .B(_00155_),
    .Y(_00237_));
 sky130_fd_sc_hd__nor2_1 _07454_ (.A(_00236_),
    .B(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand3_2 _07455_ (.A(_00238_),
    .B(_00226_),
    .C(_00229_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _07456_ (.A(_00235_),
    .B(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _07457_ (.A(_00237_),
    .B(_00236_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand3b_1 _07458_ (.A_N(_00091_),
    .B(_00234_),
    .C(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _07459_ (.A(_00240_),
    .B(_00242_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _07460_ (.A(_00234_),
    .B(_00241_),
    .Y(_00244_));
 sky130_fd_sc_hd__nor2_1 _07461_ (.A(_00091_),
    .B(_00244_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand3_2 _07462_ (.A(_00245_),
    .B(_00235_),
    .C(_00239_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _07463_ (.A(_00243_),
    .B(_00246_),
    .Y(_00247_));
 sky130_fd_sc_hd__inv_2 _07464_ (.A(_00093_),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(_00244_),
    .B(_00091_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand3_1 _07466_ (.A(_00248_),
    .B(_00242_),
    .C(_00249_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _07467_ (.A(_00247_),
    .B(_00250_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _07468_ (.A(_00242_),
    .B(_00249_),
    .Y(_00252_));
 sky130_fd_sc_hd__nor2_1 _07469_ (.A(_00093_),
    .B(_00252_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand3_1 _07470_ (.A(_00253_),
    .B(_00246_),
    .C(_00243_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand2_1 _07471_ (.A(_00252_),
    .B(_00093_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _07472_ (.A(_00255_),
    .B(_00250_),
    .Y(_00256_));
 sky130_fd_sc_hd__nor2_1 _07473_ (.A(_00095_),
    .B(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__a21oi_1 _07474_ (.A1(_00251_),
    .A2(_00254_),
    .B1(_00257_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand3_1 _07475_ (.A(_00257_),
    .B(_00251_),
    .C(_00254_),
    .Y(_00259_));
 sky130_fd_sc_hd__and2b_1 _07476_ (.A_N(_00258_),
    .B(_00259_),
    .X(_00260_));
 sky130_fd_sc_hd__clkbuf_1 _07477_ (.A(_00260_),
    .X(\m1.out[9] ));
 sky130_fd_sc_hd__a21o_1 _07478_ (.A1(_00218_),
    .A2(_00223_),
    .B1(_00216_),
    .X(_00261_));
 sky130_fd_sc_hd__a21oi_1 _07479_ (.A1(_00187_),
    .A2(_00173_),
    .B1(_00171_),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _07480_ (.A(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _07481_ (.A(_06268_),
    .B(net64),
    .Y(_00264_));
 sky130_fd_sc_hd__inv_2 _07482_ (.A(_00264_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _07483_ (.A(net1),
    .B(_06229_),
    .Y(_00266_));
 sky130_fd_sc_hd__inv_2 _07484_ (.A(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__nand2_1 _07485_ (.A(_00265_),
    .B(_00267_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _07486_ (.A(_00264_),
    .B(_00266_),
    .Y(_00269_));
 sky130_fd_sc_hd__clkbuf_8 _07487_ (.A(net63),
    .X(_00270_));
 sky130_fd_sc_hd__nand2_1 _07488_ (.A(_06392_),
    .B(_00270_),
    .Y(_00271_));
 sky130_fd_sc_hd__inv_2 _07489_ (.A(_00271_),
    .Y(_00272_));
 sky130_fd_sc_hd__a21o_1 _07490_ (.A1(_00268_),
    .A2(_00269_),
    .B1(_00272_),
    .X(_00273_));
 sky130_fd_sc_hd__nand3_1 _07491_ (.A(_00268_),
    .B(_00272_),
    .C(_00269_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _07492_ (.A(_00273_),
    .B(_00274_),
    .Y(_00275_));
 sky130_fd_sc_hd__inv_2 _07493_ (.A(_00275_),
    .Y(_00276_));
 sky130_fd_sc_hd__a21oi_2 _07494_ (.A1(_00164_),
    .A2(_00168_),
    .B1(_00163_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _07495_ (.A(_00276_),
    .B(_00277_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand2_1 _07496_ (.A(_00175_),
    .B(_06196_),
    .Y(_00279_));
 sky130_fd_sc_hd__inv_2 _07497_ (.A(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(_06260_),
    .B(_06201_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_1 _07499_ (.A(_06273_),
    .B(_06199_),
    .Y(_00282_));
 sky130_fd_sc_hd__or2_1 _07500_ (.A(_00281_),
    .B(_00282_),
    .X(_00283_));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(_00281_),
    .B(_00282_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _07502_ (.A(_00283_),
    .B(_00284_),
    .Y(_00285_));
 sky130_fd_sc_hd__xor2_2 _07503_ (.A(_00280_),
    .B(_00285_),
    .X(_00286_));
 sky130_fd_sc_hd__inv_2 _07504_ (.A(_00277_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _07505_ (.A(_00275_),
    .B(_00287_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand3_1 _07506_ (.A(_00278_),
    .B(_00286_),
    .C(_00288_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _07507_ (.A(_00276_),
    .B(_00287_),
    .Y(_00290_));
 sky130_fd_sc_hd__inv_2 _07508_ (.A(_00286_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _07509_ (.A(_00275_),
    .B(_00277_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand3_1 _07510_ (.A(_00290_),
    .B(_00291_),
    .C(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand3_1 _07511_ (.A(_00263_),
    .B(_00289_),
    .C(_00293_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _07512_ (.A(_00293_),
    .B(_00289_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _07513_ (.A(_00295_),
    .B(_00262_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _07514_ (.A(_00294_),
    .B(_00296_),
    .Y(_00297_));
 sky130_fd_sc_hd__inv_2 _07515_ (.A(_06197_),
    .Y(_00298_));
 sky130_fd_sc_hd__buf_6 _07516_ (.A(_06263_),
    .X(_00299_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_00299_),
    .B(_06210_),
    .Y(_00300_));
 sky130_fd_sc_hd__or3_1 _07518_ (.A(_00069_),
    .B(_00298_),
    .C(_00300_),
    .X(_00301_));
 sky130_fd_sc_hd__o21ai_1 _07519_ (.A1(_00069_),
    .A2(_00298_),
    .B1(_00300_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _07520_ (.A(_00301_),
    .B(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _07521_ (.A(_00193_),
    .B(_06214_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _07522_ (.A(_00303_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__inv_2 _07523_ (.A(_00304_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand3_2 _07524_ (.A(_00301_),
    .B(_00306_),
    .C(_00302_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _07525_ (.A(_00305_),
    .B(_00307_),
    .Y(_00308_));
 sky130_fd_sc_hd__o21a_1 _07526_ (.A1(_00177_),
    .A2(_00182_),
    .B1(_00180_),
    .X(_00309_));
 sky130_fd_sc_hd__nand2_1 _07527_ (.A(_00308_),
    .B(_00309_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _07528_ (.A(_00183_),
    .B(_00180_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand3_1 _07529_ (.A(_00311_),
    .B(_00305_),
    .C(_00307_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _07530_ (.A(_00200_),
    .B(_00197_),
    .Y(_00313_));
 sky130_fd_sc_hd__nand3_1 _07531_ (.A(_00310_),
    .B(_00312_),
    .C(_00313_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _07532_ (.A(_00308_),
    .B(_00311_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand3_1 _07533_ (.A(_00305_),
    .B(_00309_),
    .C(_00307_),
    .Y(_00316_));
 sky130_fd_sc_hd__inv_2 _07534_ (.A(_00313_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand3_1 _07535_ (.A(_00315_),
    .B(_00316_),
    .C(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__nand2_1 _07536_ (.A(_00314_),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _07537_ (.A(_00297_),
    .B(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__inv_2 _07538_ (.A(_00319_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand3_1 _07539_ (.A(_00294_),
    .B(_00321_),
    .C(_00296_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _07540_ (.A(_00320_),
    .B(_00322_),
    .Y(_00323_));
 sky130_fd_sc_hd__a21boi_1 _07541_ (.A1(_00213_),
    .A2(_00190_),
    .B1_N(_00191_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _07542_ (.A(_00323_),
    .B(_00324_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _07543_ (.A(_00214_),
    .B(_00191_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand3_2 _07544_ (.A(_00326_),
    .B(_00320_),
    .C(_00322_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _07545_ (.A(_00325_),
    .B(_00327_),
    .Y(_00328_));
 sky130_fd_sc_hd__inv_2 _07546_ (.A(_06287_),
    .Y(_00329_));
 sky130_fd_sc_hd__inv_2 _07547_ (.A(net2),
    .Y(_00330_));
 sky130_fd_sc_hd__inv_2 _07548_ (.A(_06207_),
    .Y(_00331_));
 sky130_fd_sc_hd__or4_2 _07549_ (.A(_00329_),
    .B(_00330_),
    .C(_06330_),
    .D(_00331_),
    .X(_00332_));
 sky130_fd_sc_hd__a22o_1 _07550_ (.A1(_06288_),
    .A2(_06206_),
    .B1(_06292_),
    .B2(_06208_),
    .X(_00333_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(_00332_),
    .B(_00333_),
    .Y(_00334_));
 sky130_fd_sc_hd__o21a_1 _07552_ (.A1(_00202_),
    .A2(_00203_),
    .B1(_00209_),
    .X(_00335_));
 sky130_fd_sc_hd__nor2_1 _07553_ (.A(_00334_),
    .B(_00335_),
    .Y(_00336_));
 sky130_fd_sc_hd__inv_2 _07554_ (.A(_00336_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _07555_ (.A(_00335_),
    .B(_00334_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _07556_ (.A(_00337_),
    .B(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _07557_ (.A(_00328_),
    .B(_00339_),
    .Y(_00340_));
 sky130_fd_sc_hd__inv_2 _07558_ (.A(_00339_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand3_2 _07559_ (.A(_00325_),
    .B(_00327_),
    .C(_00341_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand3_2 _07560_ (.A(_00261_),
    .B(_00340_),
    .C(_00342_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _07561_ (.A(_00340_),
    .B(_00342_),
    .Y(_00344_));
 sky130_fd_sc_hd__a21oi_1 _07562_ (.A1(_00218_),
    .A2(_00223_),
    .B1(_00216_),
    .Y(_00345_));
 sky130_fd_sc_hd__nand2_1 _07563_ (.A(_00344_),
    .B(_00345_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _07564_ (.A(_00343_),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_2 _07565_ (.A(_00221_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _07566_ (.A(_00347_),
    .B(_00348_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand3_1 _07567_ (.A(_00343_),
    .B(_00346_),
    .C(_00221_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _07568_ (.A(_00349_),
    .B(_00350_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _07569_ (.A(_00351_),
    .B(_00226_),
    .Y(_00352_));
 sky130_fd_sc_hd__inv_2 _07570_ (.A(_00226_),
    .Y(_00353_));
 sky130_fd_sc_hd__nand3_2 _07571_ (.A(_00349_),
    .B(_00353_),
    .C(_00350_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _07572_ (.A(_00352_),
    .B(_00354_),
    .Y(_00355_));
 sky130_fd_sc_hd__nand2_1 _07573_ (.A(_00355_),
    .B(_00239_),
    .Y(_00356_));
 sky130_fd_sc_hd__inv_2 _07574_ (.A(_00239_),
    .Y(_00357_));
 sky130_fd_sc_hd__nand3_2 _07575_ (.A(_00352_),
    .B(_00357_),
    .C(_00354_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand2_1 _07576_ (.A(_00356_),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_1 _07577_ (.A(_00359_),
    .B(_00246_),
    .Y(_00360_));
 sky130_fd_sc_hd__inv_2 _07578_ (.A(_00246_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand3_1 _07579_ (.A(_00361_),
    .B(_00356_),
    .C(_00358_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_1 _07580_ (.A(_00360_),
    .B(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__nand2_1 _07581_ (.A(_00259_),
    .B(_00254_),
    .Y(_00364_));
 sky130_fd_sc_hd__inv_2 _07582_ (.A(_00364_),
    .Y(_00365_));
 sky130_fd_sc_hd__or2_1 _07583_ (.A(_00363_),
    .B(_00365_),
    .X(_00366_));
 sky130_fd_sc_hd__nand2_1 _07584_ (.A(_00365_),
    .B(_00363_),
    .Y(_00367_));
 sky130_fd_sc_hd__and2_1 _07585_ (.A(_00366_),
    .B(_00367_),
    .X(_00368_));
 sky130_fd_sc_hd__clkbuf_1 _07586_ (.A(_00368_),
    .X(\m1.out[10] ));
 sky130_fd_sc_hd__nand2_1 _07587_ (.A(_00350_),
    .B(_00343_),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _07588_ (.A(_00342_),
    .B(_00327_),
    .Y(_00370_));
 sky130_fd_sc_hd__inv_2 _07589_ (.A(_00296_),
    .Y(_00371_));
 sky130_fd_sc_hd__o21ai_1 _07590_ (.A1(_00319_),
    .A2(_00371_),
    .B1(_00294_),
    .Y(_00372_));
 sky130_fd_sc_hd__inv_2 _07591_ (.A(_00372_),
    .Y(_00373_));
 sky130_fd_sc_hd__nand2_1 _07592_ (.A(_00293_),
    .B(_00290_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _07593_ (.A(_06327_),
    .B(_06230_),
    .Y(_00375_));
 sky130_fd_sc_hd__buf_8 _07594_ (.A(_06227_),
    .X(_00376_));
 sky130_fd_sc_hd__nand2_1 _07595_ (.A(_06270_),
    .B(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__nor2_1 _07596_ (.A(_00375_),
    .B(_00377_),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_2 _07597_ (.A(_00378_),
    .Y(_00379_));
 sky130_fd_sc_hd__nand2_1 _07598_ (.A(_00375_),
    .B(_00377_),
    .Y(_00380_));
 sky130_fd_sc_hd__nand2_1 _07599_ (.A(_06276_),
    .B(_06225_),
    .Y(_00381_));
 sky130_fd_sc_hd__inv_4 _07600_ (.A(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__a21o_1 _07601_ (.A1(_00379_),
    .A2(_00380_),
    .B1(_00382_),
    .X(_00383_));
 sky130_fd_sc_hd__nand3_1 _07602_ (.A(_00379_),
    .B(_00382_),
    .C(_00380_),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_1 _07603_ (.A(_00383_),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _07604_ (.A(_00274_),
    .B(_00268_),
    .Y(_00386_));
 sky130_fd_sc_hd__clkinvlp_2 _07605_ (.A(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _07606_ (.A(_00385_),
    .B(_00387_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand3_1 _07607_ (.A(_00383_),
    .B(_00386_),
    .C(_00384_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _07608_ (.A(_00388_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _07609_ (.A(_06260_),
    .B(net62),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_1 _07610_ (.A(_06272_),
    .B(net63),
    .Y(_00392_));
 sky130_fd_sc_hd__nor2_1 _07611_ (.A(_00391_),
    .B(_00392_),
    .Y(_00393_));
 sky130_fd_sc_hd__inv_2 _07612_ (.A(_00393_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _07613_ (.A(_00391_),
    .B(_00392_),
    .Y(_00395_));
 sky130_fd_sc_hd__nand2_1 _07614_ (.A(_06258_),
    .B(_06201_),
    .Y(_00396_));
 sky130_fd_sc_hd__inv_2 _07615_ (.A(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__a21o_1 _07616_ (.A1(_00394_),
    .A2(_00395_),
    .B1(_00397_),
    .X(_00398_));
 sky130_fd_sc_hd__nand3_1 _07617_ (.A(_00394_),
    .B(_00397_),
    .C(_00395_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _07618_ (.A(_00398_),
    .B(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _07619_ (.A(_00390_),
    .B(_00400_),
    .Y(_00401_));
 sky130_fd_sc_hd__inv_2 _07620_ (.A(_00400_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand3_1 _07621_ (.A(_00388_),
    .B(_00402_),
    .C(_00389_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand3_1 _07622_ (.A(_00374_),
    .B(_00401_),
    .C(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__a21boi_1 _07623_ (.A1(_00291_),
    .A2(_00292_),
    .B1_N(_00290_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _07624_ (.A(_00401_),
    .B(_00403_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _07625_ (.A(_00405_),
    .B(_00406_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand2_1 _07626_ (.A(_00404_),
    .B(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__nand2_1 _07627_ (.A(_06263_),
    .B(_06197_),
    .Y(_00409_));
 sky130_fd_sc_hd__inv_2 _07628_ (.A(_00409_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _07629_ (.A(net29),
    .B(net60),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _07630_ (.A(_00411_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _07631_ (.A(_00410_),
    .B(_00412_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _07632_ (.A(_00409_),
    .B(_00411_),
    .Y(_00414_));
 sky130_fd_sc_hd__nand2_1 _07633_ (.A(_06289_),
    .B(_06210_),
    .Y(_00415_));
 sky130_fd_sc_hd__inv_2 _07634_ (.A(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__a21o_1 _07635_ (.A1(_00413_),
    .A2(_00414_),
    .B1(_00416_),
    .X(_00417_));
 sky130_fd_sc_hd__nand3_1 _07636_ (.A(_00413_),
    .B(_00416_),
    .C(_00414_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _07637_ (.A(_00417_),
    .B(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__inv_2 _07638_ (.A(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__a21boi_1 _07639_ (.A1(_00280_),
    .A2(_00284_),
    .B1_N(_00283_),
    .Y(_00421_));
 sky130_fd_sc_hd__inv_2 _07640_ (.A(_00421_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _07641_ (.A(_00420_),
    .B(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _07642_ (.A(_00419_),
    .B(_00421_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _07643_ (.A(_00423_),
    .B(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _07644_ (.A(_00307_),
    .B(_00301_),
    .Y(_00426_));
 sky130_fd_sc_hd__inv_2 _07645_ (.A(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _07646_ (.A(_00425_),
    .B(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand3_1 _07647_ (.A(_00423_),
    .B(_00426_),
    .C(_00424_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _07648_ (.A(_00428_),
    .B(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _07649_ (.A(_00408_),
    .B(_00430_),
    .Y(_00431_));
 sky130_fd_sc_hd__inv_2 _07650_ (.A(_00430_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand3_1 _07651_ (.A(_00404_),
    .B(_00432_),
    .C(_00407_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _07652_ (.A(_00431_),
    .B(_00433_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _07653_ (.A(_00373_),
    .B(_00434_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand3_1 _07654_ (.A(_00372_),
    .B(_00431_),
    .C(_00433_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _07655_ (.A(_00435_),
    .B(_00436_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _07656_ (.A(_06291_),
    .B(_06207_),
    .Y(_00438_));
 sky130_fd_sc_hd__buf_4 _07657_ (.A(net2),
    .X(_00439_));
 sky130_fd_sc_hd__nand2_1 _07658_ (.A(_00439_),
    .B(_06204_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _07659_ (.A(_06287_),
    .B(_06214_),
    .Y(_00441_));
 sky130_fd_sc_hd__nor2_1 _07660_ (.A(_00440_),
    .B(_00441_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _07661_ (.A(_00440_),
    .B(_00441_),
    .Y(_00443_));
 sky130_fd_sc_hd__and2b_1 _07662_ (.A_N(_00442_),
    .B(_00443_),
    .X(_00444_));
 sky130_fd_sc_hd__xor2_1 _07663_ (.A(_00438_),
    .B(_00444_),
    .X(_00445_));
 sky130_fd_sc_hd__nor2_1 _07664_ (.A(_00445_),
    .B(_00332_),
    .Y(_00446_));
 sky130_fd_sc_hd__inv_2 _07665_ (.A(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand2_1 _07666_ (.A(_00332_),
    .B(_00445_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _07667_ (.A(_00447_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__and2_1 _07668_ (.A(_00314_),
    .B(_00312_),
    .X(_00450_));
 sky130_fd_sc_hd__nor2_1 _07669_ (.A(_00449_),
    .B(_00450_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _07670_ (.A(_00450_),
    .B(_00449_),
    .Y(_00452_));
 sky130_fd_sc_hd__and2b_1 _07671_ (.A_N(_00451_),
    .B(_00452_),
    .X(_00453_));
 sky130_fd_sc_hd__inv_2 _07672_ (.A(_00453_),
    .Y(_00454_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(_00437_),
    .B(_00454_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand3_1 _07674_ (.A(_00435_),
    .B(_00436_),
    .C(_00453_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand3_1 _07675_ (.A(_00370_),
    .B(_00455_),
    .C(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _07676_ (.A(_00455_),
    .B(_00456_),
    .Y(_00458_));
 sky130_fd_sc_hd__a21boi_1 _07677_ (.A1(_00341_),
    .A2(_00325_),
    .B1_N(_00327_),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _07678_ (.A(_00458_),
    .B(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand3_1 _07679_ (.A(_00457_),
    .B(_00336_),
    .C(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _07680_ (.A(_00457_),
    .B(_00460_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _07681_ (.A(_00462_),
    .B(_00337_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand3_2 _07682_ (.A(_00369_),
    .B(_00461_),
    .C(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _07683_ (.A(_00463_),
    .B(_00461_),
    .Y(_00465_));
 sky130_fd_sc_hd__a21boi_1 _07684_ (.A1(_00221_),
    .A2(_00346_),
    .B1_N(_00343_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _07685_ (.A(_00465_),
    .B(_00466_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _07686_ (.A(_00464_),
    .B(_00467_),
    .Y(_00468_));
 sky130_fd_sc_hd__nand2_1 _07687_ (.A(_00468_),
    .B(_00354_),
    .Y(_00469_));
 sky130_fd_sc_hd__inv_2 _07688_ (.A(_00354_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand3_4 _07689_ (.A(_00470_),
    .B(_00464_),
    .C(_00467_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _07690_ (.A(_00469_),
    .B(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__nand2_1 _07691_ (.A(_00472_),
    .B(_00358_),
    .Y(_00473_));
 sky130_fd_sc_hd__inv_2 _07692_ (.A(_00358_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand3_1 _07693_ (.A(_00474_),
    .B(_00469_),
    .C(_00471_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(_00473_),
    .B(_00475_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _07695_ (.A(_00366_),
    .B(_00362_),
    .Y(_00477_));
 sky130_fd_sc_hd__or2_1 _07696_ (.A(_00476_),
    .B(_00477_),
    .X(_00478_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(_00477_),
    .B(_00476_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _07698_ (.A(_00478_),
    .B(_00479_),
    .Y(\m1.out[11] ));
 sky130_fd_sc_hd__nor2_1 _07699_ (.A(_00363_),
    .B(_00476_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand2_1 _07700_ (.A(_00480_),
    .B(_00364_),
    .Y(_00481_));
 sky130_fd_sc_hd__inv_2 _07701_ (.A(_00362_),
    .Y(_00482_));
 sky130_fd_sc_hd__a21boi_1 _07702_ (.A1(_00482_),
    .A2(_00473_),
    .B1_N(_00475_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _07703_ (.A(_00481_),
    .B(_00483_),
    .Y(_00484_));
 sky130_fd_sc_hd__inv_2 _07704_ (.A(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__inv_2 _07705_ (.A(_00471_),
    .Y(_00486_));
 sky130_fd_sc_hd__nor2_1 _07706_ (.A(_00466_),
    .B(_00465_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_1 _07707_ (.A(_00459_),
    .B(_00458_),
    .Y(_00488_));
 sky130_fd_sc_hd__a21o_1 _07708_ (.A1(_00460_),
    .A2(_00336_),
    .B1(_00488_),
    .X(_00489_));
 sky130_fd_sc_hd__nor2_1 _07709_ (.A(_00434_),
    .B(_00373_),
    .Y(_00490_));
 sky130_fd_sc_hd__a21oi_1 _07710_ (.A1(_00435_),
    .A2(_00453_),
    .B1(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_1 _07711_ (.A(_06268_),
    .B(_00376_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _07712_ (.A(_06270_),
    .B(_06219_),
    .Y(_00493_));
 sky130_fd_sc_hd__nor2_1 _07713_ (.A(_00492_),
    .B(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _07714_ (.A(_00492_),
    .B(_00493_),
    .Y(_00495_));
 sky130_fd_sc_hd__inv_2 _07715_ (.A(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _07716_ (.A(_06275_),
    .B(_06229_),
    .Y(_00497_));
 sky130_fd_sc_hd__o21ai_1 _07717_ (.A1(_00494_),
    .A2(_00496_),
    .B1(_00497_),
    .Y(_00498_));
 sky130_fd_sc_hd__inv_2 _07718_ (.A(_00497_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand3b_1 _07719_ (.A_N(_00494_),
    .B(_00499_),
    .C(_00495_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _07720_ (.A(_00498_),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__inv_2 _07721_ (.A(_00501_),
    .Y(_00502_));
 sky130_fd_sc_hd__a21oi_2 _07722_ (.A1(_00380_),
    .A2(_00382_),
    .B1(_00378_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _07723_ (.A(_00502_),
    .B(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _07724_ (.A(_06261_),
    .B(_00270_),
    .Y(_00505_));
 sky130_fd_sc_hd__nand2_1 _07725_ (.A(_06273_),
    .B(net64),
    .Y(_00506_));
 sky130_fd_sc_hd__nor2_1 _07726_ (.A(_00505_),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(_00505_),
    .B(_00506_),
    .Y(_00508_));
 sky130_fd_sc_hd__inv_2 _07728_ (.A(_00508_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _07729_ (.A(_06258_),
    .B(_06199_),
    .Y(_00510_));
 sky130_fd_sc_hd__o21ai_1 _07730_ (.A1(_00507_),
    .A2(_00509_),
    .B1(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__inv_2 _07731_ (.A(_00510_),
    .Y(_00512_));
 sky130_fd_sc_hd__nand3b_1 _07732_ (.A_N(_00507_),
    .B(_00512_),
    .C(_00508_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _07733_ (.A(_00511_),
    .B(_00513_),
    .Y(_00514_));
 sky130_fd_sc_hd__inv_2 _07734_ (.A(_00503_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _07735_ (.A(_00501_),
    .B(_00515_),
    .Y(_00516_));
 sky130_fd_sc_hd__nand3_1 _07736_ (.A(_00504_),
    .B(_00514_),
    .C(_00516_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _07737_ (.A(_00502_),
    .B(_00515_),
    .Y(_00518_));
 sky130_fd_sc_hd__inv_2 _07738_ (.A(_00514_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _07739_ (.A(_00501_),
    .B(_00503_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand3_1 _07740_ (.A(_00518_),
    .B(_00519_),
    .C(_00520_),
    .Y(_00521_));
 sky130_fd_sc_hd__nand2_1 _07741_ (.A(_00517_),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__a21boi_2 _07742_ (.A1(_00388_),
    .A2(_00402_),
    .B1_N(_00389_),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2b_1 _07743_ (.A_N(_00522_),
    .B(_00523_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _07744_ (.A(_00399_),
    .B(_00394_),
    .Y(_00525_));
 sky130_fd_sc_hd__inv_2 _07745_ (.A(_00525_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _07746_ (.A(_00299_),
    .B(_06195_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_06265_),
    .B(_06201_),
    .Y(_00528_));
 sky130_fd_sc_hd__nor2_1 _07748_ (.A(_00527_),
    .B(_00528_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _07749_ (.A(_00527_),
    .B(_00528_),
    .Y(_00530_));
 sky130_fd_sc_hd__inv_2 _07750_ (.A(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _07751_ (.A(_06289_),
    .B(_00176_),
    .Y(_00532_));
 sky130_fd_sc_hd__o21ai_1 _07752_ (.A1(_00529_),
    .A2(_00531_),
    .B1(_00532_),
    .Y(_00533_));
 sky130_fd_sc_hd__inv_2 _07753_ (.A(_00532_),
    .Y(_00534_));
 sky130_fd_sc_hd__nand3b_1 _07754_ (.A_N(_00529_),
    .B(_00534_),
    .C(_00530_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _07755_ (.A(_00533_),
    .B(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _07756_ (.A(_00526_),
    .B(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__nand3_1 _07757_ (.A(_00525_),
    .B(_00533_),
    .C(_00535_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _07758_ (.A(_00537_),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand3_1 _07759_ (.A(_00539_),
    .B(_00413_),
    .C(_00418_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _07760_ (.A(_00418_),
    .B(_00413_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand3_1 _07761_ (.A(_00537_),
    .B(_00538_),
    .C(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _07762_ (.A(_00540_),
    .B(_00542_),
    .Y(_00543_));
 sky130_fd_sc_hd__inv_2 _07763_ (.A(_00523_),
    .Y(_00544_));
 sky130_fd_sc_hd__nand2_1 _07764_ (.A(_00544_),
    .B(_00522_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand3_1 _07765_ (.A(_00524_),
    .B(_00543_),
    .C(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__nor2_1 _07766_ (.A(_00523_),
    .B(_00522_),
    .Y(_00547_));
 sky130_fd_sc_hd__inv_2 _07767_ (.A(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__inv_2 _07768_ (.A(_00543_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _07769_ (.A(_00522_),
    .B(_00523_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand3_1 _07770_ (.A(_00548_),
    .B(_00549_),
    .C(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _07771_ (.A(_00546_),
    .B(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__nor2_1 _07772_ (.A(_00406_),
    .B(_00405_),
    .Y(_00553_));
 sky130_fd_sc_hd__a21oi_2 _07773_ (.A1(_00407_),
    .A2(_00432_),
    .B1(_00553_),
    .Y(_00554_));
 sky130_fd_sc_hd__inv_2 _07774_ (.A(_00554_),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _07775_ (.A(_00552_),
    .B(_00555_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand3_1 _07776_ (.A(_00554_),
    .B(_00546_),
    .C(_00551_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _07777_ (.A(_00556_),
    .B(_00557_),
    .Y(_00558_));
 sky130_fd_sc_hd__inv_2 _07778_ (.A(_00438_),
    .Y(_00559_));
 sky130_fd_sc_hd__a21oi_2 _07779_ (.A1(_00443_),
    .A2(_00559_),
    .B1(_00442_),
    .Y(_00560_));
 sky130_fd_sc_hd__clkbuf_8 _07780_ (.A(net3),
    .X(_00561_));
 sky130_fd_sc_hd__nand2_1 _07781_ (.A(_00561_),
    .B(_06204_),
    .Y(_00562_));
 sky130_fd_sc_hd__inv_2 _07782_ (.A(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand2_1 _07783_ (.A(_00439_),
    .B(_06214_),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_1 _07784_ (.A(_06287_),
    .B(_06211_),
    .Y(_00565_));
 sky130_fd_sc_hd__xor2_1 _07785_ (.A(_00564_),
    .B(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__or2_1 _07786_ (.A(_00563_),
    .B(_00566_),
    .X(_00567_));
 sky130_fd_sc_hd__nand2_1 _07787_ (.A(_00566_),
    .B(_00563_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _07788_ (.A(_00567_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__nor2_1 _07789_ (.A(_00560_),
    .B(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__inv_2 _07790_ (.A(_00570_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _07791_ (.A(_06280_),
    .B(_06208_),
    .Y(_00572_));
 sky130_fd_sc_hd__inv_2 _07792_ (.A(_00572_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _07793_ (.A(_00569_),
    .B(_00560_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand3_1 _07794_ (.A(_00571_),
    .B(_00573_),
    .C(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__a21o_1 _07795_ (.A1(_00567_),
    .A2(_00568_),
    .B1(_00560_),
    .X(_00576_));
 sky130_fd_sc_hd__nand3_1 _07796_ (.A(_00567_),
    .B(_00560_),
    .C(_00568_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand3_1 _07797_ (.A(_00576_),
    .B(_00577_),
    .C(_00572_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _07798_ (.A(_00575_),
    .B(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(_00429_),
    .B(_00423_),
    .Y(_00580_));
 sky130_fd_sc_hd__inv_2 _07800_ (.A(_00580_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_1 _07801_ (.A(_00579_),
    .B(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand3_1 _07802_ (.A(_00575_),
    .B(_00578_),
    .C(_00580_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(_00582_),
    .B(_00583_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _07804_ (.A(_00584_),
    .B(_00447_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand3_1 _07805_ (.A(_00582_),
    .B(_00583_),
    .C(_00446_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _07806_ (.A(_00585_),
    .B(_00586_),
    .Y(_00587_));
 sky130_fd_sc_hd__inv_2 _07807_ (.A(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _07808_ (.A(_00558_),
    .B(_00588_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand3_1 _07809_ (.A(_00587_),
    .B(_00556_),
    .C(_00557_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _07810_ (.A(_00589_),
    .B(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hd__nor2_1 _07811_ (.A(_00491_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__inv_2 _07812_ (.A(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _07813_ (.A(_00591_),
    .B(_00491_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand3_1 _07814_ (.A(_00593_),
    .B(_00451_),
    .C(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(_00593_),
    .B(_00594_),
    .Y(_00596_));
 sky130_fd_sc_hd__inv_2 _07816_ (.A(_00451_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _07817_ (.A(_00596_),
    .B(_00597_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand3_2 _07818_ (.A(_00489_),
    .B(_00595_),
    .C(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _07819_ (.A(_00598_),
    .B(_00595_),
    .Y(_00600_));
 sky130_fd_sc_hd__a21oi_1 _07820_ (.A1(_00460_),
    .A2(_00336_),
    .B1(_00488_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _07821_ (.A(_00600_),
    .B(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand3_1 _07822_ (.A(_00487_),
    .B(_00599_),
    .C(_00602_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _07823_ (.A(_00599_),
    .B(_00602_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _07824_ (.A(_00604_),
    .B(_00464_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand3_1 _07825_ (.A(_00486_),
    .B(_00603_),
    .C(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _07826_ (.A(_00605_),
    .B(_00603_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _07827_ (.A(_00607_),
    .B(_00471_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _07828_ (.A(_00606_),
    .B(_00608_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _07829_ (.A(_00485_),
    .B(_00609_),
    .Y(_00610_));
 sky130_fd_sc_hd__inv_2 _07830_ (.A(_00609_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _07831_ (.A(_00484_),
    .B(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__and2_1 _07832_ (.A(_00610_),
    .B(_00612_),
    .X(_00613_));
 sky130_fd_sc_hd__clkbuf_1 _07833_ (.A(_00613_),
    .X(\m1.out[12] ));
 sky130_fd_sc_hd__nor2_1 _07834_ (.A(_00464_),
    .B(_00604_),
    .Y(_00614_));
 sky130_fd_sc_hd__nor2_1 _07835_ (.A(_00601_),
    .B(_00600_),
    .Y(_00615_));
 sky130_fd_sc_hd__a21oi_2 _07836_ (.A1(_00549_),
    .A2(_00550_),
    .B1(_00547_),
    .Y(_00616_));
 sky130_fd_sc_hd__nor2_1 _07837_ (.A(_00503_),
    .B(_00501_),
    .Y(_00617_));
 sky130_fd_sc_hd__a21oi_2 _07838_ (.A1(_00520_),
    .A2(_00519_),
    .B1(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__nand2_1 _07839_ (.A(_06268_),
    .B(_06219_),
    .Y(_00619_));
 sky130_fd_sc_hd__inv_2 _07840_ (.A(_00619_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _07841_ (.A(net1),
    .B(_06217_),
    .Y(_00621_));
 sky130_fd_sc_hd__inv_2 _07842_ (.A(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _07843_ (.A(_00620_),
    .B(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _07844_ (.A(_00619_),
    .B(_00621_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _07845_ (.A(_00623_),
    .B(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _07846_ (.A(_06275_),
    .B(_06227_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _07847_ (.A(_00625_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__inv_2 _07848_ (.A(_00626_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand3_1 _07849_ (.A(_00623_),
    .B(_00628_),
    .C(_00624_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _07850_ (.A(_00627_),
    .B(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hd__a21oi_2 _07851_ (.A1(_00495_),
    .A2(_00499_),
    .B1(_00494_),
    .Y(_00631_));
 sky130_fd_sc_hd__inv_2 _07852_ (.A(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _07853_ (.A(_00630_),
    .B(_00632_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand3_1 _07854_ (.A(_00627_),
    .B(_00631_),
    .C(_00629_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _07855_ (.A(_00633_),
    .B(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _07856_ (.A(_06260_),
    .B(net64),
    .Y(_00636_));
 sky130_fd_sc_hd__inv_2 _07857_ (.A(_00636_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _07858_ (.A(_06272_),
    .B(_06229_),
    .Y(_00638_));
 sky130_fd_sc_hd__inv_2 _07859_ (.A(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand2_1 _07860_ (.A(_00637_),
    .B(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _07861_ (.A(_00636_),
    .B(_00638_),
    .Y(_00641_));
 sky130_fd_sc_hd__nand2_1 _07862_ (.A(_00640_),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__nand2_1 _07863_ (.A(_00175_),
    .B(_00270_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _07864_ (.A(_00642_),
    .B(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__inv_2 _07865_ (.A(_00643_),
    .Y(_00645_));
 sky130_fd_sc_hd__nand3_1 _07866_ (.A(_00640_),
    .B(_00645_),
    .C(_00641_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand2_1 _07867_ (.A(_00644_),
    .B(_00646_),
    .Y(_00647_));
 sky130_fd_sc_hd__inv_2 _07868_ (.A(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__nand2_1 _07869_ (.A(_00635_),
    .B(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__nand3_1 _07870_ (.A(_00633_),
    .B(_00634_),
    .C(_00647_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand2_1 _07871_ (.A(_00649_),
    .B(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hd__nand2b_1 _07872_ (.A_N(_00618_),
    .B(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__nand3_1 _07873_ (.A(_00618_),
    .B(_00650_),
    .C(_00649_),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _07874_ (.A(_00652_),
    .B(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _07875_ (.A(_06263_),
    .B(net61),
    .Y(_00655_));
 sky130_fd_sc_hd__inv_2 _07876_ (.A(_00655_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand2_1 _07877_ (.A(net29),
    .B(net62),
    .Y(_00657_));
 sky130_fd_sc_hd__inv_2 _07878_ (.A(_00657_),
    .Y(_00658_));
 sky130_fd_sc_hd__nand2_1 _07879_ (.A(_00656_),
    .B(_00658_),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_1 _07880_ (.A(_00655_),
    .B(_00657_),
    .Y(_00660_));
 sky130_fd_sc_hd__nand2_1 _07881_ (.A(_00659_),
    .B(_00660_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand2_1 _07882_ (.A(_00193_),
    .B(_06196_),
    .Y(_00662_));
 sky130_fd_sc_hd__nand2_1 _07883_ (.A(_00661_),
    .B(_00662_),
    .Y(_00663_));
 sky130_fd_sc_hd__nand3b_1 _07884_ (.A_N(_00662_),
    .B(_00659_),
    .C(_00660_),
    .Y(_00664_));
 sky130_fd_sc_hd__nand2_1 _07885_ (.A(_00663_),
    .B(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__a21oi_1 _07886_ (.A1(_00508_),
    .A2(_00512_),
    .B1(_00507_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand2_1 _07887_ (.A(_00665_),
    .B(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__a21o_1 _07888_ (.A1(_00508_),
    .A2(_00512_),
    .B1(_00507_),
    .X(_00668_));
 sky130_fd_sc_hd__nand3_1 _07889_ (.A(_00668_),
    .B(_00664_),
    .C(_00663_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand2_1 _07890_ (.A(_00667_),
    .B(_00669_),
    .Y(_00670_));
 sky130_fd_sc_hd__a21oi_1 _07891_ (.A1(_00530_),
    .A2(_00534_),
    .B1(_00529_),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _07892_ (.A(_00670_),
    .B(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__inv_2 _07893_ (.A(_00671_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand3_1 _07894_ (.A(_00667_),
    .B(_00669_),
    .C(_00673_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _07895_ (.A(_00672_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__inv_2 _07896_ (.A(_00675_),
    .Y(_00676_));
 sky130_fd_sc_hd__nand2_1 _07897_ (.A(_00654_),
    .B(_00676_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand3_1 _07898_ (.A(_00652_),
    .B(_00675_),
    .C(_00653_),
    .Y(_00678_));
 sky130_fd_sc_hd__nand2_1 _07899_ (.A(_00677_),
    .B(_00678_),
    .Y(_00679_));
 sky130_fd_sc_hd__nor2_1 _07900_ (.A(_00616_),
    .B(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__nor2_1 _07901_ (.A(_00536_),
    .B(_00526_),
    .Y(_00681_));
 sky130_fd_sc_hd__a21oi_2 _07902_ (.A1(_00537_),
    .A2(_00541_),
    .B1(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__inv_2 _07903_ (.A(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__nand2_1 _07904_ (.A(_00439_),
    .B(_06210_),
    .Y(_00684_));
 sky130_fd_sc_hd__nand2_1 _07905_ (.A(_06287_),
    .B(_00176_),
    .Y(_00685_));
 sky130_fd_sc_hd__nor2_1 _07906_ (.A(_00684_),
    .B(_00685_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand2_1 _07907_ (.A(_00684_),
    .B(_00685_),
    .Y(_00687_));
 sky130_fd_sc_hd__inv_2 _07908_ (.A(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand2_1 _07909_ (.A(_06291_),
    .B(_06214_),
    .Y(_00689_));
 sky130_fd_sc_hd__o21ai_1 _07910_ (.A1(_00686_),
    .A2(_00688_),
    .B1(_00689_),
    .Y(_00690_));
 sky130_fd_sc_hd__inv_2 _07911_ (.A(_00689_),
    .Y(_00691_));
 sky130_fd_sc_hd__nand3b_1 _07912_ (.A_N(_00686_),
    .B(_00691_),
    .C(_00687_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand2_1 _07913_ (.A(_00690_),
    .B(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__nand2_1 _07914_ (.A(_00564_),
    .B(_00565_),
    .Y(_00694_));
 sky130_fd_sc_hd__nor2_1 _07915_ (.A(_00564_),
    .B(_00565_),
    .Y(_00695_));
 sky130_fd_sc_hd__a21oi_1 _07916_ (.A1(_00694_),
    .A2(_00563_),
    .B1(_00695_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_1 _07917_ (.A(_00693_),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand3b_1 _07918_ (.A_N(_00696_),
    .B(_00690_),
    .C(_00692_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand2_1 _07919_ (.A(_00697_),
    .B(_00698_),
    .Y(_00699_));
 sky130_fd_sc_hd__inv_2 _07920_ (.A(net4),
    .Y(_00700_));
 sky130_fd_sc_hd__buf_6 _07921_ (.A(_06278_),
    .X(_00701_));
 sky130_fd_sc_hd__nand2_1 _07922_ (.A(_00701_),
    .B(_06207_),
    .Y(_00702_));
 sky130_fd_sc_hd__nor3_1 _07923_ (.A(_00700_),
    .B(_06330_),
    .C(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__inv_2 _07924_ (.A(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__o21ai_1 _07925_ (.A1(_00700_),
    .A2(_06330_),
    .B1(_00702_),
    .Y(_00705_));
 sky130_fd_sc_hd__nand2_1 _07926_ (.A(_00704_),
    .B(_00705_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_1 _07927_ (.A(_00699_),
    .B(_00706_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand3b_1 _07928_ (.A_N(_00706_),
    .B(_00697_),
    .C(_00698_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _07929_ (.A(_00707_),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _07930_ (.A(_00683_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand3_1 _07931_ (.A(_00682_),
    .B(_00707_),
    .C(_00708_),
    .Y(_00711_));
 sky130_fd_sc_hd__nand2_1 _07932_ (.A(_00710_),
    .B(_00711_),
    .Y(_00712_));
 sky130_fd_sc_hd__a21oi_1 _07933_ (.A1(_00574_),
    .A2(_00573_),
    .B1(_00570_),
    .Y(_00713_));
 sky130_fd_sc_hd__inv_2 _07934_ (.A(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _07935_ (.A(_00712_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__nand3_1 _07936_ (.A(_00710_),
    .B(_00711_),
    .C(_00713_),
    .Y(_00716_));
 sky130_fd_sc_hd__nand2_1 _07937_ (.A(_00715_),
    .B(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__inv_2 _07938_ (.A(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_1 _07939_ (.A(_00679_),
    .B(_00616_),
    .Y(_00719_));
 sky130_fd_sc_hd__nand3b_1 _07940_ (.A_N(_00680_),
    .B(_00718_),
    .C(_00719_),
    .Y(_00720_));
 sky130_fd_sc_hd__or2b_1 _07941_ (.A(_00616_),
    .B_N(_00679_),
    .X(_00721_));
 sky130_fd_sc_hd__nand3_1 _07942_ (.A(_00616_),
    .B(_00678_),
    .C(_00677_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand3_1 _07943_ (.A(_00721_),
    .B(_00722_),
    .C(_00717_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand2_2 _07944_ (.A(_00720_),
    .B(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__inv_2 _07945_ (.A(_00724_),
    .Y(_00725_));
 sky130_fd_sc_hd__nor2_1 _07946_ (.A(_00554_),
    .B(_00552_),
    .Y(_00726_));
 sky130_fd_sc_hd__a21oi_1 _07947_ (.A1(_00558_),
    .A2(_00588_),
    .B1(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__nand2_1 _07948_ (.A(_00725_),
    .B(_00727_),
    .Y(_00728_));
 sky130_fd_sc_hd__nand2_1 _07949_ (.A(_00586_),
    .B(_00583_),
    .Y(_00729_));
 sky130_fd_sc_hd__inv_2 _07950_ (.A(_00729_),
    .Y(_00730_));
 sky130_fd_sc_hd__o21ai_1 _07951_ (.A1(_00554_),
    .A2(_00552_),
    .B1(_00589_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _07952_ (.A(_00731_),
    .B(_00724_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand3_1 _07953_ (.A(_00728_),
    .B(_00730_),
    .C(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand2_1 _07954_ (.A(_00725_),
    .B(_00731_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _07955_ (.A(_00727_),
    .B(_00724_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand3_1 _07956_ (.A(_00734_),
    .B(_00729_),
    .C(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand2_1 _07957_ (.A(_00733_),
    .B(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__a21o_1 _07958_ (.A1(_00594_),
    .A2(_00451_),
    .B1(_00592_),
    .X(_00738_));
 sky130_fd_sc_hd__inv_2 _07959_ (.A(_00738_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _07960_ (.A(_00737_),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__nand3_1 _07961_ (.A(_00738_),
    .B(_00733_),
    .C(_00736_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand3_1 _07962_ (.A(_00615_),
    .B(_00740_),
    .C(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__nand2_1 _07963_ (.A(_00740_),
    .B(_00741_),
    .Y(_00743_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_00743_),
    .B(_00599_),
    .Y(_00744_));
 sky130_fd_sc_hd__nand3_1 _07965_ (.A(_00614_),
    .B(_00742_),
    .C(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__nand2_1 _07966_ (.A(_00742_),
    .B(_00744_),
    .Y(_00746_));
 sky130_fd_sc_hd__nand2_1 _07967_ (.A(_00746_),
    .B(_00603_),
    .Y(_00747_));
 sky130_fd_sc_hd__nand2_1 _07968_ (.A(_00745_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__inv_2 _07969_ (.A(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__nand2_1 _07970_ (.A(_00612_),
    .B(_00606_),
    .Y(_00750_));
 sky130_fd_sc_hd__xor2_1 _07971_ (.A(_00749_),
    .B(_00750_),
    .X(\m1.out[13] ));
 sky130_fd_sc_hd__nor2_1 _07972_ (.A(_00739_),
    .B(_00737_),
    .Y(_00751_));
 sky130_fd_sc_hd__nand2_1 _07973_ (.A(_00630_),
    .B(_00631_),
    .Y(_00752_));
 sky130_fd_sc_hd__nor2_1 _07974_ (.A(_00631_),
    .B(_00630_),
    .Y(_00753_));
 sky130_fd_sc_hd__a21oi_1 _07975_ (.A1(_00752_),
    .A2(_00648_),
    .B1(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__nand2_1 _07976_ (.A(net1),
    .B(net38),
    .Y(_00755_));
 sky130_fd_sc_hd__inv_2 _07977_ (.A(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__nand2_1 _07978_ (.A(_06268_),
    .B(_06217_),
    .Y(_00757_));
 sky130_fd_sc_hd__nand2_1 _07979_ (.A(_00756_),
    .B(_00757_),
    .Y(_00758_));
 sky130_fd_sc_hd__inv_2 _07980_ (.A(_00757_),
    .Y(_00759_));
 sky130_fd_sc_hd__nand2_1 _07981_ (.A(_00759_),
    .B(_00755_),
    .Y(_00760_));
 sky130_fd_sc_hd__nand2_1 _07982_ (.A(_06392_),
    .B(_06220_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand3_1 _07983_ (.A(_00758_),
    .B(_00760_),
    .C(_00761_),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _07984_ (.A(_00759_),
    .B(_00756_),
    .Y(_00763_));
 sky130_fd_sc_hd__inv_2 _07985_ (.A(_00761_),
    .Y(_00764_));
 sky130_fd_sc_hd__nand2_1 _07986_ (.A(_00757_),
    .B(_00755_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand3_1 _07987_ (.A(_00763_),
    .B(_00764_),
    .C(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hd__nand2_1 _07988_ (.A(_00762_),
    .B(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2_1 _07989_ (.A(_00619_),
    .B(_00621_),
    .Y(_00768_));
 sky130_fd_sc_hd__a21oi_2 _07990_ (.A1(_00624_),
    .A2(_00628_),
    .B1(_00768_),
    .Y(_00769_));
 sky130_fd_sc_hd__inv_2 _07991_ (.A(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hd__nand2_1 _07992_ (.A(_00767_),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__nand3_1 _07993_ (.A(_00769_),
    .B(_00762_),
    .C(_00766_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand2_1 _07994_ (.A(_06260_),
    .B(_06229_),
    .Y(_00773_));
 sky130_fd_sc_hd__inv_2 _07995_ (.A(_00773_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _07996_ (.A(_06272_),
    .B(_06227_),
    .Y(_00775_));
 sky130_fd_sc_hd__inv_2 _07997_ (.A(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand2_1 _07998_ (.A(_00774_),
    .B(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand2_1 _07999_ (.A(_00773_),
    .B(_00775_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _08000_ (.A(_00777_),
    .B(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hd__buf_4 _08001_ (.A(net64),
    .X(_00780_));
 sky130_fd_sc_hd__nand2_1 _08002_ (.A(_06258_),
    .B(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hd__nand2_1 _08003_ (.A(_00779_),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _08004_ (.A(_00781_),
    .Y(_00783_));
 sky130_fd_sc_hd__nand3_1 _08005_ (.A(_00777_),
    .B(_00783_),
    .C(_00778_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_1 _08006_ (.A(_00782_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand3_1 _08007_ (.A(_00771_),
    .B(_00772_),
    .C(_00785_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand3_1 _08008_ (.A(_00770_),
    .B(_00762_),
    .C(_00766_),
    .Y(_00787_));
 sky130_fd_sc_hd__nand2_1 _08009_ (.A(_00767_),
    .B(_00769_),
    .Y(_00788_));
 sky130_fd_sc_hd__inv_2 _08010_ (.A(_00785_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand3_1 _08011_ (.A(_00787_),
    .B(_00788_),
    .C(_00789_),
    .Y(_00790_));
 sky130_fd_sc_hd__nand3_1 _08012_ (.A(_00754_),
    .B(_00786_),
    .C(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hd__a21o_1 _08013_ (.A1(_00752_),
    .A2(_00648_),
    .B1(_00753_),
    .X(_00792_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(_00790_),
    .B(_00786_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_1 _08015_ (.A(_00792_),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand2_1 _08016_ (.A(_00791_),
    .B(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand2_1 _08017_ (.A(_00299_),
    .B(_06199_),
    .Y(_00796_));
 sky130_fd_sc_hd__inv_2 _08018_ (.A(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _08019_ (.A(_06265_),
    .B(_00270_),
    .Y(_00798_));
 sky130_fd_sc_hd__inv_2 _08020_ (.A(_00798_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_1 _08021_ (.A(_00797_),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hd__nand2_1 _08022_ (.A(_00796_),
    .B(_00798_),
    .Y(_00801_));
 sky130_fd_sc_hd__nand2_1 _08023_ (.A(_00800_),
    .B(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hd__nand2_1 _08024_ (.A(_00193_),
    .B(_06201_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand2_1 _08025_ (.A(_00802_),
    .B(_00803_),
    .Y(_00804_));
 sky130_fd_sc_hd__inv_2 _08026_ (.A(_00803_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand3_2 _08027_ (.A(_00800_),
    .B(_00805_),
    .C(_00801_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(_00804_),
    .B(_00806_),
    .Y(_00807_));
 sky130_fd_sc_hd__nor2_1 _08029_ (.A(_00636_),
    .B(_00638_),
    .Y(_00808_));
 sky130_fd_sc_hd__a21oi_1 _08030_ (.A1(_00641_),
    .A2(_00645_),
    .B1(_00808_),
    .Y(_00809_));
 sky130_fd_sc_hd__nand2_1 _08031_ (.A(_00807_),
    .B(_00809_),
    .Y(_00810_));
 sky130_fd_sc_hd__a21o_1 _08032_ (.A1(_00641_),
    .A2(_00645_),
    .B1(_00808_),
    .X(_00811_));
 sky130_fd_sc_hd__nand3_1 _08033_ (.A(_00811_),
    .B(_00806_),
    .C(_00804_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _08034_ (.A(_00664_),
    .B(_00659_),
    .Y(_00813_));
 sky130_fd_sc_hd__nand3_1 _08035_ (.A(_00810_),
    .B(_00812_),
    .C(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _08036_ (.A(_00807_),
    .B(_00811_),
    .Y(_00815_));
 sky130_fd_sc_hd__nand3_1 _08037_ (.A(_00804_),
    .B(_00809_),
    .C(_00806_),
    .Y(_00816_));
 sky130_fd_sc_hd__inv_2 _08038_ (.A(_00813_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand3_1 _08039_ (.A(_00815_),
    .B(_00816_),
    .C(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _08040_ (.A(_00814_),
    .B(_00818_),
    .Y(_00819_));
 sky130_fd_sc_hd__inv_2 _08041_ (.A(_00819_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand2_1 _08042_ (.A(_00795_),
    .B(_00820_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand3_1 _08043_ (.A(_00791_),
    .B(_00794_),
    .C(_00819_),
    .Y(_00822_));
 sky130_fd_sc_hd__nand2_2 _08044_ (.A(_00821_),
    .B(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__inv_2 _08045_ (.A(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__nand2_1 _08046_ (.A(_00618_),
    .B(_00651_),
    .Y(_00825_));
 sky130_fd_sc_hd__nor2_1 _08047_ (.A(_00651_),
    .B(_00618_),
    .Y(_00826_));
 sky130_fd_sc_hd__a21oi_2 _08048_ (.A1(_00825_),
    .A2(_00676_),
    .B1(_00826_),
    .Y(_00827_));
 sky130_fd_sc_hd__nand2_1 _08049_ (.A(_00824_),
    .B(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hd__nor2_1 _08050_ (.A(_00666_),
    .B(_00665_),
    .Y(_00829_));
 sky130_fd_sc_hd__a21oi_1 _08051_ (.A1(_00667_),
    .A2(_00673_),
    .B1(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_1 _08052_ (.A(_00439_),
    .B(_00176_),
    .Y(_00831_));
 sky130_fd_sc_hd__inv_2 _08053_ (.A(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__nand2_1 _08054_ (.A(_06287_),
    .B(_06196_),
    .Y(_00833_));
 sky130_fd_sc_hd__inv_2 _08055_ (.A(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__nand2_1 _08056_ (.A(_00832_),
    .B(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__nand2_1 _08057_ (.A(_00831_),
    .B(_00833_),
    .Y(_00836_));
 sky130_fd_sc_hd__nand2_1 _08058_ (.A(_00835_),
    .B(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__nand2_1 _08059_ (.A(_06291_),
    .B(_06211_),
    .Y(_00838_));
 sky130_fd_sc_hd__nand2_1 _08060_ (.A(_00837_),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__inv_2 _08061_ (.A(_00838_),
    .Y(_00840_));
 sky130_fd_sc_hd__nand3_1 _08062_ (.A(_00835_),
    .B(_00840_),
    .C(_00836_),
    .Y(_00841_));
 sky130_fd_sc_hd__nand2_1 _08063_ (.A(_00839_),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__a21o_1 _08064_ (.A1(_00687_),
    .A2(_00691_),
    .B1(_00686_),
    .X(_00843_));
 sky130_fd_sc_hd__nand2_1 _08065_ (.A(_00842_),
    .B(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__a21oi_1 _08066_ (.A1(_00687_),
    .A2(_00691_),
    .B1(_00686_),
    .Y(_00845_));
 sky130_fd_sc_hd__nand3_1 _08067_ (.A(_00839_),
    .B(_00845_),
    .C(_00841_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _08068_ (.A(_00701_),
    .B(_06204_),
    .Y(_00847_));
 sky130_fd_sc_hd__inv_2 _08069_ (.A(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hd__buf_6 _08070_ (.A(net4),
    .X(_00849_));
 sky130_fd_sc_hd__nand2_1 _08071_ (.A(_00849_),
    .B(_06214_),
    .Y(_00850_));
 sky130_fd_sc_hd__inv_2 _08072_ (.A(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__nand2_1 _08073_ (.A(_00848_),
    .B(_00851_),
    .Y(_00852_));
 sky130_fd_sc_hd__nand2_1 _08074_ (.A(_00847_),
    .B(_00850_),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_1 _08075_ (.A(_00852_),
    .B(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__nand2_1 _08076_ (.A(_06284_),
    .B(_06207_),
    .Y(_00855_));
 sky130_fd_sc_hd__nand2_1 _08077_ (.A(_00854_),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand3b_1 _08078_ (.A_N(_00855_),
    .B(_00852_),
    .C(_00853_),
    .Y(_00857_));
 sky130_fd_sc_hd__nand2_1 _08079_ (.A(_00856_),
    .B(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__nand3_1 _08080_ (.A(_00844_),
    .B(_00846_),
    .C(_00858_),
    .Y(_00859_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_00842_),
    .B(_00845_),
    .Y(_00860_));
 sky130_fd_sc_hd__nand3_1 _08082_ (.A(_00843_),
    .B(_00841_),
    .C(_00839_),
    .Y(_00861_));
 sky130_fd_sc_hd__nand3b_1 _08083_ (.A_N(_00858_),
    .B(_00860_),
    .C(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand3_1 _08084_ (.A(_00830_),
    .B(_00859_),
    .C(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__nand2_1 _08085_ (.A(_00862_),
    .B(_00859_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2_1 _08086_ (.A(_00674_),
    .B(_00669_),
    .Y(_00865_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(_00864_),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__nand2_1 _08088_ (.A(_00863_),
    .B(_00866_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2_1 _08089_ (.A(_00708_),
    .B(_00698_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _08090_ (.A(_00867_),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _08091_ (.A(_00868_),
    .Y(_00870_));
 sky130_fd_sc_hd__nand3_1 _08092_ (.A(_00870_),
    .B(_00863_),
    .C(_00866_),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_1 _08093_ (.A(_00869_),
    .B(_00871_),
    .Y(_00872_));
 sky130_fd_sc_hd__inv_2 _08094_ (.A(_00827_),
    .Y(_00873_));
 sky130_fd_sc_hd__nand2_1 _08095_ (.A(_00873_),
    .B(_00823_),
    .Y(_00874_));
 sky130_fd_sc_hd__nand3_1 _08096_ (.A(_00828_),
    .B(_00872_),
    .C(_00874_),
    .Y(_00875_));
 sky130_fd_sc_hd__nand2_1 _08097_ (.A(_00824_),
    .B(_00873_),
    .Y(_00876_));
 sky130_fd_sc_hd__inv_2 _08098_ (.A(_00872_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_1 _08099_ (.A(_00823_),
    .B(_00827_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand3_1 _08100_ (.A(_00876_),
    .B(_00877_),
    .C(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _08101_ (.A(_00875_),
    .B(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__a21oi_2 _08102_ (.A1(_00719_),
    .A2(_00718_),
    .B1(_00680_),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2_1 _08103_ (.A(_00880_),
    .B(_00881_),
    .Y(_00882_));
 sky130_fd_sc_hd__o21a_1 _08104_ (.A1(_00709_),
    .A2(_00682_),
    .B1(_00715_),
    .X(_00883_));
 sky130_fd_sc_hd__xor2_1 _08105_ (.A(_00704_),
    .B(_00883_),
    .X(_00884_));
 sky130_fd_sc_hd__nand2_1 _08106_ (.A(_00881_),
    .B(_00880_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand3b_1 _08107_ (.A_N(_00882_),
    .B(_00884_),
    .C(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand2b_1 _08108_ (.A_N(_00881_),
    .B(_00880_),
    .Y(_00887_));
 sky130_fd_sc_hd__nand2b_1 _08109_ (.A_N(_00880_),
    .B(_00881_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand3b_1 _08110_ (.A_N(_00884_),
    .B(_00887_),
    .C(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__nand2_1 _08111_ (.A(_00886_),
    .B(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__inv_2 _08112_ (.A(_00890_),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2_1 _08113_ (.A(_00724_),
    .B(_00727_),
    .Y(_00892_));
 sky130_fd_sc_hd__a21oi_1 _08114_ (.A1(_00735_),
    .A2(_00729_),
    .B1(_00892_),
    .Y(_00893_));
 sky130_fd_sc_hd__inv_2 _08115_ (.A(_00893_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_2 _08116_ (.A(_00891_),
    .B(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__nand2_1 _08117_ (.A(_00890_),
    .B(_00893_),
    .Y(_00896_));
 sky130_fd_sc_hd__nand3_2 _08118_ (.A(_00751_),
    .B(_00895_),
    .C(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__nand2_1 _08119_ (.A(_00895_),
    .B(_00896_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand2_1 _08120_ (.A(_00898_),
    .B(_00741_),
    .Y(_00899_));
 sky130_fd_sc_hd__nand2_1 _08121_ (.A(_00897_),
    .B(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hd__nand2_1 _08122_ (.A(_00900_),
    .B(_00742_),
    .Y(_00901_));
 sky130_fd_sc_hd__nor2_1 _08123_ (.A(_00599_),
    .B(_00743_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand3_1 _08124_ (.A(_00902_),
    .B(_00899_),
    .C(_00897_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand2_1 _08125_ (.A(_00901_),
    .B(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hd__inv_2 _08126_ (.A(_00904_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2_1 _08127_ (.A(_00611_),
    .B(_00749_),
    .Y(_00906_));
 sky130_fd_sc_hd__nor2_1 _08128_ (.A(_00471_),
    .B(_00607_),
    .Y(_00907_));
 sky130_fd_sc_hd__a21boi_1 _08129_ (.A1(_00907_),
    .A2(_00747_),
    .B1_N(_00745_),
    .Y(_00908_));
 sky130_fd_sc_hd__o21ai_1 _08130_ (.A1(_00906_),
    .A2(_00485_),
    .B1(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__or2_1 _08131_ (.A(_00905_),
    .B(_00909_),
    .X(_00910_));
 sky130_fd_sc_hd__nand2_1 _08132_ (.A(_00909_),
    .B(_00905_),
    .Y(_00911_));
 sky130_fd_sc_hd__and2_1 _08133_ (.A(_00910_),
    .B(_00911_),
    .X(_00912_));
 sky130_fd_sc_hd__clkbuf_1 _08134_ (.A(_00912_),
    .X(\m1.out[14] ));
 sky130_fd_sc_hd__a21oi_2 _08135_ (.A1(_00885_),
    .A2(_00884_),
    .B1(_00882_),
    .Y(_00913_));
 sky130_fd_sc_hd__nor2_1 _08136_ (.A(_00827_),
    .B(_00823_),
    .Y(_00914_));
 sky130_fd_sc_hd__a21oi_1 _08137_ (.A1(_00878_),
    .A2(_00877_),
    .B1(_00914_),
    .Y(_00915_));
 sky130_fd_sc_hd__nor2_1 _08138_ (.A(_00769_),
    .B(_00767_),
    .Y(_00916_));
 sky130_fd_sc_hd__a21oi_2 _08139_ (.A1(_00788_),
    .A2(_00789_),
    .B1(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__buf_6 _08140_ (.A(net39),
    .X(_00918_));
 sky130_fd_sc_hd__nand2_1 _08141_ (.A(_06270_),
    .B(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__inv_2 _08142_ (.A(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__buf_6 _08143_ (.A(net38),
    .X(_00921_));
 sky130_fd_sc_hd__nand2_2 _08144_ (.A(_06327_),
    .B(_00921_),
    .Y(_00922_));
 sky130_fd_sc_hd__nand2_1 _08145_ (.A(_00920_),
    .B(_00922_),
    .Y(_00923_));
 sky130_fd_sc_hd__inv_2 _08146_ (.A(_00922_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand2_1 _08147_ (.A(_00924_),
    .B(_00919_),
    .Y(_00925_));
 sky130_fd_sc_hd__buf_6 _08148_ (.A(_06217_),
    .X(_00926_));
 sky130_fd_sc_hd__nand2_1 _08149_ (.A(_06392_),
    .B(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand3_1 _08150_ (.A(_00923_),
    .B(_00925_),
    .C(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _08151_ (.A(_00924_),
    .B(_00920_),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _08152_ (.A(_00927_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _08153_ (.A(_00922_),
    .B(_00919_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand3_1 _08154_ (.A(_00929_),
    .B(_00930_),
    .C(_00931_),
    .Y(_00932_));
 sky130_fd_sc_hd__nand2_1 _08155_ (.A(_00928_),
    .B(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__nor2_1 _08156_ (.A(_00757_),
    .B(_00755_),
    .Y(_00934_));
 sky130_fd_sc_hd__a21oi_2 _08157_ (.A1(_00765_),
    .A2(_00764_),
    .B1(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__inv_2 _08158_ (.A(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__nand2_1 _08159_ (.A(_00933_),
    .B(_00936_),
    .Y(_00937_));
 sky130_fd_sc_hd__nand3_1 _08160_ (.A(_00935_),
    .B(_00928_),
    .C(_00932_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand2_1 _08161_ (.A(_06260_),
    .B(_06227_),
    .Y(_00939_));
 sky130_fd_sc_hd__inv_2 _08162_ (.A(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand2_1 _08163_ (.A(_06272_),
    .B(_06219_),
    .Y(_00941_));
 sky130_fd_sc_hd__inv_2 _08164_ (.A(_00941_),
    .Y(_00942_));
 sky130_fd_sc_hd__nand2_1 _08165_ (.A(_00940_),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _08166_ (.A(_00939_),
    .B(_00941_),
    .Y(_00944_));
 sky130_fd_sc_hd__nand2_1 _08167_ (.A(_00943_),
    .B(_00944_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _08168_ (.A(_06258_),
    .B(_06229_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _08169_ (.A(_00945_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__inv_2 _08170_ (.A(_00946_),
    .Y(_00948_));
 sky130_fd_sc_hd__nand3_1 _08171_ (.A(_00943_),
    .B(_00948_),
    .C(_00944_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_1 _08172_ (.A(_00947_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand3_1 _08173_ (.A(_00937_),
    .B(_00938_),
    .C(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand2_1 _08174_ (.A(_00937_),
    .B(_00938_),
    .Y(_00952_));
 sky130_fd_sc_hd__inv_2 _08175_ (.A(_00950_),
    .Y(_00953_));
 sky130_fd_sc_hd__nand2_1 _08176_ (.A(_00952_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__nand3_1 _08177_ (.A(_00917_),
    .B(_00951_),
    .C(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_1 _08178_ (.A(_00954_),
    .B(_00951_),
    .Y(_00956_));
 sky130_fd_sc_hd__nand2_1 _08179_ (.A(_00790_),
    .B(_00787_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2_1 _08180_ (.A(_00956_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hd__nand2_1 _08181_ (.A(_00955_),
    .B(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__nand2_1 _08182_ (.A(_00299_),
    .B(_00270_),
    .Y(_00960_));
 sky130_fd_sc_hd__inv_2 _08183_ (.A(_00960_),
    .Y(_00961_));
 sky130_fd_sc_hd__nand2_1 _08184_ (.A(_06265_),
    .B(net64),
    .Y(_00962_));
 sky130_fd_sc_hd__inv_2 _08185_ (.A(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _08186_ (.A(_00961_),
    .B(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__nand2_1 _08187_ (.A(_00960_),
    .B(_00962_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _08188_ (.A(_00964_),
    .B(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hd__nand2_1 _08189_ (.A(_00193_),
    .B(_06200_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand2_1 _08190_ (.A(_00966_),
    .B(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hd__inv_2 _08191_ (.A(_00967_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand3_2 _08192_ (.A(_00964_),
    .B(_00969_),
    .C(_00965_),
    .Y(_00970_));
 sky130_fd_sc_hd__nand2_1 _08193_ (.A(_00968_),
    .B(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__nor2_1 _08194_ (.A(_00773_),
    .B(_00775_),
    .Y(_00972_));
 sky130_fd_sc_hd__a21oi_2 _08195_ (.A1(_00778_),
    .A2(_00783_),
    .B1(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__inv_2 _08196_ (.A(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand2_1 _08197_ (.A(_00971_),
    .B(_00974_),
    .Y(_00975_));
 sky130_fd_sc_hd__nand3_1 _08198_ (.A(_00968_),
    .B(_00973_),
    .C(_00970_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_1 _08199_ (.A(_00975_),
    .B(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_2 _08200_ (.A(_00806_),
    .B(_00800_),
    .Y(_00978_));
 sky130_fd_sc_hd__nand2_1 _08201_ (.A(_00977_),
    .B(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__inv_2 _08202_ (.A(_00978_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand3_1 _08203_ (.A(_00975_),
    .B(_00976_),
    .C(_00980_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_1 _08204_ (.A(_00979_),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__inv_2 _08205_ (.A(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__nand2_1 _08206_ (.A(_00959_),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand3_1 _08207_ (.A(_00955_),
    .B(_00958_),
    .C(_00982_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand2_1 _08208_ (.A(_00984_),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _08209_ (.A(_00793_),
    .B(_00754_),
    .Y(_00987_));
 sky130_fd_sc_hd__nor2_1 _08210_ (.A(_00754_),
    .B(_00793_),
    .Y(_00988_));
 sky130_fd_sc_hd__a21o_1 _08211_ (.A1(_00987_),
    .A2(_00820_),
    .B1(_00988_),
    .X(_00989_));
 sky130_fd_sc_hd__nand2_1 _08212_ (.A(_00986_),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__a21oi_2 _08213_ (.A1(_00987_),
    .A2(_00820_),
    .B1(_00988_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand3_1 _08214_ (.A(_00991_),
    .B(_00984_),
    .C(_00985_),
    .Y(_00992_));
 sky130_fd_sc_hd__nor2_1 _08215_ (.A(_00809_),
    .B(_00807_),
    .Y(_00993_));
 sky130_fd_sc_hd__a21oi_2 _08216_ (.A1(_00810_),
    .A2(_00813_),
    .B1(_00993_),
    .Y(_00994_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_00439_),
    .B(_06195_),
    .Y(_00995_));
 sky130_fd_sc_hd__inv_2 _08218_ (.A(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hd__nand2_1 _08219_ (.A(_06287_),
    .B(_06201_),
    .Y(_00997_));
 sky130_fd_sc_hd__inv_2 _08220_ (.A(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hd__nand2_1 _08221_ (.A(_00996_),
    .B(_00998_),
    .Y(_00999_));
 sky130_fd_sc_hd__nand2_1 _08222_ (.A(_00995_),
    .B(_00997_),
    .Y(_01000_));
 sky130_fd_sc_hd__nand2_1 _08223_ (.A(_00999_),
    .B(_01000_),
    .Y(_01001_));
 sky130_fd_sc_hd__nand2_1 _08224_ (.A(_00561_),
    .B(_06198_),
    .Y(_01002_));
 sky130_fd_sc_hd__nand2_1 _08225_ (.A(_01001_),
    .B(_01002_),
    .Y(_01003_));
 sky130_fd_sc_hd__inv_2 _08226_ (.A(_01002_),
    .Y(_01004_));
 sky130_fd_sc_hd__nand3_2 _08227_ (.A(_00999_),
    .B(_01004_),
    .C(_01000_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _08228_ (.A(_01003_),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__nor2_1 _08229_ (.A(_00831_),
    .B(_00833_),
    .Y(_01007_));
 sky130_fd_sc_hd__a21o_1 _08230_ (.A1(_00836_),
    .A2(_00840_),
    .B1(_01007_),
    .X(_01008_));
 sky130_fd_sc_hd__nand2_1 _08231_ (.A(_01006_),
    .B(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__a21oi_1 _08232_ (.A1(_00836_),
    .A2(_00840_),
    .B1(_01007_),
    .Y(_01010_));
 sky130_fd_sc_hd__nand3_1 _08233_ (.A(_01003_),
    .B(_01010_),
    .C(_01005_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand2_1 _08234_ (.A(_06278_),
    .B(_06213_),
    .Y(_01012_));
 sky130_fd_sc_hd__inv_2 _08235_ (.A(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _08236_ (.A(_00849_),
    .B(_06210_),
    .Y(_01014_));
 sky130_fd_sc_hd__inv_2 _08237_ (.A(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _08238_ (.A(_01013_),
    .B(_01015_),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _08239_ (.A(_01012_),
    .B(_01014_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _08240_ (.A(_01016_),
    .B(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2_1 _08241_ (.A(_06284_),
    .B(_06205_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2_1 _08242_ (.A(_01018_),
    .B(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand3b_1 _08243_ (.A_N(_01019_),
    .B(_01016_),
    .C(_01017_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _08244_ (.A(_01020_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand3_1 _08245_ (.A(_01009_),
    .B(_01011_),
    .C(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__nand2_1 _08246_ (.A(_01006_),
    .B(_01010_),
    .Y(_01024_));
 sky130_fd_sc_hd__nand3_1 _08247_ (.A(_01008_),
    .B(_01005_),
    .C(_01003_),
    .Y(_01025_));
 sky130_fd_sc_hd__inv_2 _08248_ (.A(_01022_),
    .Y(_01026_));
 sky130_fd_sc_hd__nand3_1 _08249_ (.A(_01024_),
    .B(_01025_),
    .C(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__nand3_1 _08250_ (.A(_00994_),
    .B(_01023_),
    .C(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand2_1 _08251_ (.A(_00814_),
    .B(_00812_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _08252_ (.A(_01027_),
    .B(_01023_),
    .Y(_01030_));
 sky130_fd_sc_hd__nand2_1 _08253_ (.A(_01029_),
    .B(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _08254_ (.A(_01028_),
    .B(_01031_),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_1 _08255_ (.A(_00862_),
    .B(_00861_),
    .Y(_01033_));
 sky130_fd_sc_hd__nand2_1 _08256_ (.A(_01032_),
    .B(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__nand3b_1 _08257_ (.A_N(_01033_),
    .B(_01028_),
    .C(_01031_),
    .Y(_01035_));
 sky130_fd_sc_hd__nand2_1 _08258_ (.A(_01034_),
    .B(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hd__nand3_1 _08259_ (.A(_00990_),
    .B(_00992_),
    .C(_01036_),
    .Y(_01037_));
 sky130_fd_sc_hd__nand3_1 _08260_ (.A(_00989_),
    .B(_00985_),
    .C(_00984_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand2_1 _08261_ (.A(_00986_),
    .B(_00991_),
    .Y(_01039_));
 sky130_fd_sc_hd__inv_2 _08262_ (.A(_01036_),
    .Y(_01040_));
 sky130_fd_sc_hd__nand3_1 _08263_ (.A(_01038_),
    .B(_01039_),
    .C(_01040_),
    .Y(_01041_));
 sky130_fd_sc_hd__nand3_1 _08264_ (.A(_00915_),
    .B(_01037_),
    .C(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__a21o_1 _08265_ (.A1(_00878_),
    .A2(_00877_),
    .B1(_00914_),
    .X(_01043_));
 sky130_fd_sc_hd__nand2_1 _08266_ (.A(_01041_),
    .B(_01037_),
    .Y(_01044_));
 sky130_fd_sc_hd__nand2_1 _08267_ (.A(_01043_),
    .B(_01044_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand2_1 _08268_ (.A(_01042_),
    .B(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2_1 _08269_ (.A(_06282_),
    .B(_06208_),
    .Y(_01047_));
 sky130_fd_sc_hd__and2_1 _08270_ (.A(_00857_),
    .B(_00852_),
    .X(_01048_));
 sky130_fd_sc_hd__nor2_1 _08271_ (.A(_01047_),
    .B(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__inv_2 _08272_ (.A(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand2_1 _08273_ (.A(_01048_),
    .B(_01047_),
    .Y(_01051_));
 sky130_fd_sc_hd__nand2_2 _08274_ (.A(_01050_),
    .B(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__o21ai_2 _08275_ (.A1(_00864_),
    .A2(_00830_),
    .B1(_00869_),
    .Y(_01053_));
 sky130_fd_sc_hd__xnor2_2 _08276_ (.A(_01052_),
    .B(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand2_1 _08277_ (.A(_01046_),
    .B(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__nand3b_1 _08278_ (.A_N(_01054_),
    .B(_01042_),
    .C(_01045_),
    .Y(_01056_));
 sky130_fd_sc_hd__nand2_1 _08279_ (.A(_01055_),
    .B(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__nor2_1 _08280_ (.A(_00913_),
    .B(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hd__nor2_1 _08281_ (.A(_00704_),
    .B(_00883_),
    .Y(_01059_));
 sky130_fd_sc_hd__nand2_1 _08282_ (.A(_01057_),
    .B(_00913_),
    .Y(_01060_));
 sky130_fd_sc_hd__nand3b_1 _08283_ (.A_N(_01058_),
    .B(_01059_),
    .C(_01060_),
    .Y(_01061_));
 sky130_fd_sc_hd__nand2b_1 _08284_ (.A_N(_00913_),
    .B(_01057_),
    .Y(_01062_));
 sky130_fd_sc_hd__nand3_1 _08285_ (.A(_00913_),
    .B(_01056_),
    .C(_01055_),
    .Y(_01063_));
 sky130_fd_sc_hd__nand3b_1 _08286_ (.A_N(_01059_),
    .B(_01062_),
    .C(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _08287_ (.A(_01061_),
    .B(_01064_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand2_1 _08288_ (.A(_01065_),
    .B(_00895_),
    .Y(_01066_));
 sky130_fd_sc_hd__inv_2 _08289_ (.A(_00895_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand3_2 _08290_ (.A(_01061_),
    .B(_01064_),
    .C(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__nand2_1 _08291_ (.A(_01066_),
    .B(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__nand2_1 _08292_ (.A(_01069_),
    .B(_00897_),
    .Y(_01070_));
 sky130_fd_sc_hd__nand3b_1 _08293_ (.A_N(_00897_),
    .B(_01066_),
    .C(_01068_),
    .Y(_01071_));
 sky130_fd_sc_hd__nand2_1 _08294_ (.A(_01070_),
    .B(_01071_),
    .Y(_01072_));
 sky130_fd_sc_hd__nand2_1 _08295_ (.A(_00911_),
    .B(_00903_),
    .Y(_01073_));
 sky130_fd_sc_hd__xnor2_1 _08296_ (.A(_01072_),
    .B(_01073_),
    .Y(\m1.out[15] ));
 sky130_fd_sc_hd__nor2_1 _08297_ (.A(_00991_),
    .B(_00986_),
    .Y(_01074_));
 sky130_fd_sc_hd__a21oi_2 _08298_ (.A1(_01039_),
    .A2(_01040_),
    .B1(_01074_),
    .Y(_01075_));
 sky130_fd_sc_hd__nand2_1 _08299_ (.A(_00933_),
    .B(_00935_),
    .Y(_01076_));
 sky130_fd_sc_hd__nor2_1 _08300_ (.A(_00935_),
    .B(_00933_),
    .Y(_01077_));
 sky130_fd_sc_hd__a21oi_1 _08301_ (.A1(_01076_),
    .A2(_00953_),
    .B1(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand2_1 _08302_ (.A(_06270_),
    .B(_06173_),
    .Y(_01079_));
 sky130_fd_sc_hd__inv_2 _08303_ (.A(_01079_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_1 _08304_ (.A(_06268_),
    .B(net39),
    .Y(_01081_));
 sky130_fd_sc_hd__nand2_1 _08305_ (.A(_01080_),
    .B(_01081_),
    .Y(_01082_));
 sky130_fd_sc_hd__inv_2 _08306_ (.A(_01081_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand2_1 _08307_ (.A(_01083_),
    .B(_01079_),
    .Y(_01084_));
 sky130_fd_sc_hd__nand2_1 _08308_ (.A(_06275_),
    .B(net38),
    .Y(_01085_));
 sky130_fd_sc_hd__nand3_1 _08309_ (.A(_01082_),
    .B(_01084_),
    .C(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__nand2_1 _08310_ (.A(_01083_),
    .B(_01080_),
    .Y(_01087_));
 sky130_fd_sc_hd__inv_2 _08311_ (.A(_01085_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2_1 _08312_ (.A(_01081_),
    .B(_01079_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand3_1 _08313_ (.A(_01087_),
    .B(_01088_),
    .C(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__nand2_1 _08314_ (.A(_01086_),
    .B(_01090_),
    .Y(_01091_));
 sky130_fd_sc_hd__nor2_1 _08315_ (.A(_00922_),
    .B(_00919_),
    .Y(_01092_));
 sky130_fd_sc_hd__a21oi_2 _08316_ (.A1(_00931_),
    .A2(_00930_),
    .B1(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__inv_2 _08317_ (.A(_01093_),
    .Y(_01094_));
 sky130_fd_sc_hd__nand2_1 _08318_ (.A(_01091_),
    .B(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__nand3_1 _08319_ (.A(_01093_),
    .B(_01086_),
    .C(_01090_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_1 _08320_ (.A(_06260_),
    .B(_06219_),
    .Y(_01097_));
 sky130_fd_sc_hd__inv_2 _08321_ (.A(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2_1 _08322_ (.A(_06272_),
    .B(_06217_),
    .Y(_01099_));
 sky130_fd_sc_hd__inv_2 _08323_ (.A(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_1 _08324_ (.A(_01098_),
    .B(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2_1 _08325_ (.A(_01097_),
    .B(_01099_),
    .Y(_01102_));
 sky130_fd_sc_hd__nand2_1 _08326_ (.A(_01101_),
    .B(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _08327_ (.A(_00175_),
    .B(_00376_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _08328_ (.A(_01103_),
    .B(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__inv_2 _08329_ (.A(_01104_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand3_1 _08330_ (.A(_01101_),
    .B(_01106_),
    .C(_01102_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand2_1 _08331_ (.A(_01105_),
    .B(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand3_1 _08332_ (.A(_01095_),
    .B(_01096_),
    .C(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_1 _08333_ (.A(_01095_),
    .B(_01096_),
    .Y(_01110_));
 sky130_fd_sc_hd__inv_2 _08334_ (.A(_01108_),
    .Y(_01111_));
 sky130_fd_sc_hd__nand2_1 _08335_ (.A(_01110_),
    .B(_01111_),
    .Y(_01112_));
 sky130_fd_sc_hd__nand3_1 _08336_ (.A(_01078_),
    .B(_01109_),
    .C(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__a21o_1 _08337_ (.A1(_01076_),
    .A2(_00953_),
    .B1(_01077_),
    .X(_01114_));
 sky130_fd_sc_hd__nand2_1 _08338_ (.A(_01112_),
    .B(_01109_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _08339_ (.A(_01114_),
    .B(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _08340_ (.A(_01113_),
    .B(_01116_),
    .Y(_01118_));
 sky130_fd_sc_hd__nand2_1 _08341_ (.A(_00949_),
    .B(_00943_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand2_1 _08342_ (.A(_00193_),
    .B(_00270_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _08343_ (.A(_06263_),
    .B(net64),
    .Y(_01121_));
 sky130_fd_sc_hd__inv_2 _08344_ (.A(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(net29),
    .B(_06229_),
    .Y(_01123_));
 sky130_fd_sc_hd__inv_2 _08346_ (.A(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nand2_1 _08347_ (.A(_01122_),
    .B(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand2_1 _08348_ (.A(_01121_),
    .B(_01123_),
    .Y(_01126_));
 sky130_fd_sc_hd__nand3b_2 _08349_ (.A_N(_01120_),
    .B(_01125_),
    .C(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _08350_ (.A(_01125_),
    .B(_01126_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_1 _08351_ (.A(_01129_),
    .B(_01120_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand3_2 _08352_ (.A(_01119_),
    .B(_01127_),
    .C(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__inv_2 _08353_ (.A(_01119_),
    .Y(_01132_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_01130_),
    .B(_01127_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand2_2 _08355_ (.A(_01132_),
    .B(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hd__nand2_1 _08356_ (.A(_01131_),
    .B(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_2 _08357_ (.A(_00970_),
    .B(_00964_),
    .Y(_01136_));
 sky130_fd_sc_hd__inv_2 _08358_ (.A(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand2_1 _08359_ (.A(_01135_),
    .B(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand3_1 _08360_ (.A(_01131_),
    .B(_01134_),
    .C(_01136_),
    .Y(_01140_));
 sky130_fd_sc_hd__nand2_1 _08361_ (.A(_01138_),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__inv_2 _08362_ (.A(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand2_1 _08363_ (.A(_01118_),
    .B(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__nand3_1 _08364_ (.A(_01113_),
    .B(_01116_),
    .C(_01141_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand2_1 _08365_ (.A(_01143_),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand2_1 _08366_ (.A(_00956_),
    .B(_00917_),
    .Y(_01146_));
 sky130_fd_sc_hd__nor2_1 _08367_ (.A(_00917_),
    .B(_00956_),
    .Y(_01147_));
 sky130_fd_sc_hd__a21o_1 _08368_ (.A1(_01146_),
    .A2(_00983_),
    .B1(_01147_),
    .X(_01148_));
 sky130_fd_sc_hd__nand2_1 _08369_ (.A(_01145_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__a21oi_1 _08370_ (.A1(_01146_),
    .A2(_00983_),
    .B1(_01147_),
    .Y(_01151_));
 sky130_fd_sc_hd__nand3_1 _08371_ (.A(_01151_),
    .B(_01144_),
    .C(_01143_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand2_1 _08372_ (.A(_00701_),
    .B(_06210_),
    .Y(_01153_));
 sky130_fd_sc_hd__nand2_1 _08373_ (.A(_00849_),
    .B(_00176_),
    .Y(_01154_));
 sky130_fd_sc_hd__or2_1 _08374_ (.A(_01153_),
    .B(_01154_),
    .X(_01155_));
 sky130_fd_sc_hd__nand2_1 _08375_ (.A(_01153_),
    .B(_01154_),
    .Y(_01156_));
 sky130_fd_sc_hd__nand2_1 _08376_ (.A(_01155_),
    .B(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hd__buf_4 _08377_ (.A(_06283_),
    .X(_01158_));
 sky130_fd_sc_hd__nand2_1 _08378_ (.A(_01158_),
    .B(_06214_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_1 _08379_ (.A(_01157_),
    .B(_01159_),
    .Y(_01160_));
 sky130_fd_sc_hd__inv_2 _08380_ (.A(_01159_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand3_1 _08381_ (.A(_01155_),
    .B(_01162_),
    .C(_01156_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _08382_ (.A(_01160_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__nand2_1 _08383_ (.A(_01005_),
    .B(_00999_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand2_1 _08384_ (.A(net2),
    .B(net61),
    .Y(_01166_));
 sky130_fd_sc_hd__inv_2 _08385_ (.A(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand2_1 _08386_ (.A(_06286_),
    .B(net62),
    .Y(_01168_));
 sky130_fd_sc_hd__inv_2 _08387_ (.A(_01168_),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_1 _08388_ (.A(_01167_),
    .B(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__nand2_1 _08389_ (.A(_01166_),
    .B(_01168_),
    .Y(_01171_));
 sky130_fd_sc_hd__nand2_1 _08390_ (.A(_01170_),
    .B(_01171_),
    .Y(_01173_));
 sky130_fd_sc_hd__nand2_1 _08391_ (.A(net3),
    .B(net60),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_1 _08392_ (.A(_01173_),
    .B(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__inv_2 _08393_ (.A(_01174_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand3_1 _08394_ (.A(_01170_),
    .B(_01176_),
    .C(_01171_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand3_1 _08395_ (.A(_01165_),
    .B(_01175_),
    .C(_01177_),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_1 _08396_ (.A(_01175_),
    .B(_01177_),
    .Y(_01179_));
 sky130_fd_sc_hd__a21boi_1 _08397_ (.A1(_01004_),
    .A2(_01000_),
    .B1_N(_00999_),
    .Y(_01180_));
 sky130_fd_sc_hd__nand2_1 _08398_ (.A(_01179_),
    .B(_01180_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand3b_1 _08399_ (.A_N(_01164_),
    .B(_01178_),
    .C(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__nand2_1 _08400_ (.A(_01178_),
    .B(_01181_),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _08401_ (.A(_01184_),
    .B(_01164_),
    .Y(_01185_));
 sky130_fd_sc_hd__nand2_1 _08402_ (.A(_01182_),
    .B(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _08403_ (.A(_00971_),
    .B(_00973_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_1 _08404_ (.A(_00973_),
    .B(_00971_),
    .Y(_01188_));
 sky130_fd_sc_hd__a21oi_4 _08405_ (.A1(_01187_),
    .A2(_00978_),
    .B1(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__inv_2 _08406_ (.A(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _08407_ (.A(_01186_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__nand3_1 _08408_ (.A(_01189_),
    .B(_01182_),
    .C(_01185_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _08409_ (.A(_01191_),
    .B(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_1 _08410_ (.A(_01027_),
    .B(_01025_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _08411_ (.A(_01193_),
    .B(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__nand3b_1 _08412_ (.A_N(_01195_),
    .B(_01191_),
    .C(_01192_),
    .Y(_01197_));
 sky130_fd_sc_hd__nand2_1 _08413_ (.A(_01196_),
    .B(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand3_1 _08414_ (.A(_01149_),
    .B(_01152_),
    .C(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__nand3_1 _08415_ (.A(_01148_),
    .B(_01144_),
    .C(_01143_),
    .Y(_01200_));
 sky130_fd_sc_hd__inv_2 _08416_ (.A(_01198_),
    .Y(_01201_));
 sky130_fd_sc_hd__nand2_1 _08417_ (.A(_01145_),
    .B(_01151_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand3_1 _08418_ (.A(_01200_),
    .B(_01201_),
    .C(_01202_),
    .Y(_01203_));
 sky130_fd_sc_hd__nand3_1 _08419_ (.A(_01075_),
    .B(_01199_),
    .C(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _08420_ (.A(_01203_),
    .B(_01199_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_1 _08421_ (.A(_01041_),
    .B(_01038_),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _08422_ (.A(_01206_),
    .B(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__nand2_1 _08423_ (.A(_01204_),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__and2_1 _08424_ (.A(_01021_),
    .B(_01016_),
    .X(_01210_));
 sky130_fd_sc_hd__buf_4 _08425_ (.A(_06237_),
    .X(_01211_));
 sky130_fd_sc_hd__and4_1 _08426_ (.A(_06282_),
    .B(_01211_),
    .C(_06204_),
    .D(_06207_),
    .X(_01212_));
 sky130_fd_sc_hd__inv_2 _08427_ (.A(_01212_),
    .Y(_01213_));
 sky130_fd_sc_hd__a22o_1 _08428_ (.A1(_06282_),
    .A2(_06205_),
    .B1(_06238_),
    .B2(_06208_),
    .X(_01214_));
 sky130_fd_sc_hd__nand2_1 _08429_ (.A(_01213_),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__nor2_1 _08430_ (.A(_01210_),
    .B(_01215_),
    .Y(_01217_));
 sky130_fd_sc_hd__inv_2 _08431_ (.A(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hd__nand2_1 _08432_ (.A(_01215_),
    .B(_01210_),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_1 _08433_ (.A(_01218_),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__or2_1 _08434_ (.A(_01050_),
    .B(_01220_),
    .X(_01221_));
 sky130_fd_sc_hd__nand2_1 _08435_ (.A(_01220_),
    .B(_01050_),
    .Y(_01222_));
 sky130_fd_sc_hd__nand2_1 _08436_ (.A(_01221_),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__o21a_1 _08437_ (.A1(_01030_),
    .A2(_00994_),
    .B1(_01034_),
    .X(_01224_));
 sky130_fd_sc_hd__nor2_2 _08438_ (.A(_01223_),
    .B(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_1 _08439_ (.A(_01224_),
    .B(_01223_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2b_1 _08440_ (.A(_01225_),
    .B_N(_01226_),
    .Y(_01228_));
 sky130_fd_sc_hd__nand2_1 _08441_ (.A(_01209_),
    .B(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__or2b_1 _08442_ (.A(_01225_),
    .B_N(_01226_),
    .X(_01230_));
 sky130_fd_sc_hd__nand3_1 _08443_ (.A(_01204_),
    .B(_01208_),
    .C(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_01229_),
    .B(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand2_1 _08445_ (.A(_01044_),
    .B(_00915_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_1 _08446_ (.A(_00915_),
    .B(_01044_),
    .Y(_01234_));
 sky130_fd_sc_hd__a21oi_4 _08447_ (.A1(_01233_),
    .A2(_01054_),
    .B1(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hd__inv_2 _08448_ (.A(_01235_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _08449_ (.A(_01232_),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand3_2 _08450_ (.A(_01235_),
    .B(_01229_),
    .C(_01231_),
    .Y(_01239_));
 sky130_fd_sc_hd__nand2_1 _08451_ (.A(_01237_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__inv_2 _08452_ (.A(_01053_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_2 _08453_ (.A(_01052_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__inv_2 _08454_ (.A(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__nand2_1 _08455_ (.A(_01240_),
    .B(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand3_1 _08456_ (.A(_01237_),
    .B(_01239_),
    .C(_01242_),
    .Y(_01245_));
 sky130_fd_sc_hd__nand2_1 _08457_ (.A(_01244_),
    .B(_01245_),
    .Y(_01246_));
 sky130_fd_sc_hd__a21o_1 _08458_ (.A1(_01060_),
    .A2(_01059_),
    .B1(_01058_),
    .X(_01247_));
 sky130_fd_sc_hd__nand2_1 _08459_ (.A(_01246_),
    .B(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__nand2_1 _08460_ (.A(_01240_),
    .B(_01242_),
    .Y(_01250_));
 sky130_fd_sc_hd__nand3_1 _08461_ (.A(_01237_),
    .B(_01239_),
    .C(_01243_),
    .Y(_01251_));
 sky130_fd_sc_hd__nand2_1 _08462_ (.A(_01250_),
    .B(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__a21oi_1 _08463_ (.A1(_01060_),
    .A2(_01059_),
    .B1(_01058_),
    .Y(_01253_));
 sky130_fd_sc_hd__nand2_1 _08464_ (.A(_01252_),
    .B(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__nand2_1 _08465_ (.A(_01248_),
    .B(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__nor2_1 _08466_ (.A(_01068_),
    .B(_01255_),
    .Y(_01256_));
 sky130_fd_sc_hd__inv_2 _08467_ (.A(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _08468_ (.A(_01255_),
    .B(_01068_),
    .Y(_01258_));
 sky130_fd_sc_hd__nand2_1 _08469_ (.A(_01257_),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__inv_2 _08470_ (.A(_01259_),
    .Y(_01261_));
 sky130_fd_sc_hd__o21ai_1 _08471_ (.A1(_00903_),
    .A2(_01072_),
    .B1(_01071_),
    .Y(_01262_));
 sky130_fd_sc_hd__nand3_1 _08472_ (.A(_00905_),
    .B(_01071_),
    .C(_01070_),
    .Y(_01263_));
 sky130_fd_sc_hd__nor2_1 _08473_ (.A(_00908_),
    .B(_01263_),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_1 _08474_ (.A(_01262_),
    .B(_01264_),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _08475_ (.A(_00906_),
    .B(_01263_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _08476_ (.A(_00484_),
    .B(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_4 _08477_ (.A(_01265_),
    .B(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__or2_1 _08478_ (.A(_01261_),
    .B(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__nand2_1 _08479_ (.A(_01268_),
    .B(_01261_),
    .Y(_01270_));
 sky130_fd_sc_hd__and2_1 _08480_ (.A(_01269_),
    .B(_01270_),
    .X(_01272_));
 sky130_fd_sc_hd__clkbuf_1 _08481_ (.A(_01272_),
    .X(\m1.out[16] ));
 sky130_fd_sc_hd__nand2_1 _08482_ (.A(_01232_),
    .B(_01235_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor2_1 _08483_ (.A(_01235_),
    .B(_01232_),
    .Y(_01274_));
 sky130_fd_sc_hd__a21o_1 _08484_ (.A1(_01273_),
    .A2(_01242_),
    .B1(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__nor2_1 _08485_ (.A(_01151_),
    .B(_01145_),
    .Y(_01276_));
 sky130_fd_sc_hd__a21oi_2 _08486_ (.A1(_01201_),
    .A2(_01202_),
    .B1(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__buf_4 _08487_ (.A(net40),
    .X(_01278_));
 sky130_fd_sc_hd__nand2_1 _08488_ (.A(_06327_),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__buf_4 _08489_ (.A(net41),
    .X(_01280_));
 sky130_fd_sc_hd__nand2_1 _08490_ (.A(_06270_),
    .B(_01280_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor2_1 _08491_ (.A(_01279_),
    .B(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_1 _08492_ (.A(_06392_),
    .B(_00918_),
    .Y(_01284_));
 sky130_fd_sc_hd__inv_2 _08493_ (.A(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__nand2_1 _08494_ (.A(_01279_),
    .B(_01282_),
    .Y(_01286_));
 sky130_fd_sc_hd__nand3b_1 _08495_ (.A_N(_01283_),
    .B(_01285_),
    .C(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__nand2b_1 _08496_ (.A_N(_01282_),
    .B(_01279_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand2b_1 _08497_ (.A_N(_01279_),
    .B(_01282_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand3_1 _08498_ (.A(_01288_),
    .B(_01289_),
    .C(_01284_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand2_1 _08499_ (.A(_01287_),
    .B(_01290_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_1 _08500_ (.A(_01081_),
    .B(_01079_),
    .Y(_01293_));
 sky130_fd_sc_hd__a21oi_4 _08501_ (.A1(_01089_),
    .A2(_01088_),
    .B1(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__nand2_1 _08502_ (.A(_01291_),
    .B(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__clkinvlp_2 _08503_ (.A(_01294_),
    .Y(_01296_));
 sky130_fd_sc_hd__nand3_1 _08504_ (.A(_01287_),
    .B(_01296_),
    .C(_01290_),
    .Y(_01297_));
 sky130_fd_sc_hd__nand2_1 _08505_ (.A(_06261_),
    .B(_06217_),
    .Y(_01298_));
 sky130_fd_sc_hd__nand2_1 _08506_ (.A(_06273_),
    .B(net38),
    .Y(_01299_));
 sky130_fd_sc_hd__nor2_1 _08507_ (.A(_01298_),
    .B(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__inv_2 _08508_ (.A(_01300_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_1 _08509_ (.A(_01298_),
    .B(_01299_),
    .Y(_01302_));
 sky130_fd_sc_hd__nand2_1 _08510_ (.A(_01301_),
    .B(_01302_),
    .Y(_01304_));
 sky130_fd_sc_hd__nand2_1 _08511_ (.A(_00175_),
    .B(_06220_),
    .Y(_01305_));
 sky130_fd_sc_hd__nand2_1 _08512_ (.A(_01304_),
    .B(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__inv_2 _08513_ (.A(_01305_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand3_1 _08514_ (.A(_01301_),
    .B(_01307_),
    .C(_01302_),
    .Y(_01308_));
 sky130_fd_sc_hd__nand2_1 _08515_ (.A(_01306_),
    .B(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__inv_2 _08516_ (.A(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand3_1 _08517_ (.A(_01295_),
    .B(_01297_),
    .C(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__nand2_1 _08518_ (.A(_01291_),
    .B(_01296_),
    .Y(_01312_));
 sky130_fd_sc_hd__nand3_1 _08519_ (.A(_01287_),
    .B(_01290_),
    .C(_01294_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand3_1 _08520_ (.A(_01312_),
    .B(_01309_),
    .C(_01313_),
    .Y(_01315_));
 sky130_fd_sc_hd__nand2_1 _08521_ (.A(_01311_),
    .B(_01315_),
    .Y(_01316_));
 sky130_fd_sc_hd__nand2_1 _08522_ (.A(_01091_),
    .B(_01093_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_1 _08523_ (.A(_01093_),
    .B(_01091_),
    .Y(_01318_));
 sky130_fd_sc_hd__a21oi_4 _08524_ (.A1(_01317_),
    .A2(_01111_),
    .B1(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__inv_2 _08525_ (.A(_01319_),
    .Y(_01320_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(_01316_),
    .B(_01320_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand3_1 _08527_ (.A(_01319_),
    .B(_01311_),
    .C(_01315_),
    .Y(_01322_));
 sky130_fd_sc_hd__nand2_1 _08528_ (.A(_01321_),
    .B(_01322_),
    .Y(_01323_));
 sky130_fd_sc_hd__nand2_1 _08529_ (.A(_01107_),
    .B(_01101_),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2_1 _08530_ (.A(_00299_),
    .B(_06229_),
    .Y(_01326_));
 sky130_fd_sc_hd__inv_2 _08531_ (.A(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__nand2_1 _08532_ (.A(_06265_),
    .B(_06227_),
    .Y(_01328_));
 sky130_fd_sc_hd__inv_2 _08533_ (.A(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__nand2_1 _08534_ (.A(_01327_),
    .B(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand2_1 _08535_ (.A(_01326_),
    .B(_01328_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _08536_ (.A(_01330_),
    .B(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand2_1 _08537_ (.A(_00193_),
    .B(_06225_),
    .Y(_01333_));
 sky130_fd_sc_hd__nand2_1 _08538_ (.A(_01332_),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__nand3b_2 _08539_ (.A_N(_01333_),
    .B(_01330_),
    .C(_01331_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand3_1 _08540_ (.A(_01324_),
    .B(_01334_),
    .C(_01335_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand2_1 _08541_ (.A(_01334_),
    .B(_01335_),
    .Y(_01338_));
 sky130_fd_sc_hd__a21boi_1 _08542_ (.A1(_01106_),
    .A2(_01102_),
    .B1_N(_01101_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand2_2 _08543_ (.A(_01338_),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _08544_ (.A(_01337_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand2_2 _08545_ (.A(_01127_),
    .B(_01125_),
    .Y(_01342_));
 sky130_fd_sc_hd__inv_2 _08546_ (.A(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hd__nand2_1 _08547_ (.A(_01341_),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand3_1 _08548_ (.A(_01337_),
    .B(_01340_),
    .C(_01342_),
    .Y(_01345_));
 sky130_fd_sc_hd__nand2_2 _08549_ (.A(_01344_),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__inv_2 _08550_ (.A(_01346_),
    .Y(_01348_));
 sky130_fd_sc_hd__nand2_1 _08551_ (.A(_01323_),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__nand3_1 _08552_ (.A(_01321_),
    .B(_01322_),
    .C(_01346_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand2_1 _08553_ (.A(_01349_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2_1 _08554_ (.A(_01115_),
    .B(_01078_),
    .Y(_01352_));
 sky130_fd_sc_hd__nor2_1 _08555_ (.A(_01078_),
    .B(_01115_),
    .Y(_01353_));
 sky130_fd_sc_hd__a21oi_4 _08556_ (.A1(_01142_),
    .A2(_01352_),
    .B1(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__inv_2 _08557_ (.A(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(_01351_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__nand3_1 _08559_ (.A(_01354_),
    .B(_01349_),
    .C(_01350_),
    .Y(_01357_));
 sky130_fd_sc_hd__nand2_1 _08560_ (.A(_01182_),
    .B(_01178_),
    .Y(_01359_));
 sky130_fd_sc_hd__nand2_1 _08561_ (.A(_06278_),
    .B(_06197_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _08562_ (.A(net4),
    .B(_06195_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2_1 _08563_ (.A(_01360_),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__inv_2 _08564_ (.A(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__nand2_1 _08565_ (.A(_01360_),
    .B(_01361_),
    .Y(_01364_));
 sky130_fd_sc_hd__nand2_1 _08566_ (.A(_01363_),
    .B(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_1 _08567_ (.A(_06283_),
    .B(_06210_),
    .Y(_01366_));
 sky130_fd_sc_hd__nand2_1 _08568_ (.A(_01365_),
    .B(_01366_),
    .Y(_01367_));
 sky130_fd_sc_hd__inv_2 _08569_ (.A(_01366_),
    .Y(_01368_));
 sky130_fd_sc_hd__nand3_1 _08570_ (.A(_01363_),
    .B(_01368_),
    .C(_01364_),
    .Y(_01370_));
 sky130_fd_sc_hd__nand2_1 _08571_ (.A(_01367_),
    .B(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__nand2_1 _08572_ (.A(net2),
    .B(net62),
    .Y(_01372_));
 sky130_fd_sc_hd__nand2_1 _08573_ (.A(_06286_),
    .B(net63),
    .Y(_01373_));
 sky130_fd_sc_hd__nor2_1 _08574_ (.A(_01372_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__inv_2 _08575_ (.A(_01374_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _08576_ (.A(_01372_),
    .B(_01373_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _08577_ (.A(_01375_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _08578_ (.A(net3),
    .B(_06201_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _08579_ (.A(_01377_),
    .B(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__inv_2 _08580_ (.A(_01378_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand3_2 _08581_ (.A(_01375_),
    .B(_01381_),
    .C(_01376_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand2_1 _08582_ (.A(_01379_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _08583_ (.A(_01166_),
    .B(_01168_),
    .Y(_01384_));
 sky130_fd_sc_hd__a21oi_2 _08584_ (.A1(_01171_),
    .A2(_01176_),
    .B1(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_1 _08585_ (.A(_01383_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__inv_2 _08586_ (.A(_01385_),
    .Y(_01387_));
 sky130_fd_sc_hd__nand3_1 _08587_ (.A(_01387_),
    .B(_01379_),
    .C(_01382_),
    .Y(_01388_));
 sky130_fd_sc_hd__nand3b_1 _08588_ (.A_N(_01371_),
    .B(_01386_),
    .C(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__nand2_1 _08589_ (.A(_01383_),
    .B(_01387_),
    .Y(_01390_));
 sky130_fd_sc_hd__nand3_1 _08590_ (.A(_01379_),
    .B(_01382_),
    .C(_01385_),
    .Y(_01392_));
 sky130_fd_sc_hd__nand3_1 _08591_ (.A(_01390_),
    .B(_01392_),
    .C(_01371_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand2_1 _08592_ (.A(_01389_),
    .B(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__inv_2 _08593_ (.A(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__a21boi_4 _08594_ (.A1(_01136_),
    .A2(_01134_),
    .B1_N(_01131_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand2_1 _08595_ (.A(_01395_),
    .B(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__inv_2 _08596_ (.A(_01396_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand2_1 _08597_ (.A(_01398_),
    .B(_01394_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand3b_1 _08598_ (.A_N(_01359_),
    .B(_01397_),
    .C(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2_1 _08599_ (.A(_01395_),
    .B(_01398_),
    .Y(_01401_));
 sky130_fd_sc_hd__nand2_1 _08600_ (.A(_01394_),
    .B(_01396_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand3_1 _08601_ (.A(_01401_),
    .B(_01359_),
    .C(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__nand2_1 _08602_ (.A(_01400_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hd__nand3_1 _08603_ (.A(_01356_),
    .B(_01357_),
    .C(_01405_),
    .Y(_01406_));
 sky130_fd_sc_hd__nand2_1 _08604_ (.A(_01356_),
    .B(_01357_),
    .Y(_01407_));
 sky130_fd_sc_hd__inv_2 _08605_ (.A(_01405_),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_1 _08606_ (.A(_01407_),
    .B(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand3_1 _08607_ (.A(_01277_),
    .B(_01406_),
    .C(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2_1 _08608_ (.A(_01409_),
    .B(_01406_),
    .Y(_01411_));
 sky130_fd_sc_hd__nand2_1 _08609_ (.A(_01203_),
    .B(_01200_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2_1 _08610_ (.A(_01411_),
    .B(_01412_),
    .Y(_01414_));
 sky130_fd_sc_hd__nand2_1 _08611_ (.A(_01410_),
    .B(_01414_),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2_1 _08612_ (.A(_01186_),
    .B(_01189_),
    .Y(_01416_));
 sky130_fd_sc_hd__nor2_1 _08613_ (.A(_01189_),
    .B(_01186_),
    .Y(_01417_));
 sky130_fd_sc_hd__a21oi_1 _08614_ (.A1(_01416_),
    .A2(_01195_),
    .B1(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__inv_2 _08615_ (.A(_01418_),
    .Y(_01419_));
 sky130_fd_sc_hd__nand2_1 _08616_ (.A(_06238_),
    .B(_06205_),
    .Y(_01420_));
 sky130_fd_sc_hd__nand3b_1 _08617_ (.A_N(_01420_),
    .B(_06282_),
    .C(_06215_),
    .Y(_01421_));
 sky130_fd_sc_hd__inv_2 _08618_ (.A(_06281_),
    .Y(_01422_));
 sky130_fd_sc_hd__o21ai_1 _08619_ (.A1(_01422_),
    .A2(_06331_),
    .B1(_01420_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _08620_ (.A(_01421_),
    .B(_01423_),
    .Y(_01425_));
 sky130_fd_sc_hd__nand2_1 _08621_ (.A(_06236_),
    .B(_06207_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _08622_ (.A(_01425_),
    .B(_01426_),
    .Y(_01427_));
 sky130_fd_sc_hd__nand3b_1 _08623_ (.A_N(_01426_),
    .B(_01421_),
    .C(_01423_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_1 _08624_ (.A(_01427_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_2 _08625_ (.A(_01163_),
    .B(_01155_),
    .Y(_01430_));
 sky130_fd_sc_hd__inv_2 _08626_ (.A(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_1 _08627_ (.A(_01429_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__nand3_1 _08628_ (.A(_01430_),
    .B(_01428_),
    .C(_01427_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _08629_ (.A(_01432_),
    .B(_01433_),
    .Y(_01434_));
 sky130_fd_sc_hd__nand2_1 _08630_ (.A(_01434_),
    .B(_01213_),
    .Y(_01436_));
 sky130_fd_sc_hd__nand3_1 _08631_ (.A(_01432_),
    .B(_01433_),
    .C(_01212_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _08632_ (.A(_01436_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__nand2_1 _08633_ (.A(_01438_),
    .B(_01218_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand3_2 _08634_ (.A(_01436_),
    .B(_01437_),
    .C(_01217_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand2_2 _08635_ (.A(_01439_),
    .B(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__inv_2 _08636_ (.A(_01441_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _08637_ (.A(_01419_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__nand2_1 _08638_ (.A(_01418_),
    .B(_01441_),
    .Y(_01444_));
 sky130_fd_sc_hd__nand2_1 _08639_ (.A(_01443_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _08640_ (.A(_01445_),
    .B(_01221_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand3b_1 _08641_ (.A_N(_01221_),
    .B(_01443_),
    .C(_01444_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _08642_ (.A(_01447_),
    .B(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__inv_2 _08643_ (.A(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand2_1 _08644_ (.A(_01415_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__nand3_1 _08645_ (.A(_01410_),
    .B(_01414_),
    .C(_01449_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand2_1 _08646_ (.A(_01451_),
    .B(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(_01206_),
    .B(_01075_),
    .Y(_01454_));
 sky130_fd_sc_hd__nor2_1 _08648_ (.A(_01075_),
    .B(_01206_),
    .Y(_01455_));
 sky130_fd_sc_hd__a21oi_2 _08649_ (.A1(_01454_),
    .A2(_01228_),
    .B1(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__inv_2 _08650_ (.A(_01456_),
    .Y(_01458_));
 sky130_fd_sc_hd__nand2_1 _08651_ (.A(_01453_),
    .B(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand3_1 _08652_ (.A(_01456_),
    .B(_01451_),
    .C(_01452_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand3b_1 _08653_ (.A_N(_01225_),
    .B(_01459_),
    .C(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand2_1 _08654_ (.A(_01459_),
    .B(_01460_),
    .Y(_01462_));
 sky130_fd_sc_hd__nand2_1 _08655_ (.A(_01462_),
    .B(_01225_),
    .Y(_01463_));
 sky130_fd_sc_hd__nand3_2 _08656_ (.A(_01275_),
    .B(_01461_),
    .C(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _08657_ (.A(_01463_),
    .B(_01461_),
    .Y(_01465_));
 sky130_fd_sc_hd__a21oi_1 _08658_ (.A1(_01273_),
    .A2(_01242_),
    .B1(_01274_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_1 _08659_ (.A(_01465_),
    .B(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _08660_ (.A(_01464_),
    .B(_01467_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(_01469_),
    .B(_01248_),
    .Y(_01470_));
 sky130_fd_sc_hd__nor2_1 _08662_ (.A(_01253_),
    .B(_01252_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand3_1 _08663_ (.A(_01464_),
    .B(_01471_),
    .C(_01467_),
    .Y(_01472_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(_01470_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__nand2_1 _08665_ (.A(_01270_),
    .B(_01257_),
    .Y(_01474_));
 sky130_fd_sc_hd__xnor2_1 _08666_ (.A(_01473_),
    .B(_01474_),
    .Y(\m1.out[17] ));
 sky130_fd_sc_hd__nor2_1 _08667_ (.A(_01294_),
    .B(_01291_),
    .Y(_01475_));
 sky130_fd_sc_hd__a21oi_2 _08668_ (.A1(_01295_),
    .A2(_01310_),
    .B1(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__nand2_1 _08669_ (.A(_06327_),
    .B(_06171_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2_1 _08670_ (.A(_06270_),
    .B(_06178_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_1 _08671_ (.A(_01477_),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2_1 _08672_ (.A(_01477_),
    .B(_01479_),
    .Y(_01481_));
 sky130_fd_sc_hd__inv_2 _08673_ (.A(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _08674_ (.A(_06392_),
    .B(_01278_),
    .Y(_01483_));
 sky130_fd_sc_hd__o21ai_1 _08675_ (.A1(_01480_),
    .A2(_01482_),
    .B1(_01483_),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_1 _08676_ (.A(_01480_),
    .B(_01482_),
    .Y(_01485_));
 sky130_fd_sc_hd__inv_2 _08677_ (.A(_01483_),
    .Y(_01486_));
 sky130_fd_sc_hd__nand2_1 _08678_ (.A(_01485_),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_1 _08679_ (.A(_01484_),
    .B(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__a21oi_2 _08680_ (.A1(_01286_),
    .A2(_01285_),
    .B1(_01283_),
    .Y(_01490_));
 sky130_fd_sc_hd__inv_2 _08681_ (.A(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _08682_ (.A(_01488_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand3_1 _08683_ (.A(_01484_),
    .B(_01487_),
    .C(_01490_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_06262_),
    .B(_00921_),
    .Y(_01494_));
 sky130_fd_sc_hd__nand2_1 _08685_ (.A(_06274_),
    .B(_00918_),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_1 _08686_ (.A(_01494_),
    .B(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand2_1 _08687_ (.A(_01494_),
    .B(_01495_),
    .Y(_01497_));
 sky130_fd_sc_hd__inv_2 _08688_ (.A(_01497_),
    .Y(_01498_));
 sky130_fd_sc_hd__nand2_1 _08689_ (.A(_00175_),
    .B(_00926_),
    .Y(_01499_));
 sky130_fd_sc_hd__o21ai_1 _08690_ (.A1(_01496_),
    .A2(_01498_),
    .B1(_01499_),
    .Y(_01501_));
 sky130_fd_sc_hd__inv_2 _08691_ (.A(_01499_),
    .Y(_01502_));
 sky130_fd_sc_hd__nand3b_1 _08692_ (.A_N(_01496_),
    .B(_01502_),
    .C(_01497_),
    .Y(_01503_));
 sky130_fd_sc_hd__nand2_1 _08693_ (.A(_01501_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__nand3_1 _08694_ (.A(_01492_),
    .B(_01493_),
    .C(_01504_),
    .Y(_01505_));
 sky130_fd_sc_hd__nand2_1 _08695_ (.A(_01492_),
    .B(_01493_),
    .Y(_01506_));
 sky130_fd_sc_hd__inv_2 _08696_ (.A(_01504_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(_01506_),
    .B(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__nand3_1 _08698_ (.A(_01476_),
    .B(_01505_),
    .C(_01508_),
    .Y(_01509_));
 sky130_fd_sc_hd__nand2_1 _08699_ (.A(_01508_),
    .B(_01505_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand2_1 _08700_ (.A(_01311_),
    .B(_01297_),
    .Y(_01512_));
 sky130_fd_sc_hd__nand2_1 _08701_ (.A(_01510_),
    .B(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_1 _08702_ (.A(_01509_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__nand2_1 _08703_ (.A(_01308_),
    .B(_01301_),
    .Y(_01515_));
 sky130_fd_sc_hd__inv_2 _08704_ (.A(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand2_1 _08705_ (.A(_06264_),
    .B(_00376_),
    .Y(_01517_));
 sky130_fd_sc_hd__nand2_1 _08706_ (.A(_06266_),
    .B(_06220_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor2_1 _08707_ (.A(_01517_),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand2_1 _08708_ (.A(_01517_),
    .B(_01518_),
    .Y(_01520_));
 sky130_fd_sc_hd__inv_2 _08709_ (.A(_01520_),
    .Y(_01521_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_06290_),
    .B(_06231_),
    .Y(_01523_));
 sky130_fd_sc_hd__o21ai_1 _08711_ (.A1(_01519_),
    .A2(_01521_),
    .B1(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__inv_2 _08712_ (.A(_01523_),
    .Y(_01525_));
 sky130_fd_sc_hd__nand3b_1 _08713_ (.A_N(_01519_),
    .B(_01525_),
    .C(_01520_),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_1 _08714_ (.A(_01524_),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand2_1 _08715_ (.A(_01516_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__nand3_1 _08716_ (.A(_01515_),
    .B(_01524_),
    .C(_01526_),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_1 _08717_ (.A(_01528_),
    .B(_01529_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand2_2 _08718_ (.A(_01335_),
    .B(_01330_),
    .Y(_01531_));
 sky130_fd_sc_hd__inv_2 _08719_ (.A(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand2_1 _08720_ (.A(_01530_),
    .B(_01532_),
    .Y(_01534_));
 sky130_fd_sc_hd__nand3_1 _08721_ (.A(_01528_),
    .B(_01529_),
    .C(_01531_),
    .Y(_01535_));
 sky130_fd_sc_hd__nand2_1 _08722_ (.A(_01534_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__inv_2 _08723_ (.A(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__nand2_1 _08724_ (.A(_01514_),
    .B(_01537_),
    .Y(_01538_));
 sky130_fd_sc_hd__nand3_1 _08725_ (.A(_01509_),
    .B(_01513_),
    .C(_01536_),
    .Y(_01539_));
 sky130_fd_sc_hd__nand2_1 _08726_ (.A(_01538_),
    .B(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand2_1 _08727_ (.A(_01316_),
    .B(_01319_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _08728_ (.A(_01319_),
    .B(_01316_),
    .Y(_01542_));
 sky130_fd_sc_hd__a21oi_4 _08729_ (.A1(_01541_),
    .A2(_01348_),
    .B1(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__inv_2 _08730_ (.A(_01543_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_1 _08731_ (.A(_01540_),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand3_1 _08732_ (.A(_01543_),
    .B(_01538_),
    .C(_01539_),
    .Y(_01547_));
 sky130_fd_sc_hd__nand2_1 _08733_ (.A(_01546_),
    .B(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__nand2_1 _08734_ (.A(_01382_),
    .B(_01375_),
    .Y(_01549_));
 sky130_fd_sc_hd__inv_2 _08735_ (.A(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__nand2_1 _08736_ (.A(_00439_),
    .B(_00270_),
    .Y(_01551_));
 sky130_fd_sc_hd__nand2_1 _08737_ (.A(_06287_),
    .B(_00780_),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _08738_ (.A(_01551_),
    .B(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_1 _08739_ (.A(_01551_),
    .B(_01552_),
    .Y(_01554_));
 sky130_fd_sc_hd__inv_2 _08740_ (.A(_01554_),
    .Y(_01556_));
 sky130_fd_sc_hd__nand2_1 _08741_ (.A(net3),
    .B(_06199_),
    .Y(_01557_));
 sky130_fd_sc_hd__o21ai_1 _08742_ (.A1(_01553_),
    .A2(_01556_),
    .B1(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__inv_2 _08743_ (.A(_01557_),
    .Y(_01559_));
 sky130_fd_sc_hd__nand3b_1 _08744_ (.A_N(_01553_),
    .B(_01559_),
    .C(_01554_),
    .Y(_01560_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(_01558_),
    .B(_01560_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _08746_ (.A(_01550_),
    .B(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__nand3_1 _08747_ (.A(_01549_),
    .B(_01558_),
    .C(_01560_),
    .Y(_01563_));
 sky130_fd_sc_hd__nand2_1 _08748_ (.A(_01562_),
    .B(_01563_),
    .Y(_01564_));
 sky130_fd_sc_hd__nand2_1 _08749_ (.A(_06279_),
    .B(_06196_),
    .Y(_01565_));
 sky130_fd_sc_hd__nand2_1 _08750_ (.A(_06280_),
    .B(_06202_),
    .Y(_01567_));
 sky130_fd_sc_hd__nor2_1 _08751_ (.A(_01565_),
    .B(_01567_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand2_1 _08752_ (.A(_01565_),
    .B(_01567_),
    .Y(_01569_));
 sky130_fd_sc_hd__inv_2 _08753_ (.A(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(_06284_),
    .B(_06198_),
    .Y(_01571_));
 sky130_fd_sc_hd__o21ai_1 _08755_ (.A1(_01568_),
    .A2(_01570_),
    .B1(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__inv_2 _08756_ (.A(_01571_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand3b_1 _08757_ (.A_N(_01568_),
    .B(_01573_),
    .C(_01569_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _08758_ (.A(_01572_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(_01564_),
    .B(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__nand3b_1 _08760_ (.A_N(_01575_),
    .B(_01562_),
    .C(_01563_),
    .Y(_01578_));
 sky130_fd_sc_hd__nand2_1 _08761_ (.A(_01576_),
    .B(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__a21boi_4 _08762_ (.A1(_01342_),
    .A2(_01340_),
    .B1_N(_01337_),
    .Y(_01580_));
 sky130_fd_sc_hd__inv_2 _08763_ (.A(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__nand2_1 _08764_ (.A(_01579_),
    .B(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__nand3_1 _08765_ (.A(_01580_),
    .B(_01576_),
    .C(_01578_),
    .Y(_01583_));
 sky130_fd_sc_hd__nand2_1 _08766_ (.A(_01582_),
    .B(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_1 _08767_ (.A(_01389_),
    .B(_01388_),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _08768_ (.A(_01584_),
    .B(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hd__nand3b_1 _08769_ (.A_N(_01585_),
    .B(_01582_),
    .C(_01583_),
    .Y(_01587_));
 sky130_fd_sc_hd__nand2_1 _08770_ (.A(_01586_),
    .B(_01587_),
    .Y(_01589_));
 sky130_fd_sc_hd__inv_2 _08771_ (.A(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__nand2_1 _08772_ (.A(_01548_),
    .B(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__nand3_1 _08773_ (.A(_01546_),
    .B(_01547_),
    .C(_01589_),
    .Y(_01592_));
 sky130_fd_sc_hd__nand2_1 _08774_ (.A(_01591_),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__nand2_1 _08775_ (.A(_01351_),
    .B(_01354_),
    .Y(_01594_));
 sky130_fd_sc_hd__nor2_1 _08776_ (.A(_01354_),
    .B(_01351_),
    .Y(_01595_));
 sky130_fd_sc_hd__a21o_1 _08777_ (.A1(_01408_),
    .A2(_01594_),
    .B1(_01595_),
    .X(_01596_));
 sky130_fd_sc_hd__nand2_1 _08778_ (.A(_01593_),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__a21oi_2 _08779_ (.A1(_01408_),
    .A2(_01594_),
    .B1(_01595_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand3_1 _08780_ (.A(_01598_),
    .B(_01592_),
    .C(_01591_),
    .Y(_01600_));
 sky130_fd_sc_hd__nand2_1 _08781_ (.A(_01597_),
    .B(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__nand2_1 _08782_ (.A(_01437_),
    .B(_01433_),
    .Y(_01602_));
 sky130_fd_sc_hd__nand2_1 _08783_ (.A(_01370_),
    .B(_01363_),
    .Y(_01603_));
 sky130_fd_sc_hd__inv_2 _08784_ (.A(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _08785_ (.A(_06238_),
    .B(_06215_),
    .Y(_01605_));
 sky130_fd_sc_hd__nand2_1 _08786_ (.A(_06282_),
    .B(_06211_),
    .Y(_01606_));
 sky130_fd_sc_hd__nor2_1 _08787_ (.A(_01605_),
    .B(_01606_),
    .Y(_01607_));
 sky130_fd_sc_hd__nand2_1 _08788_ (.A(_01605_),
    .B(_01606_),
    .Y(_01608_));
 sky130_fd_sc_hd__inv_2 _08789_ (.A(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_1 _08790_ (.A(_06235_),
    .B(_06204_),
    .Y(_01611_));
 sky130_fd_sc_hd__o21ai_1 _08791_ (.A1(_01607_),
    .A2(_01609_),
    .B1(_01611_),
    .Y(_01612_));
 sky130_fd_sc_hd__inv_2 _08792_ (.A(_01611_),
    .Y(_01613_));
 sky130_fd_sc_hd__nand3b_1 _08793_ (.A_N(_01607_),
    .B(_01613_),
    .C(_01608_),
    .Y(_01614_));
 sky130_fd_sc_hd__nand2_1 _08794_ (.A(_01612_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__nand2_1 _08795_ (.A(_01604_),
    .B(_01615_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand3_1 _08796_ (.A(_01603_),
    .B(_01612_),
    .C(_01614_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_01616_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _08798_ (.A(_01428_),
    .B(_01421_),
    .Y(_01619_));
 sky130_fd_sc_hd__inv_2 _08799_ (.A(_01619_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_1 _08800_ (.A(_01618_),
    .B(_01620_),
    .Y(_01622_));
 sky130_fd_sc_hd__nand3_1 _08801_ (.A(_01616_),
    .B(_01617_),
    .C(_01619_),
    .Y(_01623_));
 sky130_fd_sc_hd__nand3_1 _08802_ (.A(_01602_),
    .B(_01622_),
    .C(_01623_),
    .Y(_01624_));
 sky130_fd_sc_hd__a21boi_1 _08803_ (.A1(_01432_),
    .A2(_01212_),
    .B1_N(_01433_),
    .Y(_01625_));
 sky130_fd_sc_hd__nand2_1 _08804_ (.A(_01622_),
    .B(_01623_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_01625_),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__nand2_1 _08806_ (.A(_01624_),
    .B(_01627_),
    .Y(_01628_));
 sky130_fd_sc_hd__nand2_1 _08807_ (.A(_06243_),
    .B(_06209_),
    .Y(_01629_));
 sky130_fd_sc_hd__nand2_1 _08808_ (.A(_01628_),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__inv_2 _08809_ (.A(_01629_),
    .Y(_01631_));
 sky130_fd_sc_hd__nand3_1 _08810_ (.A(_01624_),
    .B(_01631_),
    .C(_01627_),
    .Y(_01633_));
 sky130_fd_sc_hd__nand2_1 _08811_ (.A(_01630_),
    .B(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__nand2_2 _08812_ (.A(_01404_),
    .B(_01401_),
    .Y(_01635_));
 sky130_fd_sc_hd__inv_2 _08813_ (.A(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__nand2_1 _08814_ (.A(_01634_),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__nand3_1 _08815_ (.A(_01635_),
    .B(_01630_),
    .C(_01633_),
    .Y(_01638_));
 sky130_fd_sc_hd__nand2_1 _08816_ (.A(_01637_),
    .B(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2_1 _08817_ (.A(_01639_),
    .B(_01440_),
    .Y(_01640_));
 sky130_fd_sc_hd__nand3b_1 _08818_ (.A_N(_01440_),
    .B(_01637_),
    .C(_01638_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _08819_ (.A(_01640_),
    .B(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__inv_2 _08820_ (.A(_01642_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _08821_ (.A(_01601_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__nand3_1 _08822_ (.A(_01597_),
    .B(_01600_),
    .C(_01642_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _08823_ (.A(_01645_),
    .B(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__nand2_1 _08824_ (.A(_01411_),
    .B(_01277_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_1 _08825_ (.A(_01277_),
    .B(_01411_),
    .Y(_01649_));
 sky130_fd_sc_hd__a21oi_4 _08826_ (.A1(_01648_),
    .A2(_01450_),
    .B1(_01649_),
    .Y(_01650_));
 sky130_fd_sc_hd__inv_2 _08827_ (.A(_01650_),
    .Y(_01651_));
 sky130_fd_sc_hd__nand2_1 _08828_ (.A(_01647_),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand3_1 _08829_ (.A(_01650_),
    .B(_01645_),
    .C(_01646_),
    .Y(_01653_));
 sky130_fd_sc_hd__nand2_1 _08830_ (.A(_01652_),
    .B(_01653_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_2 _08831_ (.A(_01448_),
    .B(_01443_),
    .Y(_01656_));
 sky130_fd_sc_hd__nand2_1 _08832_ (.A(_01655_),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__inv_2 _08833_ (.A(_01656_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand3_1 _08834_ (.A(_01652_),
    .B(_01653_),
    .C(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _08835_ (.A(_01657_),
    .B(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _08836_ (.A(_01453_),
    .B(_01456_),
    .Y(_01661_));
 sky130_fd_sc_hd__nor2_1 _08837_ (.A(_01456_),
    .B(_01453_),
    .Y(_01662_));
 sky130_fd_sc_hd__a21oi_2 _08838_ (.A1(_01661_),
    .A2(_01225_),
    .B1(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__nand2_1 _08839_ (.A(_01660_),
    .B(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__nand2_1 _08840_ (.A(_01655_),
    .B(_01658_),
    .Y(_01666_));
 sky130_fd_sc_hd__nand3_1 _08841_ (.A(_01652_),
    .B(_01653_),
    .C(_01656_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _08842_ (.A(_01666_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__inv_2 _08843_ (.A(_01663_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand2_2 _08844_ (.A(_01668_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _08845_ (.A(_01664_),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _08846_ (.A(_01671_),
    .B(_01464_),
    .Y(_01672_));
 sky130_fd_sc_hd__nor2_1 _08847_ (.A(_01466_),
    .B(_01465_),
    .Y(_01673_));
 sky130_fd_sc_hd__nand3_1 _08848_ (.A(_01664_),
    .B(_01670_),
    .C(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_1 _08849_ (.A(_01672_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__inv_2 _08850_ (.A(_01675_),
    .Y(_01677_));
 sky130_fd_sc_hd__nor2_1 _08851_ (.A(_01473_),
    .B(_01259_),
    .Y(_01678_));
 sky130_fd_sc_hd__nand3_1 _08852_ (.A(_01470_),
    .B(_01256_),
    .C(_01472_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _08853_ (.A(_01679_),
    .B(_01472_),
    .Y(_01680_));
 sky130_fd_sc_hd__a21o_1 _08854_ (.A1(_01268_),
    .A2(_01678_),
    .B1(_01680_),
    .X(_01681_));
 sky130_fd_sc_hd__or2_1 _08855_ (.A(_01677_),
    .B(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__nand2_1 _08856_ (.A(_01681_),
    .B(_01677_),
    .Y(_01683_));
 sky130_fd_sc_hd__and2_1 _08857_ (.A(_01682_),
    .B(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__clkbuf_1 _08858_ (.A(_01684_),
    .X(\m1.out[18] ));
 sky130_fd_sc_hd__nor2_1 _08859_ (.A(_01598_),
    .B(_01593_),
    .Y(_01685_));
 sky130_fd_sc_hd__inv_2 _08860_ (.A(_01685_),
    .Y(_01687_));
 sky130_fd_sc_hd__nand2_1 _08861_ (.A(_01645_),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__nand2_1 _08862_ (.A(_01540_),
    .B(_01543_),
    .Y(_01689_));
 sky130_fd_sc_hd__nor2_1 _08863_ (.A(_01543_),
    .B(_01540_),
    .Y(_01690_));
 sky130_fd_sc_hd__a21oi_2 _08864_ (.A1(_01689_),
    .A2(_01590_),
    .B1(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__buf_6 _08865_ (.A(_06175_),
    .X(_01692_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_06270_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__inv_2 _08867_ (.A(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _08868_ (.A(_06327_),
    .B(_06178_),
    .Y(_01695_));
 sky130_fd_sc_hd__nand2_1 _08869_ (.A(_01694_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__inv_2 _08870_ (.A(_01695_),
    .Y(_01698_));
 sky130_fd_sc_hd__nand2_1 _08871_ (.A(_01698_),
    .B(_01693_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _08872_ (.A(_06276_),
    .B(_06172_),
    .Y(_01700_));
 sky130_fd_sc_hd__nand3_1 _08873_ (.A(_01696_),
    .B(_01699_),
    .C(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(_01698_),
    .B(_01694_),
    .Y(_01702_));
 sky130_fd_sc_hd__inv_2 _08875_ (.A(_01700_),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(_01695_),
    .B(_01693_),
    .Y(_01704_));
 sky130_fd_sc_hd__nand3_1 _08877_ (.A(_01702_),
    .B(_01703_),
    .C(_01704_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_1 _08878_ (.A(_01701_),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__a21oi_2 _08879_ (.A1(_01481_),
    .A2(_01486_),
    .B1(_01480_),
    .Y(_01707_));
 sky130_fd_sc_hd__inv_2 _08880_ (.A(_01707_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_1 _08881_ (.A(_01706_),
    .B(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand3_1 _08882_ (.A(_01707_),
    .B(_01701_),
    .C(_01705_),
    .Y(_01711_));
 sky130_fd_sc_hd__nand2_1 _08883_ (.A(_01710_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__nand2_1 _08884_ (.A(_06274_),
    .B(_01278_),
    .Y(_01713_));
 sky130_fd_sc_hd__inv_2 _08885_ (.A(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__nand2_1 _08886_ (.A(_06262_),
    .B(_00918_),
    .Y(_01715_));
 sky130_fd_sc_hd__nand2_1 _08887_ (.A(_01714_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__inv_2 _08888_ (.A(_01715_),
    .Y(_01717_));
 sky130_fd_sc_hd__nand2_1 _08889_ (.A(_01717_),
    .B(_01713_),
    .Y(_01718_));
 sky130_fd_sc_hd__nand2_1 _08890_ (.A(_06259_),
    .B(_06223_),
    .Y(_01720_));
 sky130_fd_sc_hd__nand3_1 _08891_ (.A(_01716_),
    .B(_01718_),
    .C(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__nand2_1 _08892_ (.A(_01717_),
    .B(_01714_),
    .Y(_01722_));
 sky130_fd_sc_hd__inv_2 _08893_ (.A(_01720_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_1 _08894_ (.A(_01715_),
    .B(_01713_),
    .Y(_01724_));
 sky130_fd_sc_hd__nand3_1 _08895_ (.A(_01722_),
    .B(_01723_),
    .C(_01724_),
    .Y(_01725_));
 sky130_fd_sc_hd__nand2_2 _08896_ (.A(_01721_),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__inv_2 _08897_ (.A(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand2_1 _08898_ (.A(_01712_),
    .B(_01727_),
    .Y(_01728_));
 sky130_fd_sc_hd__nand3_1 _08899_ (.A(_01710_),
    .B(_01711_),
    .C(_01726_),
    .Y(_01729_));
 sky130_fd_sc_hd__nand2_1 _08900_ (.A(_01728_),
    .B(_01729_),
    .Y(_01731_));
 sky130_fd_sc_hd__nand2_1 _08901_ (.A(_01488_),
    .B(_01490_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_1 _08902_ (.A(_01490_),
    .B(_01488_),
    .Y(_01733_));
 sky130_fd_sc_hd__a21oi_2 _08903_ (.A1(_01732_),
    .A2(_01507_),
    .B1(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__or2_1 _08904_ (.A(_01731_),
    .B(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__nand2_2 _08905_ (.A(_06265_),
    .B(_06217_),
    .Y(_01736_));
 sky130_fd_sc_hd__inv_2 _08906_ (.A(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_1 _08907_ (.A(_00299_),
    .B(_06220_),
    .Y(_01738_));
 sky130_fd_sc_hd__nand2_1 _08908_ (.A(_01737_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__inv_2 _08909_ (.A(_01738_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand2_1 _08910_ (.A(_01740_),
    .B(_01736_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand2_1 _08911_ (.A(_00193_),
    .B(_00376_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand3_1 _08912_ (.A(_01739_),
    .B(_01742_),
    .C(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__nand2_1 _08913_ (.A(_01740_),
    .B(_01737_),
    .Y(_01745_));
 sky130_fd_sc_hd__inv_2 _08914_ (.A(_01743_),
    .Y(_01746_));
 sky130_fd_sc_hd__nand2_1 _08915_ (.A(_01738_),
    .B(_01736_),
    .Y(_01747_));
 sky130_fd_sc_hd__nand3_2 _08916_ (.A(_01745_),
    .B(_01746_),
    .C(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nand2_1 _08917_ (.A(_01744_),
    .B(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__a21oi_2 _08918_ (.A1(_01497_),
    .A2(_01502_),
    .B1(_01496_),
    .Y(_01750_));
 sky130_fd_sc_hd__inv_2 _08919_ (.A(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_1 _08920_ (.A(_01749_),
    .B(_01751_),
    .Y(_01753_));
 sky130_fd_sc_hd__nand3_1 _08921_ (.A(_01750_),
    .B(_01744_),
    .C(_01748_),
    .Y(_01754_));
 sky130_fd_sc_hd__nand2_1 _08922_ (.A(_01753_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__a21o_1 _08923_ (.A1(_01520_),
    .A2(_01525_),
    .B1(_01519_),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_1 _08924_ (.A(_01755_),
    .B(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand3b_1 _08925_ (.A_N(_01756_),
    .B(_01753_),
    .C(_01754_),
    .Y(_01758_));
 sky130_fd_sc_hd__nand2_1 _08926_ (.A(_01757_),
    .B(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__inv_2 _08927_ (.A(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__nand2_1 _08928_ (.A(_01734_),
    .B(_01731_),
    .Y(_01761_));
 sky130_fd_sc_hd__nand3_1 _08929_ (.A(_01735_),
    .B(_01760_),
    .C(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2b_1 _08930_ (.A_N(_01734_),
    .B(_01731_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand3_1 _08931_ (.A(_01734_),
    .B(_01729_),
    .C(_01728_),
    .Y(_01765_));
 sky130_fd_sc_hd__nand3_1 _08932_ (.A(_01764_),
    .B(_01759_),
    .C(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__nand2_1 _08933_ (.A(_01762_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__nand2_1 _08934_ (.A(_01510_),
    .B(_01476_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _08935_ (.A(_01476_),
    .B(_01510_),
    .Y(_01769_));
 sky130_fd_sc_hd__a21o_1 _08936_ (.A1(_01768_),
    .A2(_01537_),
    .B1(_01769_),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_1 _08937_ (.A(_01767_),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__a21oi_2 _08938_ (.A1(_01768_),
    .A2(_01537_),
    .B1(_01769_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand3_1 _08939_ (.A(_01772_),
    .B(_01762_),
    .C(_01766_),
    .Y(_01773_));
 sky130_fd_sc_hd__nor2_1 _08940_ (.A(_01527_),
    .B(_01516_),
    .Y(_01775_));
 sky130_fd_sc_hd__a21oi_2 _08941_ (.A1(_01528_),
    .A2(_01531_),
    .B1(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__nand2_1 _08942_ (.A(_00439_),
    .B(_00780_),
    .Y(_01777_));
 sky130_fd_sc_hd__nand2_1 _08943_ (.A(_06286_),
    .B(_06230_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _08944_ (.A(_01777_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__nand2_1 _08945_ (.A(_01777_),
    .B(_01778_),
    .Y(_01780_));
 sky130_fd_sc_hd__inv_2 _08946_ (.A(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _08947_ (.A(net3),
    .B(net63),
    .Y(_01782_));
 sky130_fd_sc_hd__o21ai_1 _08948_ (.A1(_01779_),
    .A2(_01781_),
    .B1(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__inv_2 _08949_ (.A(_01782_),
    .Y(_01784_));
 sky130_fd_sc_hd__nand3b_1 _08950_ (.A_N(_01779_),
    .B(_01784_),
    .C(_01780_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _08951_ (.A(_01783_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__a21oi_2 _08952_ (.A1(_01554_),
    .A2(_01559_),
    .B1(_01553_),
    .Y(_01788_));
 sky130_fd_sc_hd__inv_2 _08953_ (.A(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _08954_ (.A(_01787_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__nand3_1 _08955_ (.A(_01783_),
    .B(_01786_),
    .C(_01788_),
    .Y(_01791_));
 sky130_fd_sc_hd__nand2_1 _08956_ (.A(_06278_),
    .B(_06201_),
    .Y(_01792_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(net4),
    .B(_06199_),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _08958_ (.A(_01792_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__nand2_1 _08959_ (.A(_01792_),
    .B(_01793_),
    .Y(_01795_));
 sky130_fd_sc_hd__inv_2 _08960_ (.A(_01795_),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_1 _08961_ (.A(_06283_),
    .B(_06195_),
    .Y(_01798_));
 sky130_fd_sc_hd__o21ai_1 _08962_ (.A1(_01794_),
    .A2(_01797_),
    .B1(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__inv_2 _08963_ (.A(_01798_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand3b_1 _08964_ (.A_N(_01794_),
    .B(_01800_),
    .C(_01795_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _08965_ (.A(_01799_),
    .B(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__nand3_1 _08966_ (.A(_01790_),
    .B(_01791_),
    .C(_01802_),
    .Y(_01803_));
 sky130_fd_sc_hd__nand2_1 _08967_ (.A(_01787_),
    .B(_01788_),
    .Y(_01804_));
 sky130_fd_sc_hd__nand3_1 _08968_ (.A(_01783_),
    .B(_01786_),
    .C(_01789_),
    .Y(_01805_));
 sky130_fd_sc_hd__inv_2 _08969_ (.A(_01802_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand3_1 _08970_ (.A(_01804_),
    .B(_01805_),
    .C(_01806_),
    .Y(_01808_));
 sky130_fd_sc_hd__nand3_1 _08971_ (.A(_01776_),
    .B(_01803_),
    .C(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__inv_2 _08972_ (.A(_01776_),
    .Y(_01810_));
 sky130_fd_sc_hd__nand2_1 _08973_ (.A(_01808_),
    .B(_01803_),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(_01810_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__nand2_1 _08975_ (.A(_01809_),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__nand2_1 _08976_ (.A(_01578_),
    .B(_01563_),
    .Y(_01814_));
 sky130_fd_sc_hd__nand2_1 _08977_ (.A(_01813_),
    .B(_01814_),
    .Y(_01815_));
 sky130_fd_sc_hd__nand3b_1 _08978_ (.A_N(_01814_),
    .B(_01809_),
    .C(_01812_),
    .Y(_01816_));
 sky130_fd_sc_hd__nand2_2 _08979_ (.A(_01815_),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__nand3_1 _08980_ (.A(_01771_),
    .B(_01773_),
    .C(_01817_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand3_1 _08981_ (.A(_01770_),
    .B(_01766_),
    .C(_01762_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2_1 _08982_ (.A(_01767_),
    .B(_01772_),
    .Y(_01821_));
 sky130_fd_sc_hd__inv_2 _08983_ (.A(_01817_),
    .Y(_01822_));
 sky130_fd_sc_hd__nand3_1 _08984_ (.A(_01820_),
    .B(_01821_),
    .C(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__nand3_1 _08985_ (.A(_01691_),
    .B(_01819_),
    .C(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand2_1 _08986_ (.A(_01823_),
    .B(_01819_),
    .Y(_01825_));
 sky130_fd_sc_hd__a21o_1 _08987_ (.A1(_01689_),
    .A2(_01590_),
    .B1(_01690_),
    .X(_01826_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(_01825_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__a21boi_1 _08989_ (.A1(_01619_),
    .A2(_01616_),
    .B1_N(_01617_),
    .Y(_01828_));
 sky130_fd_sc_hd__nand2_1 _08990_ (.A(_01211_),
    .B(_06211_),
    .Y(_01830_));
 sky130_fd_sc_hd__clkbuf_8 _08991_ (.A(_06281_),
    .X(_01831_));
 sky130_fd_sc_hd__nand2_1 _08992_ (.A(_01831_),
    .B(_06198_),
    .Y(_01832_));
 sky130_fd_sc_hd__nor2_1 _08993_ (.A(_01830_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_1 _08994_ (.A(_01830_),
    .B(_01832_),
    .Y(_01834_));
 sky130_fd_sc_hd__inv_2 _08995_ (.A(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__nand2_1 _08996_ (.A(_06234_),
    .B(_06213_),
    .Y(_01836_));
 sky130_fd_sc_hd__o21ai_1 _08997_ (.A1(_01833_),
    .A2(_01835_),
    .B1(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__nor2_1 _08998_ (.A(_01833_),
    .B(_01835_),
    .Y(_01838_));
 sky130_fd_sc_hd__inv_2 _08999_ (.A(_01836_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand2_1 _09000_ (.A(_01838_),
    .B(_01839_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _09001_ (.A(_01837_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__a21oi_2 _09002_ (.A1(_01569_),
    .A2(_01573_),
    .B1(_01568_),
    .Y(_01843_));
 sky130_fd_sc_hd__nand2_1 _09003_ (.A(_01842_),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__inv_2 _09004_ (.A(_01843_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand3_1 _09005_ (.A(_01837_),
    .B(_01845_),
    .C(_01841_),
    .Y(_01846_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(_01844_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__a21oi_1 _09007_ (.A1(_01608_),
    .A2(_01613_),
    .B1(_01607_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _09008_ (.A(_01847_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__inv_2 _09009_ (.A(_01848_),
    .Y(_01850_));
 sky130_fd_sc_hd__nand3_1 _09010_ (.A(_01844_),
    .B(_01846_),
    .C(_01850_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand3_1 _09011_ (.A(_01828_),
    .B(_01849_),
    .C(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_1 _09012_ (.A(_01623_),
    .B(_01617_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand2_1 _09013_ (.A(_01849_),
    .B(_01852_),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _09014_ (.A(_01854_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_01853_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__buf_4 _09016_ (.A(net11),
    .X(_01858_));
 sky130_fd_sc_hd__and4_1 _09017_ (.A(_01858_),
    .B(_06242_),
    .C(_06204_),
    .D(_06207_),
    .X(_01859_));
 sky130_fd_sc_hd__inv_2 _09018_ (.A(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__a22o_1 _09019_ (.A1(_06240_),
    .A2(_06209_),
    .B1(_06243_),
    .B2(_06206_),
    .X(_01861_));
 sky130_fd_sc_hd__and2_1 _09020_ (.A(_01860_),
    .B(_01861_),
    .X(_01863_));
 sky130_fd_sc_hd__nand2_1 _09021_ (.A(_01857_),
    .B(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__nand3b_1 _09022_ (.A_N(_01863_),
    .B(_01853_),
    .C(_01856_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _09023_ (.A(_01864_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand2_1 _09024_ (.A(_01579_),
    .B(_01580_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor2_1 _09025_ (.A(_01580_),
    .B(_01579_),
    .Y(_01868_));
 sky130_fd_sc_hd__a21oi_2 _09026_ (.A1(_01867_),
    .A2(_01585_),
    .B1(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__inv_2 _09027_ (.A(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hd__nand2_1 _09028_ (.A(_01866_),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__nand3_1 _09029_ (.A(_01869_),
    .B(_01864_),
    .C(_01865_),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_1 _09030_ (.A(_01871_),
    .B(_01872_),
    .Y(_01874_));
 sky130_fd_sc_hd__nand2_1 _09031_ (.A(_01633_),
    .B(_01624_),
    .Y(_01875_));
 sky130_fd_sc_hd__nand2_1 _09032_ (.A(_01874_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__inv_2 _09033_ (.A(_01875_),
    .Y(_01877_));
 sky130_fd_sc_hd__nand3_1 _09034_ (.A(_01871_),
    .B(_01872_),
    .C(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _09035_ (.A(_01876_),
    .B(_01878_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand3_1 _09036_ (.A(_01824_),
    .B(_01827_),
    .C(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _09037_ (.A(_01824_),
    .B(_01827_),
    .Y(_01881_));
 sky130_fd_sc_hd__inv_2 _09038_ (.A(_01879_),
    .Y(_01882_));
 sky130_fd_sc_hd__nand2_1 _09039_ (.A(_01881_),
    .B(_01882_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand3_1 _09040_ (.A(_01688_),
    .B(_01880_),
    .C(_01883_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_1 _09041_ (.A(_01883_),
    .B(_01880_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _09042_ (.A(_01593_),
    .B(_01598_),
    .Y(_01887_));
 sky130_fd_sc_hd__a21oi_1 _09043_ (.A1(_01644_),
    .A2(_01887_),
    .B1(_01685_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_1 _09044_ (.A(_01886_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__nand2_1 _09045_ (.A(_01641_),
    .B(_01638_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand3_2 _09046_ (.A(_01885_),
    .B(_01889_),
    .C(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__nand3_1 _09047_ (.A(_01888_),
    .B(_01880_),
    .C(_01883_),
    .Y(_01892_));
 sky130_fd_sc_hd__nand2_1 _09048_ (.A(_01886_),
    .B(_01688_),
    .Y(_01893_));
 sky130_fd_sc_hd__inv_2 _09049_ (.A(_01890_),
    .Y(_01894_));
 sky130_fd_sc_hd__nand3_1 _09050_ (.A(_01892_),
    .B(_01893_),
    .C(_01894_),
    .Y(_01896_));
 sky130_fd_sc_hd__nand2_1 _09051_ (.A(_01891_),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_1 _09052_ (.A(_01647_),
    .B(_01650_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _09053_ (.A(_01650_),
    .B(_01647_),
    .Y(_01899_));
 sky130_fd_sc_hd__a21oi_1 _09054_ (.A1(_01898_),
    .A2(_01656_),
    .B1(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hd__inv_2 _09055_ (.A(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _09056_ (.A(_01897_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__nand3_1 _09057_ (.A(_01900_),
    .B(_01891_),
    .C(_01896_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _09058_ (.A(_01902_),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__inv_2 _09059_ (.A(_01670_),
    .Y(_01905_));
 sky130_fd_sc_hd__nand2_1 _09060_ (.A(_01904_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__nand3_1 _09061_ (.A(_01902_),
    .B(_01903_),
    .C(_01670_),
    .Y(_01907_));
 sky130_fd_sc_hd__nand2_1 _09062_ (.A(_01906_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__nand2_1 _09063_ (.A(_01683_),
    .B(_01674_),
    .Y(_01909_));
 sky130_fd_sc_hd__xnor2_1 _09064_ (.A(_01908_),
    .B(_01909_),
    .Y(\m1.out[19] ));
 sky130_fd_sc_hd__nand2b_1 _09065_ (.A_N(_01897_),
    .B(_01901_),
    .Y(_01910_));
 sky130_fd_sc_hd__a21boi_1 _09066_ (.A1(_01890_),
    .A2(_01889_),
    .B1_N(_01885_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand2_1 _09067_ (.A(_01825_),
    .B(_01691_),
    .Y(_01912_));
 sky130_fd_sc_hd__nor2_1 _09068_ (.A(_01691_),
    .B(_01825_),
    .Y(_01913_));
 sky130_fd_sc_hd__a21oi_1 _09069_ (.A1(_01882_),
    .A2(_01912_),
    .B1(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _09070_ (.A(_01772_),
    .B(_01767_),
    .Y(_01916_));
 sky130_fd_sc_hd__a21oi_1 _09071_ (.A1(_01821_),
    .A2(_01822_),
    .B1(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _09072_ (.A(_01706_),
    .B(_01707_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _09073_ (.A(_01707_),
    .B(_01706_),
    .Y(_01919_));
 sky130_fd_sc_hd__a21oi_1 _09074_ (.A1(_01918_),
    .A2(_01727_),
    .B1(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__buf_6 _09075_ (.A(_06187_),
    .X(_01921_));
 sky130_fd_sc_hd__buf_6 _09076_ (.A(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__nand2_1 _09077_ (.A(_06271_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__inv_2 _09078_ (.A(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _09079_ (.A(_06327_),
    .B(_01692_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_1 _09080_ (.A(_01924_),
    .B(_01925_),
    .Y(_01927_));
 sky130_fd_sc_hd__inv_2 _09081_ (.A(_01925_),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _09082_ (.A(_01928_),
    .B(_01923_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_1 _09083_ (.A(_06276_),
    .B(_06178_),
    .Y(_01930_));
 sky130_fd_sc_hd__nand3_1 _09084_ (.A(_01927_),
    .B(_01929_),
    .C(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__nand2_1 _09085_ (.A(_01928_),
    .B(_01924_),
    .Y(_01932_));
 sky130_fd_sc_hd__inv_2 _09086_ (.A(_01930_),
    .Y(_01933_));
 sky130_fd_sc_hd__nand2_1 _09087_ (.A(_01925_),
    .B(_01923_),
    .Y(_01934_));
 sky130_fd_sc_hd__nand3_1 _09088_ (.A(_01932_),
    .B(_01933_),
    .C(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__nand2_1 _09089_ (.A(_01931_),
    .B(_01935_),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _09090_ (.A(_01695_),
    .B(_01693_),
    .Y(_01938_));
 sky130_fd_sc_hd__a21o_1 _09091_ (.A1(_01704_),
    .A2(_01703_),
    .B1(_01938_),
    .X(_01939_));
 sky130_fd_sc_hd__nand2_1 _09092_ (.A(_01936_),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__a21oi_1 _09093_ (.A1(_01704_),
    .A2(_01703_),
    .B1(_01938_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand3_1 _09094_ (.A(_01941_),
    .B(_01931_),
    .C(_01935_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _09095_ (.A(_06261_),
    .B(_01278_),
    .Y(_01943_));
 sky130_fd_sc_hd__inv_2 _09096_ (.A(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__nand2_1 _09097_ (.A(_06273_),
    .B(_06171_),
    .Y(_01945_));
 sky130_fd_sc_hd__inv_2 _09098_ (.A(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__nand2_1 _09099_ (.A(_01944_),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__nand2_1 _09100_ (.A(_01943_),
    .B(_01945_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_1 _09101_ (.A(_01947_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__nand2_1 _09102_ (.A(_06258_),
    .B(net39),
    .Y(_01951_));
 sky130_fd_sc_hd__nand2_1 _09103_ (.A(_01950_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__inv_2 _09104_ (.A(_01951_),
    .Y(_01953_));
 sky130_fd_sc_hd__nand3_1 _09105_ (.A(_01947_),
    .B(_01953_),
    .C(_01949_),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_2 _09106_ (.A(_01952_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand3_1 _09107_ (.A(_01940_),
    .B(_01942_),
    .C(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__nand3_1 _09108_ (.A(_01939_),
    .B(_01931_),
    .C(_01935_),
    .Y(_01957_));
 sky130_fd_sc_hd__nand2_1 _09109_ (.A(_01936_),
    .B(_01941_),
    .Y(_01958_));
 sky130_fd_sc_hd__inv_2 _09110_ (.A(_01955_),
    .Y(_01960_));
 sky130_fd_sc_hd__nand3_1 _09111_ (.A(_01957_),
    .B(_01958_),
    .C(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand3_1 _09112_ (.A(_01920_),
    .B(_01956_),
    .C(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__a21o_1 _09113_ (.A1(_01918_),
    .A2(_01727_),
    .B1(_01919_),
    .X(_01963_));
 sky130_fd_sc_hd__nand2_1 _09114_ (.A(_01961_),
    .B(_01956_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _09115_ (.A(_01963_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__nand2_1 _09116_ (.A(_01962_),
    .B(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _09117_ (.A(_00299_),
    .B(_00926_),
    .Y(_01967_));
 sky130_fd_sc_hd__inv_2 _09118_ (.A(_01967_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _09119_ (.A(_06266_),
    .B(_00921_),
    .Y(_01969_));
 sky130_fd_sc_hd__inv_2 _09120_ (.A(_01969_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand2_1 _09121_ (.A(_01968_),
    .B(_01971_),
    .Y(_01972_));
 sky130_fd_sc_hd__nand2_1 _09122_ (.A(_01967_),
    .B(_01969_),
    .Y(_01973_));
 sky130_fd_sc_hd__nand2_1 _09123_ (.A(_01972_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__nand2_1 _09124_ (.A(_06290_),
    .B(_06220_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _09125_ (.A(_01974_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__inv_2 _09126_ (.A(_01975_),
    .Y(_01977_));
 sky130_fd_sc_hd__nand3_2 _09127_ (.A(_01972_),
    .B(_01977_),
    .C(_01973_),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(_01976_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _09129_ (.A(_01715_),
    .B(_01713_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21oi_1 _09130_ (.A1(_01724_),
    .A2(_01723_),
    .B1(_01980_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand2_1 _09131_ (.A(_01979_),
    .B(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hd__a21o_1 _09132_ (.A1(_01724_),
    .A2(_01723_),
    .B1(_01980_),
    .X(_01984_));
 sky130_fd_sc_hd__nand3_1 _09133_ (.A(_01984_),
    .B(_01976_),
    .C(_01978_),
    .Y(_01985_));
 sky130_fd_sc_hd__nand2_1 _09134_ (.A(_01748_),
    .B(_01745_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand3_1 _09135_ (.A(_01983_),
    .B(_01985_),
    .C(_01986_),
    .Y(_01987_));
 sky130_fd_sc_hd__nand2_1 _09136_ (.A(_01979_),
    .B(_01984_),
    .Y(_01988_));
 sky130_fd_sc_hd__nand3_1 _09137_ (.A(_01976_),
    .B(_01982_),
    .C(_01978_),
    .Y(_01989_));
 sky130_fd_sc_hd__inv_2 _09138_ (.A(_01986_),
    .Y(_01990_));
 sky130_fd_sc_hd__nand3_1 _09139_ (.A(_01988_),
    .B(_01989_),
    .C(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_2 _09140_ (.A(_01987_),
    .B(_01991_),
    .Y(_01993_));
 sky130_fd_sc_hd__inv_2 _09141_ (.A(_01993_),
    .Y(_01994_));
 sky130_fd_sc_hd__nand2_1 _09142_ (.A(_01966_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__nand3_1 _09143_ (.A(_01962_),
    .B(_01965_),
    .C(_01993_),
    .Y(_01996_));
 sky130_fd_sc_hd__nand2_2 _09144_ (.A(_01995_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__inv_2 _09145_ (.A(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__nor2_1 _09146_ (.A(_01731_),
    .B(_01734_),
    .Y(_01999_));
 sky130_fd_sc_hd__a21oi_2 _09147_ (.A1(_01761_),
    .A2(_01760_),
    .B1(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__nand2_1 _09148_ (.A(_01998_),
    .B(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__inv_2 _09149_ (.A(_02000_),
    .Y(_02002_));
 sky130_fd_sc_hd__nand2_1 _09150_ (.A(_02002_),
    .B(_01997_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand2_1 _09151_ (.A(_01808_),
    .B(_01805_),
    .Y(_02005_));
 sky130_fd_sc_hd__nand2_2 _09152_ (.A(_06286_),
    .B(_06227_),
    .Y(_02006_));
 sky130_fd_sc_hd__inv_2 _09153_ (.A(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_2 _09154_ (.A(net2),
    .B(_06229_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2_1 _09155_ (.A(_02007_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__inv_2 _09156_ (.A(_02008_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _09157_ (.A(_02010_),
    .B(_02006_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2_1 _09158_ (.A(_00561_),
    .B(_00780_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand3_1 _09159_ (.A(_02009_),
    .B(_02011_),
    .C(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_1 _09160_ (.A(_02010_),
    .B(_02007_),
    .Y(_02015_));
 sky130_fd_sc_hd__inv_2 _09161_ (.A(_02012_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_1 _09162_ (.A(_02008_),
    .B(_02006_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand3_1 _09163_ (.A(_02015_),
    .B(_02016_),
    .C(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__nand2_1 _09164_ (.A(_02013_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__a21oi_2 _09165_ (.A1(_01780_),
    .A2(_01784_),
    .B1(_01779_),
    .Y(_02020_));
 sky130_fd_sc_hd__inv_2 _09166_ (.A(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__nand2_1 _09167_ (.A(_02019_),
    .B(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__nand3_1 _09168_ (.A(_02020_),
    .B(_02013_),
    .C(_02018_),
    .Y(_02023_));
 sky130_fd_sc_hd__nand2_1 _09169_ (.A(_02022_),
    .B(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_1 _09170_ (.A(_06278_),
    .B(net62),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _09171_ (.A(net4),
    .B(net63),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _09172_ (.A(_02026_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__inv_2 _09173_ (.A(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__nand2_1 _09174_ (.A(_02026_),
    .B(_02027_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand2_1 _09175_ (.A(_02029_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__nand2_1 _09176_ (.A(_06283_),
    .B(_06201_),
    .Y(_02032_));
 sky130_fd_sc_hd__nand2_1 _09177_ (.A(_02031_),
    .B(_02032_),
    .Y(_02033_));
 sky130_fd_sc_hd__inv_2 _09178_ (.A(_02032_),
    .Y(_02034_));
 sky130_fd_sc_hd__nand3_1 _09179_ (.A(_02029_),
    .B(_02034_),
    .C(_02030_),
    .Y(_02035_));
 sky130_fd_sc_hd__nand2_1 _09180_ (.A(_02033_),
    .B(_02035_),
    .Y(_02037_));
 sky130_fd_sc_hd__inv_2 _09181_ (.A(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _09182_ (.A(_02024_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand3_1 _09183_ (.A(_02022_),
    .B(_02023_),
    .C(_02037_),
    .Y(_02040_));
 sky130_fd_sc_hd__nand2_1 _09184_ (.A(_02039_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _09185_ (.A(_01749_),
    .B(_01750_),
    .Y(_02042_));
 sky130_fd_sc_hd__nor2_1 _09186_ (.A(_01750_),
    .B(_01749_),
    .Y(_02043_));
 sky130_fd_sc_hd__a21o_1 _09187_ (.A1(_02042_),
    .A2(_01756_),
    .B1(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__nand2_1 _09188_ (.A(_02041_),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__a21oi_1 _09189_ (.A1(_02042_),
    .A2(_01756_),
    .B1(_02043_),
    .Y(_02046_));
 sky130_fd_sc_hd__nand3_1 _09190_ (.A(_02046_),
    .B(_02040_),
    .C(_02039_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand3b_1 _09191_ (.A_N(_02005_),
    .B(_02045_),
    .C(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__nand2_1 _09192_ (.A(_02048_),
    .B(_02045_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_1 _09193_ (.A(_02050_),
    .B(_02005_),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_02049_),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__nand3_1 _09195_ (.A(_02001_),
    .B(_02004_),
    .C(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_1 _09196_ (.A(_01998_),
    .B(_02002_),
    .Y(_02054_));
 sky130_fd_sc_hd__inv_2 _09197_ (.A(_02052_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _09198_ (.A(_01997_),
    .B(_02000_),
    .Y(_02056_));
 sky130_fd_sc_hd__nand3_1 _09199_ (.A(_02054_),
    .B(_02055_),
    .C(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand3_1 _09200_ (.A(_01917_),
    .B(_02053_),
    .C(_02057_),
    .Y(_02059_));
 sky130_fd_sc_hd__nand2_1 _09201_ (.A(_01823_),
    .B(_01820_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand2_1 _09202_ (.A(_02057_),
    .B(_02053_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _09203_ (.A(_02060_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _09204_ (.A(_01843_),
    .B(_01842_),
    .Y(_02063_));
 sky130_fd_sc_hd__a21oi_1 _09205_ (.A1(_01844_),
    .A2(_01850_),
    .B1(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__a21oi_2 _09206_ (.A1(_01795_),
    .A2(_01800_),
    .B1(_01794_),
    .Y(_02065_));
 sky130_fd_sc_hd__inv_2 _09207_ (.A(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand2_1 _09208_ (.A(_06237_),
    .B(_06197_),
    .Y(_02067_));
 sky130_fd_sc_hd__inv_2 _09209_ (.A(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _09210_ (.A(_06281_),
    .B(_06195_),
    .Y(_02070_));
 sky130_fd_sc_hd__nand2_1 _09211_ (.A(_02068_),
    .B(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__inv_2 _09212_ (.A(_02070_),
    .Y(_02072_));
 sky130_fd_sc_hd__nand2_1 _09213_ (.A(_02072_),
    .B(_02067_),
    .Y(_02073_));
 sky130_fd_sc_hd__nand2_1 _09214_ (.A(_06234_),
    .B(_06210_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand3_1 _09215_ (.A(_02071_),
    .B(_02073_),
    .C(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_1 _09216_ (.A(_02068_),
    .B(_02072_),
    .Y(_02076_));
 sky130_fd_sc_hd__inv_2 _09217_ (.A(_02074_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(_02067_),
    .B(_02070_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand3_1 _09219_ (.A(_02076_),
    .B(_02077_),
    .C(_02078_),
    .Y(_02079_));
 sky130_fd_sc_hd__nand3_1 _09220_ (.A(_02066_),
    .B(_02075_),
    .C(_02079_),
    .Y(_02081_));
 sky130_fd_sc_hd__nand2_1 _09221_ (.A(_02075_),
    .B(_02079_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _09222_ (.A(_02082_),
    .B(_02065_),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _09223_ (.A(_02081_),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__a21oi_1 _09224_ (.A1(_01834_),
    .A2(_01839_),
    .B1(_01833_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand2_1 _09225_ (.A(_02084_),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__inv_2 _09226_ (.A(_02085_),
    .Y(_02087_));
 sky130_fd_sc_hd__nand3_1 _09227_ (.A(_02081_),
    .B(_02083_),
    .C(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand3_1 _09228_ (.A(_02064_),
    .B(_02086_),
    .C(_02088_),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_1 _09229_ (.A(_01852_),
    .B(_01846_),
    .Y(_02090_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(_02086_),
    .B(_02088_),
    .Y(_02092_));
 sky130_fd_sc_hd__nand2_1 _09231_ (.A(_02090_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__nand2_1 _09232_ (.A(_02089_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__buf_6 _09233_ (.A(net13),
    .X(_02095_));
 sky130_fd_sc_hd__nand2_1 _09234_ (.A(_02095_),
    .B(net33),
    .Y(_02096_));
 sky130_fd_sc_hd__nand2_1 _09235_ (.A(_06239_),
    .B(net44),
    .Y(_02097_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(_06241_),
    .B(_06213_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_1 _09237_ (.A(_02097_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__nand2_1 _09238_ (.A(_02097_),
    .B(_02098_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2b_1 _09239_ (.A(_02099_),
    .B_N(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__xor2_1 _09240_ (.A(_02096_),
    .B(_02101_),
    .X(_02103_));
 sky130_fd_sc_hd__or2_1 _09241_ (.A(_01860_),
    .B(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__nand2_1 _09242_ (.A(_02103_),
    .B(_01860_),
    .Y(_02105_));
 sky130_fd_sc_hd__nand2_1 _09243_ (.A(_02104_),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__inv_2 _09244_ (.A(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand2_1 _09245_ (.A(_02094_),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__nand3_1 _09246_ (.A(_02089_),
    .B(_02093_),
    .C(_02106_),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _09247_ (.A(_02108_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__nand2_1 _09248_ (.A(_01811_),
    .B(_01776_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor2_1 _09249_ (.A(_01776_),
    .B(_01811_),
    .Y(_02112_));
 sky130_fd_sc_hd__a21oi_2 _09250_ (.A1(_02111_),
    .A2(_01814_),
    .B1(_02112_),
    .Y(_02114_));
 sky130_fd_sc_hd__inv_2 _09251_ (.A(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _09252_ (.A(_02110_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__nand3_1 _09253_ (.A(_02114_),
    .B(_02108_),
    .C(_02109_),
    .Y(_02117_));
 sky130_fd_sc_hd__nand2_1 _09254_ (.A(_02116_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__nand2_1 _09255_ (.A(_01828_),
    .B(_01855_),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _09256_ (.A(_01855_),
    .B(_01828_),
    .Y(_02120_));
 sky130_fd_sc_hd__a21oi_1 _09257_ (.A1(_02119_),
    .A2(_01863_),
    .B1(_02120_),
    .Y(_02121_));
 sky130_fd_sc_hd__inv_2 _09258_ (.A(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_02118_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand3_1 _09260_ (.A(_02116_),
    .B(_02117_),
    .C(_02121_),
    .Y(_02125_));
 sky130_fd_sc_hd__nand2_1 _09261_ (.A(_02123_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand3_1 _09262_ (.A(_02059_),
    .B(_02062_),
    .C(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__nand2_1 _09263_ (.A(_02059_),
    .B(_02062_),
    .Y(_02128_));
 sky130_fd_sc_hd__inv_2 _09264_ (.A(_02126_),
    .Y(_02129_));
 sky130_fd_sc_hd__nand2_1 _09265_ (.A(_02128_),
    .B(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand3_1 _09266_ (.A(_01914_),
    .B(_02127_),
    .C(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__a21o_1 _09267_ (.A1(_01882_),
    .A2(_01912_),
    .B1(_01913_),
    .X(_02132_));
 sky130_fd_sc_hd__nand2_1 _09268_ (.A(_02130_),
    .B(_02127_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand2_1 _09269_ (.A(_02132_),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__nand2_1 _09270_ (.A(_02131_),
    .B(_02134_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand3_1 _09271_ (.A(_01870_),
    .B(_01865_),
    .C(_01864_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_2 _09272_ (.A(_01876_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__nand2_1 _09273_ (.A(_02136_),
    .B(_02138_),
    .Y(_02139_));
 sky130_fd_sc_hd__inv_2 _09274_ (.A(_02138_),
    .Y(_02140_));
 sky130_fd_sc_hd__nand3_1 _09275_ (.A(_02131_),
    .B(_02134_),
    .C(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nand2_1 _09276_ (.A(_02139_),
    .B(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__nand2_1 _09277_ (.A(_01911_),
    .B(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__nand2_1 _09278_ (.A(_02136_),
    .B(_02140_),
    .Y(_02144_));
 sky130_fd_sc_hd__nand3_1 _09279_ (.A(_02131_),
    .B(_02134_),
    .C(_02138_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand2_1 _09280_ (.A(_02144_),
    .B(_02145_),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_1 _09281_ (.A(_01891_),
    .B(_01885_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand2_1 _09282_ (.A(_02147_),
    .B(_02148_),
    .Y(_02149_));
 sky130_fd_sc_hd__nand2_1 _09283_ (.A(_02143_),
    .B(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hd__nor2_1 _09284_ (.A(_01910_),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__inv_2 _09285_ (.A(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_1 _09286_ (.A(_02150_),
    .B(_01910_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_02152_),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__inv_2 _09288_ (.A(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _09289_ (.A(_01675_),
    .B(_01908_),
    .Y(_02156_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(_01680_),
    .B(_02156_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _09291_ (.A(_01464_),
    .B(_01671_),
    .Y(_02159_));
 sky130_fd_sc_hd__a21boi_1 _09292_ (.A1(_02159_),
    .A2(_01907_),
    .B1_N(_01906_),
    .Y(_02160_));
 sky130_fd_sc_hd__nand2_1 _09293_ (.A(_02158_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__a31o_1 _09294_ (.A1(_01268_),
    .A2(_01678_),
    .A3(_02156_),
    .B1(_02161_),
    .X(_02162_));
 sky130_fd_sc_hd__or2_1 _09295_ (.A(_02155_),
    .B(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__nand2_1 _09296_ (.A(_02162_),
    .B(_02155_),
    .Y(_02164_));
 sky130_fd_sc_hd__and2_1 _09297_ (.A(_02163_),
    .B(_02164_),
    .X(_02165_));
 sky130_fd_sc_hd__clkbuf_1 _09298_ (.A(_02165_),
    .X(\m1.out[20] ));
 sky130_fd_sc_hd__nand2_1 _09299_ (.A(_02133_),
    .B(_01914_),
    .Y(_02166_));
 sky130_fd_sc_hd__nor2_1 _09300_ (.A(_01914_),
    .B(_02133_),
    .Y(_02168_));
 sky130_fd_sc_hd__a21o_1 _09301_ (.A1(_02166_),
    .A2(_02138_),
    .B1(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__or2_1 _09302_ (.A(_02114_),
    .B(_02110_),
    .X(_02170_));
 sky130_fd_sc_hd__and2_1 _09303_ (.A(_02123_),
    .B(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__nor2_1 _09304_ (.A(_02104_),
    .B(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _09305_ (.A(_02171_),
    .B(_02104_),
    .Y(_02173_));
 sky130_fd_sc_hd__nor2b_1 _09306_ (.A(_02172_),
    .B_N(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_1 _09307_ (.A(_02000_),
    .B(_01997_),
    .Y(_02175_));
 sky130_fd_sc_hd__a21oi_1 _09308_ (.A1(_02056_),
    .A2(_02055_),
    .B1(_02175_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _09309_ (.A(_01941_),
    .B(_01936_),
    .Y(_02177_));
 sky130_fd_sc_hd__a21oi_1 _09310_ (.A1(_01958_),
    .A2(_01960_),
    .B1(_02177_),
    .Y(_02179_));
 sky130_fd_sc_hd__buf_6 _09311_ (.A(net46),
    .X(_02180_));
 sky130_fd_sc_hd__buf_6 _09312_ (.A(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__nand2_1 _09313_ (.A(_06270_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__inv_2 _09314_ (.A(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__nand2_2 _09315_ (.A(_06327_),
    .B(_01921_),
    .Y(_02184_));
 sky130_fd_sc_hd__nand2_1 _09316_ (.A(_02183_),
    .B(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hd__inv_2 _09317_ (.A(_02184_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _09318_ (.A(_02186_),
    .B(_02182_),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _09319_ (.A(_06276_),
    .B(_06176_),
    .Y(_02188_));
 sky130_fd_sc_hd__nand3_1 _09320_ (.A(_02185_),
    .B(_02187_),
    .C(_02188_),
    .Y(_02190_));
 sky130_fd_sc_hd__nand2_1 _09321_ (.A(_02186_),
    .B(_02183_),
    .Y(_02191_));
 sky130_fd_sc_hd__inv_2 _09322_ (.A(_02188_),
    .Y(_02192_));
 sky130_fd_sc_hd__nand2_1 _09323_ (.A(_02184_),
    .B(_02182_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand3_1 _09324_ (.A(_02191_),
    .B(_02192_),
    .C(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__nand2_1 _09325_ (.A(_02190_),
    .B(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__nor2_1 _09326_ (.A(_01925_),
    .B(_01923_),
    .Y(_02196_));
 sky130_fd_sc_hd__a21o_1 _09327_ (.A1(_01934_),
    .A2(_01933_),
    .B1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__nand2_1 _09328_ (.A(_02195_),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__a21oi_1 _09329_ (.A1(_01934_),
    .A2(_01933_),
    .B1(_02196_),
    .Y(_02199_));
 sky130_fd_sc_hd__nand3_1 _09330_ (.A(_02199_),
    .B(_02190_),
    .C(_02194_),
    .Y(_02201_));
 sky130_fd_sc_hd__nand2_1 _09331_ (.A(_06274_),
    .B(_06178_),
    .Y(_02202_));
 sky130_fd_sc_hd__inv_2 _09332_ (.A(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2_1 _09333_ (.A(_06262_),
    .B(_06171_),
    .Y(_02204_));
 sky130_fd_sc_hd__nand2_1 _09334_ (.A(_02203_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__inv_2 _09335_ (.A(_02204_),
    .Y(_02206_));
 sky130_fd_sc_hd__nand2_1 _09336_ (.A(_02206_),
    .B(_02202_),
    .Y(_02207_));
 sky130_fd_sc_hd__nand2_1 _09337_ (.A(_06259_),
    .B(_06174_),
    .Y(_02208_));
 sky130_fd_sc_hd__nand3_1 _09338_ (.A(_02205_),
    .B(_02207_),
    .C(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__nand2_1 _09339_ (.A(_02206_),
    .B(_02203_),
    .Y(_02210_));
 sky130_fd_sc_hd__inv_2 _09340_ (.A(_02208_),
    .Y(_02212_));
 sky130_fd_sc_hd__nand2_1 _09341_ (.A(_02204_),
    .B(_02202_),
    .Y(_02213_));
 sky130_fd_sc_hd__nand3_1 _09342_ (.A(_02210_),
    .B(_02212_),
    .C(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hd__nand2_2 _09343_ (.A(_02209_),
    .B(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__nand3_1 _09344_ (.A(_02198_),
    .B(_02201_),
    .C(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__nand3_1 _09345_ (.A(_02197_),
    .B(_02190_),
    .C(_02194_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _09346_ (.A(_02195_),
    .B(_02199_),
    .Y(_02218_));
 sky130_fd_sc_hd__inv_2 _09347_ (.A(_02215_),
    .Y(_02219_));
 sky130_fd_sc_hd__nand3_1 _09348_ (.A(_02217_),
    .B(_02218_),
    .C(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__nand3_1 _09349_ (.A(_02179_),
    .B(_02216_),
    .C(_02220_),
    .Y(_02221_));
 sky130_fd_sc_hd__nand2_1 _09350_ (.A(_02220_),
    .B(_02216_),
    .Y(_02223_));
 sky130_fd_sc_hd__nand2_1 _09351_ (.A(_01961_),
    .B(_01957_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_1 _09352_ (.A(_02223_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hd__nand2_1 _09353_ (.A(_02221_),
    .B(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _09354_ (.A(_06264_),
    .B(_00921_),
    .Y(_02227_));
 sky130_fd_sc_hd__inv_2 _09355_ (.A(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(_06266_),
    .B(_00918_),
    .Y(_02229_));
 sky130_fd_sc_hd__nand2_1 _09357_ (.A(_02228_),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__inv_2 _09358_ (.A(_02229_),
    .Y(_02231_));
 sky130_fd_sc_hd__nand2_1 _09359_ (.A(_02231_),
    .B(_02227_),
    .Y(_02232_));
 sky130_fd_sc_hd__nand2_1 _09360_ (.A(_06290_),
    .B(_00926_),
    .Y(_02233_));
 sky130_fd_sc_hd__nand3_1 _09361_ (.A(_02230_),
    .B(_02232_),
    .C(_02233_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2_1 _09362_ (.A(_02228_),
    .B(_02231_),
    .Y(_02235_));
 sky130_fd_sc_hd__inv_2 _09363_ (.A(_02233_),
    .Y(_02236_));
 sky130_fd_sc_hd__nand2_1 _09364_ (.A(_02227_),
    .B(_02229_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand3_1 _09365_ (.A(_02235_),
    .B(_02236_),
    .C(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(_02234_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _09367_ (.A(_01943_),
    .B(_01945_),
    .Y(_02240_));
 sky130_fd_sc_hd__a21oi_2 _09368_ (.A1(_01949_),
    .A2(_01953_),
    .B1(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__inv_2 _09369_ (.A(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__nand2_1 _09370_ (.A(_02239_),
    .B(_02242_),
    .Y(_02244_));
 sky130_fd_sc_hd__nand3_1 _09371_ (.A(_02241_),
    .B(_02234_),
    .C(_02238_),
    .Y(_02245_));
 sky130_fd_sc_hd__nand2_1 _09372_ (.A(_02244_),
    .B(_02245_),
    .Y(_02246_));
 sky130_fd_sc_hd__nand2_1 _09373_ (.A(_01978_),
    .B(_01972_),
    .Y(_02247_));
 sky130_fd_sc_hd__nand2_1 _09374_ (.A(_02246_),
    .B(_02247_),
    .Y(_02248_));
 sky130_fd_sc_hd__nand3b_1 _09375_ (.A_N(_02247_),
    .B(_02244_),
    .C(_02245_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_2 _09376_ (.A(_02248_),
    .B(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__inv_2 _09377_ (.A(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(_02226_),
    .B(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__nand3_1 _09379_ (.A(_02221_),
    .B(_02225_),
    .C(_02250_),
    .Y(_02253_));
 sky130_fd_sc_hd__nand2_1 _09380_ (.A(_02252_),
    .B(_02253_),
    .Y(_02255_));
 sky130_fd_sc_hd__nand2_1 _09381_ (.A(_01964_),
    .B(_01920_),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_1 _09382_ (.A(_01920_),
    .B(_01964_),
    .Y(_02257_));
 sky130_fd_sc_hd__a21o_1 _09383_ (.A1(_02256_),
    .A2(_01994_),
    .B1(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__nand2_1 _09384_ (.A(_02255_),
    .B(_02258_),
    .Y(_02259_));
 sky130_fd_sc_hd__a21oi_1 _09385_ (.A1(_02256_),
    .A2(_01994_),
    .B1(_02257_),
    .Y(_02260_));
 sky130_fd_sc_hd__nand3_1 _09386_ (.A(_02260_),
    .B(_02252_),
    .C(_02253_),
    .Y(_02261_));
 sky130_fd_sc_hd__nor2_1 _09387_ (.A(_01982_),
    .B(_01979_),
    .Y(_02262_));
 sky130_fd_sc_hd__a21oi_2 _09388_ (.A1(_01983_),
    .A2(_01986_),
    .B1(_02262_),
    .Y(_02263_));
 sky130_fd_sc_hd__nand2_1 _09389_ (.A(_06292_),
    .B(_06228_),
    .Y(_02264_));
 sky130_fd_sc_hd__inv_2 _09390_ (.A(_02264_),
    .Y(_02266_));
 sky130_fd_sc_hd__nand2_1 _09391_ (.A(_06288_),
    .B(_06220_),
    .Y(_02267_));
 sky130_fd_sc_hd__nand2_1 _09392_ (.A(_02266_),
    .B(_02267_),
    .Y(_02268_));
 sky130_fd_sc_hd__inv_2 _09393_ (.A(_02267_),
    .Y(_02269_));
 sky130_fd_sc_hd__nand2_1 _09394_ (.A(_02269_),
    .B(_02264_),
    .Y(_02270_));
 sky130_fd_sc_hd__nand2_1 _09395_ (.A(_06291_),
    .B(_06231_),
    .Y(_02271_));
 sky130_fd_sc_hd__nand3_1 _09396_ (.A(_02268_),
    .B(_02270_),
    .C(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__nand2_1 _09397_ (.A(_02266_),
    .B(_02269_),
    .Y(_02273_));
 sky130_fd_sc_hd__inv_2 _09398_ (.A(_02271_),
    .Y(_02274_));
 sky130_fd_sc_hd__nand2_1 _09399_ (.A(_02264_),
    .B(_02267_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand3_1 _09400_ (.A(_02273_),
    .B(_02274_),
    .C(_02275_),
    .Y(_02277_));
 sky130_fd_sc_hd__nand2_1 _09401_ (.A(_02272_),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__nor2_1 _09402_ (.A(_02008_),
    .B(_02006_),
    .Y(_02279_));
 sky130_fd_sc_hd__a21oi_1 _09403_ (.A1(_02017_),
    .A2(_02016_),
    .B1(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hd__inv_2 _09404_ (.A(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2_1 _09405_ (.A(_02278_),
    .B(_02281_),
    .Y(_02282_));
 sky130_fd_sc_hd__nand3_1 _09406_ (.A(_02280_),
    .B(_02272_),
    .C(_02277_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _09407_ (.A(_00701_),
    .B(_06226_),
    .Y(_02284_));
 sky130_fd_sc_hd__nand2_1 _09408_ (.A(_06280_),
    .B(_00780_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _09409_ (.A(_02284_),
    .B(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__nand2_2 _09410_ (.A(_02284_),
    .B(_02285_),
    .Y(_02288_));
 sky130_fd_sc_hd__inv_2 _09411_ (.A(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _09412_ (.A(_06284_),
    .B(_06200_),
    .Y(_02290_));
 sky130_fd_sc_hd__o21ai_1 _09413_ (.A1(_02286_),
    .A2(_02289_),
    .B1(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__inv_2 _09414_ (.A(_02290_),
    .Y(_02292_));
 sky130_fd_sc_hd__nand3b_1 _09415_ (.A_N(_02286_),
    .B(_02292_),
    .C(_02288_),
    .Y(_02293_));
 sky130_fd_sc_hd__nand2_1 _09416_ (.A(_02291_),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand3_1 _09417_ (.A(_02282_),
    .B(_02283_),
    .C(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__nand2_1 _09418_ (.A(_02282_),
    .B(_02283_),
    .Y(_02296_));
 sky130_fd_sc_hd__inv_2 _09419_ (.A(_02294_),
    .Y(_02297_));
 sky130_fd_sc_hd__nand2_1 _09420_ (.A(_02296_),
    .B(_02297_),
    .Y(_02299_));
 sky130_fd_sc_hd__nand3_1 _09421_ (.A(_02263_),
    .B(_02295_),
    .C(_02299_),
    .Y(_02300_));
 sky130_fd_sc_hd__inv_2 _09422_ (.A(_02263_),
    .Y(_02301_));
 sky130_fd_sc_hd__nand2_1 _09423_ (.A(_02299_),
    .B(_02295_),
    .Y(_02302_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(_02301_),
    .B(_02302_),
    .Y(_02303_));
 sky130_fd_sc_hd__nand2_1 _09425_ (.A(_02300_),
    .B(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__o21ai_2 _09426_ (.A1(_02020_),
    .A2(_02019_),
    .B1(_02039_),
    .Y(_02305_));
 sky130_fd_sc_hd__nand2_1 _09427_ (.A(_02304_),
    .B(_02305_),
    .Y(_02306_));
 sky130_fd_sc_hd__nand3b_1 _09428_ (.A_N(_02305_),
    .B(_02300_),
    .C(_02303_),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_2 _09429_ (.A(_02306_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__nand3_1 _09430_ (.A(_02259_),
    .B(_02261_),
    .C(_02308_),
    .Y(_02310_));
 sky130_fd_sc_hd__nand3_1 _09431_ (.A(_02258_),
    .B(_02253_),
    .C(_02252_),
    .Y(_02311_));
 sky130_fd_sc_hd__nand2_1 _09432_ (.A(_02255_),
    .B(_02260_),
    .Y(_02312_));
 sky130_fd_sc_hd__inv_2 _09433_ (.A(_02308_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand3_1 _09434_ (.A(_02311_),
    .B(_02312_),
    .C(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__nand3_1 _09435_ (.A(_02176_),
    .B(_02310_),
    .C(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__nand2_1 _09436_ (.A(_02314_),
    .B(_02310_),
    .Y(_02316_));
 sky130_fd_sc_hd__a21o_1 _09437_ (.A1(_02056_),
    .A2(_02055_),
    .B1(_02175_),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_1 _09438_ (.A(_02316_),
    .B(_02317_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _09439_ (.A(_02315_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _09440_ (.A(_06237_),
    .B(_06195_),
    .Y(_02321_));
 sky130_fd_sc_hd__inv_2 _09441_ (.A(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__nand2_1 _09442_ (.A(_01831_),
    .B(_06201_),
    .Y(_02323_));
 sky130_fd_sc_hd__inv_2 _09443_ (.A(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_02322_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__nand2_1 _09445_ (.A(_02321_),
    .B(_02323_),
    .Y(_02326_));
 sky130_fd_sc_hd__nand2_1 _09446_ (.A(_02325_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__nand2_1 _09447_ (.A(_06236_),
    .B(_06198_),
    .Y(_02328_));
 sky130_fd_sc_hd__nand2_1 _09448_ (.A(_02327_),
    .B(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand3b_2 _09449_ (.A_N(_02328_),
    .B(_02325_),
    .C(_02326_),
    .Y(_02330_));
 sky130_fd_sc_hd__nand2_1 _09450_ (.A(_02329_),
    .B(_02330_),
    .Y(_02332_));
 sky130_fd_sc_hd__a21oi_2 _09451_ (.A1(_02030_),
    .A2(_02034_),
    .B1(_02028_),
    .Y(_02333_));
 sky130_fd_sc_hd__nand2_1 _09452_ (.A(_02332_),
    .B(_02333_),
    .Y(_02334_));
 sky130_fd_sc_hd__a21o_1 _09453_ (.A1(_02030_),
    .A2(_02034_),
    .B1(_02028_),
    .X(_02335_));
 sky130_fd_sc_hd__nand3_1 _09454_ (.A(_02335_),
    .B(_02330_),
    .C(_02329_),
    .Y(_02336_));
 sky130_fd_sc_hd__nand2_1 _09455_ (.A(_02079_),
    .B(_02076_),
    .Y(_02337_));
 sky130_fd_sc_hd__nand3_2 _09456_ (.A(_02334_),
    .B(_02336_),
    .C(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__nand2_1 _09457_ (.A(_02332_),
    .B(_02335_),
    .Y(_02339_));
 sky130_fd_sc_hd__nand3_1 _09458_ (.A(_02329_),
    .B(_02330_),
    .C(_02333_),
    .Y(_02340_));
 sky130_fd_sc_hd__inv_2 _09459_ (.A(_02337_),
    .Y(_02341_));
 sky130_fd_sc_hd__nand3_1 _09460_ (.A(_02339_),
    .B(_02340_),
    .C(_02341_),
    .Y(_02343_));
 sky130_fd_sc_hd__nand2_1 _09461_ (.A(_02338_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__nor2_1 _09462_ (.A(_02065_),
    .B(_02082_),
    .Y(_02345_));
 sky130_fd_sc_hd__a21oi_1 _09463_ (.A1(_02083_),
    .A2(_02087_),
    .B1(_02345_),
    .Y(_02346_));
 sky130_fd_sc_hd__inv_2 _09464_ (.A(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _09465_ (.A(_02344_),
    .B(_02347_),
    .Y(_02348_));
 sky130_fd_sc_hd__nand3_1 _09466_ (.A(_02346_),
    .B(_02343_),
    .C(_02338_),
    .Y(_02349_));
 sky130_fd_sc_hd__nand2_1 _09467_ (.A(_02348_),
    .B(_02349_),
    .Y(_02350_));
 sky130_fd_sc_hd__inv_2 _09468_ (.A(_02096_),
    .Y(_02351_));
 sky130_fd_sc_hd__a21oi_1 _09469_ (.A1(_02100_),
    .A2(_02351_),
    .B1(_02099_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _09470_ (.A(_06239_),
    .B(_06213_),
    .Y(_02354_));
 sky130_fd_sc_hd__inv_2 _09471_ (.A(_02354_),
    .Y(_02355_));
 sky130_fd_sc_hd__nand3_2 _09472_ (.A(_02355_),
    .B(_06243_),
    .C(_06212_),
    .Y(_02356_));
 sky130_fd_sc_hd__nand2_1 _09473_ (.A(_06242_),
    .B(_06212_),
    .Y(_02357_));
 sky130_fd_sc_hd__nand2_1 _09474_ (.A(_02354_),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__nand2_1 _09475_ (.A(_02356_),
    .B(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _09476_ (.A(_02095_),
    .B(_06204_),
    .Y(_02360_));
 sky130_fd_sc_hd__nand2_1 _09477_ (.A(_02359_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__inv_2 _09478_ (.A(_02360_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand3_2 _09479_ (.A(_02356_),
    .B(_02362_),
    .C(_02358_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand3b_1 _09480_ (.A_N(_02352_),
    .B(_02361_),
    .C(_02363_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _09481_ (.A(_02361_),
    .B(_02363_),
    .Y(_02366_));
 sky130_fd_sc_hd__nand2_1 _09482_ (.A(_02366_),
    .B(_02352_),
    .Y(_02367_));
 sky130_fd_sc_hd__nand2_1 _09483_ (.A(_02365_),
    .B(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__nand2_1 _09484_ (.A(_06247_),
    .B(_06208_),
    .Y(_02369_));
 sky130_fd_sc_hd__nand2_1 _09485_ (.A(_02368_),
    .B(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__nand3b_1 _09486_ (.A_N(_02369_),
    .B(_02365_),
    .C(_02367_),
    .Y(_02371_));
 sky130_fd_sc_hd__nand2_1 _09487_ (.A(_02370_),
    .B(_02371_),
    .Y(_02372_));
 sky130_fd_sc_hd__inv_2 _09488_ (.A(_02372_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_1 _09489_ (.A(_02350_),
    .B(_02373_),
    .Y(_02374_));
 sky130_fd_sc_hd__nand3_1 _09490_ (.A(_02348_),
    .B(_02349_),
    .C(_02372_),
    .Y(_02376_));
 sky130_fd_sc_hd__nand2_1 _09491_ (.A(_02374_),
    .B(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_1 _09492_ (.A(_02041_),
    .B(_02046_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _09493_ (.A(_02046_),
    .B(_02041_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21oi_2 _09494_ (.A1(_02378_),
    .A2(_02005_),
    .B1(_02379_),
    .Y(_02380_));
 sky130_fd_sc_hd__inv_2 _09495_ (.A(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__nand2_1 _09496_ (.A(_02377_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__nand3_1 _09497_ (.A(_02380_),
    .B(_02374_),
    .C(_02376_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _09498_ (.A(_02382_),
    .B(_02383_),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _09499_ (.A(_02092_),
    .B(_02064_),
    .Y(_02385_));
 sky130_fd_sc_hd__nor2_1 _09500_ (.A(_02064_),
    .B(_02092_),
    .Y(_02387_));
 sky130_fd_sc_hd__a21oi_1 _09501_ (.A1(_02107_),
    .A2(_02385_),
    .B1(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__inv_2 _09502_ (.A(_02388_),
    .Y(_02389_));
 sky130_fd_sc_hd__nand2_1 _09503_ (.A(_02384_),
    .B(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__nand3_1 _09504_ (.A(_02382_),
    .B(_02383_),
    .C(_02388_),
    .Y(_02391_));
 sky130_fd_sc_hd__nand2_1 _09505_ (.A(_02390_),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__inv_2 _09506_ (.A(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__nand2_1 _09507_ (.A(_02319_),
    .B(_02393_),
    .Y(_02394_));
 sky130_fd_sc_hd__nand3_1 _09508_ (.A(_02315_),
    .B(_02318_),
    .C(_02392_),
    .Y(_02395_));
 sky130_fd_sc_hd__nand2_1 _09509_ (.A(_02394_),
    .B(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__nand2_1 _09510_ (.A(_01917_),
    .B(_02061_),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _09511_ (.A(_02061_),
    .B(_01917_),
    .Y(_02399_));
 sky130_fd_sc_hd__a21oi_2 _09512_ (.A1(_02398_),
    .A2(_02129_),
    .B1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__nand2b_1 _09513_ (.A_N(_02396_),
    .B(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__nand2b_1 _09514_ (.A_N(_02400_),
    .B(_02396_),
    .Y(_02402_));
 sky130_fd_sc_hd__nand3b_1 _09515_ (.A_N(_02174_),
    .B(_02401_),
    .C(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _09516_ (.A(_02400_),
    .B(_02396_),
    .Y(_02404_));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(_02396_),
    .B(_02400_),
    .Y(_02405_));
 sky130_fd_sc_hd__nand3b_1 _09518_ (.A_N(_02404_),
    .B(_02174_),
    .C(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__nand3_2 _09519_ (.A(_02169_),
    .B(_02403_),
    .C(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _09520_ (.A(_02406_),
    .B(_02403_),
    .Y(_02409_));
 sky130_fd_sc_hd__a21oi_1 _09521_ (.A1(_02166_),
    .A2(_02138_),
    .B1(_02168_),
    .Y(_02410_));
 sky130_fd_sc_hd__nand2_1 _09522_ (.A(_02409_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__nand2_1 _09523_ (.A(_02407_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _09524_ (.A(_02412_),
    .B(_02149_),
    .Y(_02413_));
 sky130_fd_sc_hd__inv_2 _09525_ (.A(_02149_),
    .Y(_02414_));
 sky130_fd_sc_hd__nand3_1 _09526_ (.A(_02414_),
    .B(_02407_),
    .C(_02411_),
    .Y(_02415_));
 sky130_fd_sc_hd__nand2_1 _09527_ (.A(_02413_),
    .B(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__nand2_1 _09528_ (.A(_02164_),
    .B(_02152_),
    .Y(_02417_));
 sky130_fd_sc_hd__xnor2_1 _09529_ (.A(_02416_),
    .B(_02417_),
    .Y(\m1.out[21] ));
 sky130_fd_sc_hd__nor2_1 _09530_ (.A(_02260_),
    .B(_02255_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21oi_1 _09531_ (.A1(_02312_),
    .A2(_02313_),
    .B1(_02419_),
    .Y(_02420_));
 sky130_fd_sc_hd__nor2_1 _09532_ (.A(_02199_),
    .B(_02195_),
    .Y(_02421_));
 sky130_fd_sc_hd__a21oi_1 _09533_ (.A1(_02218_),
    .A2(_02219_),
    .B1(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__buf_4 _09534_ (.A(net47),
    .X(_02423_));
 sky130_fd_sc_hd__nand2_1 _09535_ (.A(_06270_),
    .B(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__inv_2 _09536_ (.A(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__nand2_1 _09537_ (.A(_06269_),
    .B(_02181_),
    .Y(_02426_));
 sky130_fd_sc_hd__nand2_1 _09538_ (.A(_02425_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__inv_2 _09539_ (.A(_02426_),
    .Y(_02428_));
 sky130_fd_sc_hd__nand2_1 _09540_ (.A(_02428_),
    .B(_02424_),
    .Y(_02430_));
 sky130_fd_sc_hd__nand2_1 _09541_ (.A(_06392_),
    .B(_01921_),
    .Y(_02431_));
 sky130_fd_sc_hd__nand3_2 _09542_ (.A(_02427_),
    .B(_02430_),
    .C(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(_02428_),
    .B(_02425_),
    .Y(_02433_));
 sky130_fd_sc_hd__inv_2 _09544_ (.A(_02431_),
    .Y(_02434_));
 sky130_fd_sc_hd__nand2_1 _09545_ (.A(_02426_),
    .B(_02424_),
    .Y(_02435_));
 sky130_fd_sc_hd__nand3_2 _09546_ (.A(_02433_),
    .B(_02434_),
    .C(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__nand2_1 _09547_ (.A(_02432_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__nor2_1 _09548_ (.A(_02184_),
    .B(_02182_),
    .Y(_02438_));
 sky130_fd_sc_hd__a21oi_2 _09549_ (.A1(_02193_),
    .A2(_02192_),
    .B1(_02438_),
    .Y(_02439_));
 sky130_fd_sc_hd__inv_2 _09550_ (.A(_02439_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_1 _09551_ (.A(_02437_),
    .B(_02441_),
    .Y(_02442_));
 sky130_fd_sc_hd__nand3_1 _09552_ (.A(_02439_),
    .B(_02432_),
    .C(_02436_),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _09553_ (.A(_06262_),
    .B(_06178_),
    .Y(_02444_));
 sky130_fd_sc_hd__inv_2 _09554_ (.A(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__nand2_1 _09555_ (.A(_06273_),
    .B(_01692_),
    .Y(_02446_));
 sky130_fd_sc_hd__inv_2 _09556_ (.A(_02446_),
    .Y(_02447_));
 sky130_fd_sc_hd__nand2_1 _09557_ (.A(_02445_),
    .B(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__nand2_1 _09558_ (.A(_02444_),
    .B(_02446_),
    .Y(_02449_));
 sky130_fd_sc_hd__nand2_1 _09559_ (.A(_02448_),
    .B(_02449_),
    .Y(_02450_));
 sky130_fd_sc_hd__nand2_1 _09560_ (.A(_06259_),
    .B(_06171_),
    .Y(_02451_));
 sky130_fd_sc_hd__nand2_1 _09561_ (.A(_02450_),
    .B(_02451_),
    .Y(_02452_));
 sky130_fd_sc_hd__inv_2 _09562_ (.A(_02451_),
    .Y(_02453_));
 sky130_fd_sc_hd__nand3_1 _09563_ (.A(_02448_),
    .B(_02453_),
    .C(_02449_),
    .Y(_02454_));
 sky130_fd_sc_hd__nand2_2 _09564_ (.A(_02452_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__nand3_1 _09565_ (.A(_02442_),
    .B(_02443_),
    .C(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__nand2_1 _09566_ (.A(_02442_),
    .B(_02443_),
    .Y(_02457_));
 sky130_fd_sc_hd__inv_2 _09567_ (.A(_02455_),
    .Y(_02458_));
 sky130_fd_sc_hd__nand2_1 _09568_ (.A(_02457_),
    .B(_02458_),
    .Y(_02459_));
 sky130_fd_sc_hd__nand3_1 _09569_ (.A(_02422_),
    .B(_02456_),
    .C(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__nand2_1 _09570_ (.A(_02459_),
    .B(_02456_),
    .Y(_02462_));
 sky130_fd_sc_hd__nand2_1 _09571_ (.A(_02220_),
    .B(_02217_),
    .Y(_02463_));
 sky130_fd_sc_hd__nand2_1 _09572_ (.A(_02462_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__nand2_1 _09573_ (.A(_02460_),
    .B(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__nand2_1 _09574_ (.A(_00299_),
    .B(net39),
    .Y(_02466_));
 sky130_fd_sc_hd__inv_2 _09575_ (.A(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__nand2_1 _09576_ (.A(_06265_),
    .B(_06173_),
    .Y(_02468_));
 sky130_fd_sc_hd__nand2_1 _09577_ (.A(_02467_),
    .B(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__inv_2 _09578_ (.A(_02468_),
    .Y(_02470_));
 sky130_fd_sc_hd__nand2_1 _09579_ (.A(_02470_),
    .B(_02466_),
    .Y(_02471_));
 sky130_fd_sc_hd__nand2_1 _09580_ (.A(_00193_),
    .B(_00921_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand3_1 _09581_ (.A(_02469_),
    .B(_02471_),
    .C(_02473_),
    .Y(_02474_));
 sky130_fd_sc_hd__nand2_1 _09582_ (.A(_02467_),
    .B(_02470_),
    .Y(_02475_));
 sky130_fd_sc_hd__inv_2 _09583_ (.A(_02473_),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_1 _09584_ (.A(_02466_),
    .B(_02468_),
    .Y(_02477_));
 sky130_fd_sc_hd__nand3_1 _09585_ (.A(_02475_),
    .B(_02476_),
    .C(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_02474_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _09587_ (.A(_02204_),
    .B(_02202_),
    .Y(_02480_));
 sky130_fd_sc_hd__a21oi_2 _09588_ (.A1(_02213_),
    .A2(_02212_),
    .B1(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hd__inv_2 _09589_ (.A(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__nand2_1 _09590_ (.A(_02479_),
    .B(_02482_),
    .Y(_02484_));
 sky130_fd_sc_hd__nand3_1 _09591_ (.A(_02481_),
    .B(_02474_),
    .C(_02478_),
    .Y(_02485_));
 sky130_fd_sc_hd__nand2_1 _09592_ (.A(_02484_),
    .B(_02485_),
    .Y(_02486_));
 sky130_fd_sc_hd__nand2_1 _09593_ (.A(_02238_),
    .B(_02235_),
    .Y(_02487_));
 sky130_fd_sc_hd__nand2_1 _09594_ (.A(_02486_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__nand3b_1 _09595_ (.A_N(_02487_),
    .B(_02484_),
    .C(_02485_),
    .Y(_02489_));
 sky130_fd_sc_hd__nand2_2 _09596_ (.A(_02488_),
    .B(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__inv_2 _09597_ (.A(_02490_),
    .Y(_02491_));
 sky130_fd_sc_hd__nand2_1 _09598_ (.A(_02465_),
    .B(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__nand3_1 _09599_ (.A(_02460_),
    .B(_02464_),
    .C(_02490_),
    .Y(_02493_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_02492_),
    .B(_02493_),
    .Y(_02495_));
 sky130_fd_sc_hd__nand2_1 _09601_ (.A(_02223_),
    .B(_02179_),
    .Y(_02496_));
 sky130_fd_sc_hd__nor2_1 _09602_ (.A(_02179_),
    .B(_02223_),
    .Y(_02497_));
 sky130_fd_sc_hd__a21oi_2 _09603_ (.A1(_02496_),
    .A2(_02251_),
    .B1(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__inv_2 _09604_ (.A(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__nand2_1 _09605_ (.A(_02495_),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__nand3_1 _09606_ (.A(_02498_),
    .B(_02492_),
    .C(_02493_),
    .Y(_02501_));
 sky130_fd_sc_hd__nand2_1 _09607_ (.A(_02239_),
    .B(_02241_),
    .Y(_02502_));
 sky130_fd_sc_hd__nor2_1 _09608_ (.A(_02241_),
    .B(_02239_),
    .Y(_02503_));
 sky130_fd_sc_hd__a21oi_2 _09609_ (.A1(_02502_),
    .A2(_02247_),
    .B1(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__inv_2 _09610_ (.A(_02504_),
    .Y(_02506_));
 sky130_fd_sc_hd__nor2_1 _09611_ (.A(_02264_),
    .B(_02267_),
    .Y(_02507_));
 sky130_fd_sc_hd__a21oi_2 _09612_ (.A1(_02275_),
    .A2(_02274_),
    .B1(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__inv_2 _09613_ (.A(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__nand2_1 _09614_ (.A(_06292_),
    .B(_06221_),
    .Y(_02510_));
 sky130_fd_sc_hd__inv_2 _09615_ (.A(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2_1 _09616_ (.A(_06288_),
    .B(_06218_),
    .Y(_02512_));
 sky130_fd_sc_hd__nand2_1 _09617_ (.A(_02511_),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__inv_2 _09618_ (.A(_02512_),
    .Y(_02514_));
 sky130_fd_sc_hd__nand2_1 _09619_ (.A(_02514_),
    .B(_02510_),
    .Y(_02515_));
 sky130_fd_sc_hd__nand2_1 _09620_ (.A(_06291_),
    .B(_06228_),
    .Y(_02517_));
 sky130_fd_sc_hd__nand3_1 _09621_ (.A(_02513_),
    .B(_02515_),
    .C(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__nand2_1 _09622_ (.A(_02511_),
    .B(_02514_),
    .Y(_02519_));
 sky130_fd_sc_hd__inv_2 _09623_ (.A(_02517_),
    .Y(_02520_));
 sky130_fd_sc_hd__nand2_1 _09624_ (.A(_02510_),
    .B(_02512_),
    .Y(_02521_));
 sky130_fd_sc_hd__nand3_1 _09625_ (.A(_02519_),
    .B(_02520_),
    .C(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__nand3_1 _09626_ (.A(_02509_),
    .B(_02518_),
    .C(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _09627_ (.A(_02518_),
    .B(_02522_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand2_1 _09628_ (.A(_02524_),
    .B(_02508_),
    .Y(_02525_));
 sky130_fd_sc_hd__nand2_1 _09629_ (.A(_00701_),
    .B(_06225_),
    .Y(_02526_));
 sky130_fd_sc_hd__inv_2 _09630_ (.A(_02526_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand2_1 _09631_ (.A(_06280_),
    .B(_06231_),
    .Y(_02529_));
 sky130_fd_sc_hd__inv_2 _09632_ (.A(_02529_),
    .Y(_02530_));
 sky130_fd_sc_hd__nand2_1 _09633_ (.A(_02528_),
    .B(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _09634_ (.A(_02526_),
    .B(_02529_),
    .Y(_02532_));
 sky130_fd_sc_hd__nand2_1 _09635_ (.A(_02531_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__nand2_1 _09636_ (.A(_06284_),
    .B(_06226_),
    .Y(_02534_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_02533_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__inv_2 _09638_ (.A(_02534_),
    .Y(_02536_));
 sky130_fd_sc_hd__nand3_1 _09639_ (.A(_02531_),
    .B(_02536_),
    .C(_02532_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2_1 _09640_ (.A(_02535_),
    .B(_02537_),
    .Y(_02539_));
 sky130_fd_sc_hd__inv_2 _09641_ (.A(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand3_2 _09642_ (.A(_02523_),
    .B(_02525_),
    .C(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__nand2_1 _09643_ (.A(_02524_),
    .B(_02509_),
    .Y(_02542_));
 sky130_fd_sc_hd__nand3_1 _09644_ (.A(_02508_),
    .B(_02518_),
    .C(_02522_),
    .Y(_02543_));
 sky130_fd_sc_hd__nand3_1 _09645_ (.A(_02542_),
    .B(_02543_),
    .C(_02539_),
    .Y(_02544_));
 sky130_fd_sc_hd__nand2_1 _09646_ (.A(_02541_),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__nand2_1 _09647_ (.A(_02506_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand3_1 _09648_ (.A(_02504_),
    .B(_02544_),
    .C(_02541_),
    .Y(_02547_));
 sky130_fd_sc_hd__nand2_1 _09649_ (.A(_02546_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__or2_1 _09650_ (.A(_02280_),
    .B(_02278_),
    .X(_02550_));
 sky130_fd_sc_hd__nand2_1 _09651_ (.A(_02299_),
    .B(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__nand2_1 _09652_ (.A(_02548_),
    .B(_02551_),
    .Y(_02552_));
 sky130_fd_sc_hd__nand3b_1 _09653_ (.A_N(_02551_),
    .B(_02546_),
    .C(_02547_),
    .Y(_02553_));
 sky130_fd_sc_hd__nand2_1 _09654_ (.A(_02552_),
    .B(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__nand3_1 _09655_ (.A(_02500_),
    .B(_02501_),
    .C(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__nand2_1 _09656_ (.A(_02500_),
    .B(_02501_),
    .Y(_02556_));
 sky130_fd_sc_hd__inv_2 _09657_ (.A(_02554_),
    .Y(_02557_));
 sky130_fd_sc_hd__nand2_1 _09658_ (.A(_02556_),
    .B(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand3_1 _09659_ (.A(_02420_),
    .B(_02555_),
    .C(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_1 _09660_ (.A(_02558_),
    .B(_02555_),
    .Y(_02561_));
 sky130_fd_sc_hd__nand2_1 _09661_ (.A(_02314_),
    .B(_02311_),
    .Y(_02562_));
 sky130_fd_sc_hd__nand2_1 _09662_ (.A(_02561_),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand2_1 _09663_ (.A(_02559_),
    .B(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__nand2_1 _09664_ (.A(_02302_),
    .B(_02263_),
    .Y(_02565_));
 sky130_fd_sc_hd__nor2_1 _09665_ (.A(_02263_),
    .B(_02302_),
    .Y(_02566_));
 sky130_fd_sc_hd__a21oi_2 _09666_ (.A1(_02565_),
    .A2(_02305_),
    .B1(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__inv_2 _09667_ (.A(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__nor2_1 _09668_ (.A(_02333_),
    .B(_02332_),
    .Y(_02569_));
 sky130_fd_sc_hd__a21oi_1 _09669_ (.A1(_02334_),
    .A2(_02337_),
    .B1(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _09670_ (.A(_01211_),
    .B(_06202_),
    .Y(_02572_));
 sky130_fd_sc_hd__inv_2 _09671_ (.A(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__nand2_1 _09672_ (.A(_01831_),
    .B(_06200_),
    .Y(_02574_));
 sky130_fd_sc_hd__inv_2 _09673_ (.A(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__nand2_1 _09674_ (.A(_02573_),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__nand2_1 _09675_ (.A(_02572_),
    .B(_02574_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_1 _09676_ (.A(_02576_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__nand2_1 _09677_ (.A(_06236_),
    .B(_06196_),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _09678_ (.A(_02578_),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__nand3b_2 _09679_ (.A_N(_02579_),
    .B(_02576_),
    .C(_02577_),
    .Y(_02581_));
 sky130_fd_sc_hd__nand2_1 _09680_ (.A(_02580_),
    .B(_02581_),
    .Y(_02583_));
 sky130_fd_sc_hd__a21o_1 _09681_ (.A1(_02288_),
    .A2(_02292_),
    .B1(_02286_),
    .X(_02584_));
 sky130_fd_sc_hd__nand2_1 _09682_ (.A(_02583_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__a21oi_2 _09683_ (.A1(_02288_),
    .A2(_02292_),
    .B1(_02286_),
    .Y(_02586_));
 sky130_fd_sc_hd__nand3_1 _09684_ (.A(_02580_),
    .B(_02581_),
    .C(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand2_2 _09685_ (.A(_02330_),
    .B(_02325_),
    .Y(_02588_));
 sky130_fd_sc_hd__inv_2 _09686_ (.A(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__nand3_1 _09687_ (.A(_02585_),
    .B(_02587_),
    .C(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__nand2_1 _09688_ (.A(_02583_),
    .B(_02586_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand3_1 _09689_ (.A(_02584_),
    .B(_02581_),
    .C(_02580_),
    .Y(_02592_));
 sky130_fd_sc_hd__nand3_2 _09690_ (.A(_02591_),
    .B(_02592_),
    .C(_02588_),
    .Y(_02594_));
 sky130_fd_sc_hd__nand3_1 _09691_ (.A(_02570_),
    .B(_02590_),
    .C(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_1 _09692_ (.A(_01858_),
    .B(_06211_),
    .Y(_02596_));
 sky130_fd_sc_hd__nand2_1 _09693_ (.A(_06242_),
    .B(_06198_),
    .Y(_02597_));
 sky130_fd_sc_hd__nor2_1 _09694_ (.A(_02596_),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__inv_2 _09695_ (.A(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__nand2_1 _09696_ (.A(_02596_),
    .B(_02597_),
    .Y(_02600_));
 sky130_fd_sc_hd__nand2_1 _09697_ (.A(_02599_),
    .B(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand2_1 _09698_ (.A(_02095_),
    .B(_06214_),
    .Y(_02602_));
 sky130_fd_sc_hd__nand2_1 _09699_ (.A(_02601_),
    .B(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hd__inv_2 _09700_ (.A(_02602_),
    .Y(_02605_));
 sky130_fd_sc_hd__nand3_1 _09701_ (.A(_02599_),
    .B(_02600_),
    .C(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__nand2_1 _09702_ (.A(_02603_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand3_1 _09703_ (.A(_02607_),
    .B(_02356_),
    .C(_02363_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_1 _09704_ (.A(_02363_),
    .B(_02356_),
    .Y(_02609_));
 sky130_fd_sc_hd__nand3_1 _09705_ (.A(_02609_),
    .B(_02603_),
    .C(_02606_),
    .Y(_02610_));
 sky130_fd_sc_hd__nand2_1 _09706_ (.A(_02608_),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__and4_1 _09707_ (.A(_06246_),
    .B(_06298_),
    .C(_06205_),
    .D(_06207_),
    .X(_02612_));
 sky130_fd_sc_hd__inv_2 _09708_ (.A(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hd__a22o_1 _09709_ (.A1(_06247_),
    .A2(_06206_),
    .B1(_06299_),
    .B2(_06208_),
    .X(_02614_));
 sky130_fd_sc_hd__nand2_1 _09710_ (.A(_02613_),
    .B(_02614_),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _09711_ (.A(_02611_),
    .B(_02616_),
    .Y(_02617_));
 sky130_fd_sc_hd__nand3b_1 _09712_ (.A_N(_02616_),
    .B(_02608_),
    .C(_02610_),
    .Y(_02618_));
 sky130_fd_sc_hd__nand2_1 _09713_ (.A(_02617_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__nand2_1 _09714_ (.A(_02338_),
    .B(_02336_),
    .Y(_02620_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(_02594_),
    .B(_02590_),
    .Y(_02621_));
 sky130_fd_sc_hd__nand2_1 _09716_ (.A(_02620_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__nand3_1 _09717_ (.A(_02595_),
    .B(_02619_),
    .C(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_1 _09718_ (.A(_02595_),
    .B(_02622_),
    .Y(_02624_));
 sky130_fd_sc_hd__inv_2 _09719_ (.A(_02619_),
    .Y(_02625_));
 sky130_fd_sc_hd__nand2_1 _09720_ (.A(_02624_),
    .B(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand3_1 _09721_ (.A(_02568_),
    .B(_02623_),
    .C(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__nand2_1 _09722_ (.A(_02626_),
    .B(_02623_),
    .Y(_02628_));
 sky130_fd_sc_hd__nand2_1 _09723_ (.A(_02628_),
    .B(_02567_),
    .Y(_02629_));
 sky130_fd_sc_hd__nand2_1 _09724_ (.A(_02627_),
    .B(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand3_1 _09725_ (.A(_02347_),
    .B(_02343_),
    .C(_02338_),
    .Y(_02631_));
 sky130_fd_sc_hd__nand2_1 _09726_ (.A(_02374_),
    .B(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__inv_2 _09727_ (.A(_02632_),
    .Y(_02633_));
 sky130_fd_sc_hd__nand2_1 _09728_ (.A(_02630_),
    .B(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__nand3_1 _09729_ (.A(_02627_),
    .B(_02629_),
    .C(_02632_),
    .Y(_02635_));
 sky130_fd_sc_hd__nand2_1 _09730_ (.A(_02634_),
    .B(_02635_),
    .Y(_02637_));
 sky130_fd_sc_hd__inv_2 _09731_ (.A(_02637_),
    .Y(_02638_));
 sky130_fd_sc_hd__nand2_1 _09732_ (.A(_02564_),
    .B(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hd__nand3_1 _09733_ (.A(_02559_),
    .B(_02563_),
    .C(_02637_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _09734_ (.A(_02639_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__nand2_1 _09735_ (.A(_02316_),
    .B(_02176_),
    .Y(_02642_));
 sky130_fd_sc_hd__nor2_1 _09736_ (.A(_02176_),
    .B(_02316_),
    .Y(_02643_));
 sky130_fd_sc_hd__a21oi_2 _09737_ (.A1(_02642_),
    .A2(_02393_),
    .B1(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__inv_2 _09738_ (.A(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand2_1 _09739_ (.A(_02641_),
    .B(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand3_1 _09740_ (.A(_02644_),
    .B(_02639_),
    .C(_02640_),
    .Y(_02648_));
 sky130_fd_sc_hd__nand2_1 _09741_ (.A(_02646_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__and2_1 _09742_ (.A(_02371_),
    .B(_02365_),
    .X(_02650_));
 sky130_fd_sc_hd__o21a_1 _09743_ (.A1(_02377_),
    .A2(_02380_),
    .B1(_02390_),
    .X(_02651_));
 sky130_fd_sc_hd__nor2_1 _09744_ (.A(_02650_),
    .B(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hd__inv_2 _09745_ (.A(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__nand2_1 _09746_ (.A(_02651_),
    .B(_02650_),
    .Y(_02654_));
 sky130_fd_sc_hd__nand2_1 _09747_ (.A(_02653_),
    .B(_02654_),
    .Y(_02655_));
 sky130_fd_sc_hd__inv_2 _09748_ (.A(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2_1 _09749_ (.A(_02649_),
    .B(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hd__nand3_1 _09750_ (.A(_02646_),
    .B(_02648_),
    .C(_02655_),
    .Y(_02659_));
 sky130_fd_sc_hd__nand2_1 _09751_ (.A(_02657_),
    .B(_02659_),
    .Y(_02660_));
 sky130_fd_sc_hd__a21o_1 _09752_ (.A1(_02405_),
    .A2(_02174_),
    .B1(_02404_),
    .X(_02661_));
 sky130_fd_sc_hd__nand2_1 _09753_ (.A(_02660_),
    .B(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__a21oi_1 _09754_ (.A1(_02405_),
    .A2(_02174_),
    .B1(_02404_),
    .Y(_02663_));
 sky130_fd_sc_hd__nand3_1 _09755_ (.A(_02663_),
    .B(_02657_),
    .C(_02659_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand2_1 _09756_ (.A(_02662_),
    .B(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _09757_ (.A(_02665_),
    .B(_02172_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand3b_1 _09758_ (.A_N(_02172_),
    .B(_02662_),
    .C(_02664_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand2_1 _09759_ (.A(_02666_),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__nand2_1 _09760_ (.A(_02668_),
    .B(_02407_),
    .Y(_02670_));
 sky130_fd_sc_hd__inv_2 _09761_ (.A(_02407_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand3_1 _09762_ (.A(_02666_),
    .B(_02667_),
    .C(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand2_1 _09763_ (.A(_02670_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__inv_2 _09764_ (.A(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__nor2_1 _09765_ (.A(_02416_),
    .B(_02154_),
    .Y(_02675_));
 sky130_fd_sc_hd__nand3_1 _09766_ (.A(_02151_),
    .B(_02413_),
    .C(_02415_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _09767_ (.A(_02676_),
    .B(_02415_),
    .Y(_02677_));
 sky130_fd_sc_hd__a21o_1 _09768_ (.A1(_02162_),
    .A2(_02675_),
    .B1(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__or2_1 _09769_ (.A(_02674_),
    .B(_02678_),
    .X(_02679_));
 sky130_fd_sc_hd__nand2_1 _09770_ (.A(_02678_),
    .B(_02674_),
    .Y(_02681_));
 sky130_fd_sc_hd__and2_1 _09771_ (.A(_02679_),
    .B(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__clkbuf_1 _09772_ (.A(_02682_),
    .X(\m1.out[22] ));
 sky130_fd_sc_hd__nand2_1 _09773_ (.A(_02561_),
    .B(_02420_),
    .Y(_02683_));
 sky130_fd_sc_hd__nor2_1 _09774_ (.A(_02420_),
    .B(_02561_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21oi_1 _09775_ (.A1(_02638_),
    .A2(_02683_),
    .B1(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__nand2_1 _09776_ (.A(_02495_),
    .B(_02498_),
    .Y(_02686_));
 sky130_fd_sc_hd__nor2_1 _09777_ (.A(_02498_),
    .B(_02495_),
    .Y(_02687_));
 sky130_fd_sc_hd__a21oi_1 _09778_ (.A1(_02686_),
    .A2(_02557_),
    .B1(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__nand2_1 _09779_ (.A(_02462_),
    .B(_02422_),
    .Y(_02689_));
 sky130_fd_sc_hd__nor2_1 _09780_ (.A(_02422_),
    .B(_02462_),
    .Y(_02691_));
 sky130_fd_sc_hd__a21oi_1 _09781_ (.A1(_02689_),
    .A2(_02491_),
    .B1(_02691_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _09782_ (.A(_02437_),
    .B(_02439_),
    .Y(_02693_));
 sky130_fd_sc_hd__nor2_1 _09783_ (.A(_02439_),
    .B(_02437_),
    .Y(_02694_));
 sky130_fd_sc_hd__a21oi_1 _09784_ (.A1(_02693_),
    .A2(_02458_),
    .B1(_02694_),
    .Y(_02695_));
 sky130_fd_sc_hd__nor2_1 _09785_ (.A(_02426_),
    .B(_02424_),
    .Y(_02696_));
 sky130_fd_sc_hd__a21oi_2 _09786_ (.A1(_02435_),
    .A2(_02434_),
    .B1(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__nand2_1 _09787_ (.A(_06327_),
    .B(_02423_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_1 _09788_ (.A(_02698_),
    .B(_06329_),
    .Y(_02699_));
 sky130_fd_sc_hd__nand3_1 _09789_ (.A(_06269_),
    .B(_06271_),
    .C(_02423_),
    .Y(_02700_));
 sky130_fd_sc_hd__nand2_1 _09790_ (.A(_02699_),
    .B(_02700_),
    .Y(_02702_));
 sky130_fd_sc_hd__nand2_1 _09791_ (.A(_06392_),
    .B(_02180_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand2_1 _09792_ (.A(_02702_),
    .B(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__inv_2 _09793_ (.A(_02703_),
    .Y(_02705_));
 sky130_fd_sc_hd__nand3_1 _09794_ (.A(_02699_),
    .B(_02700_),
    .C(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hd__nand3_1 _09795_ (.A(_02697_),
    .B(_02704_),
    .C(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__inv_2 _09796_ (.A(_02697_),
    .Y(_02708_));
 sky130_fd_sc_hd__nand2_1 _09797_ (.A(_02704_),
    .B(_02706_),
    .Y(_02709_));
 sky130_fd_sc_hd__nand2_1 _09798_ (.A(_02708_),
    .B(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(_06273_),
    .B(_01921_),
    .Y(_02711_));
 sky130_fd_sc_hd__inv_2 _09800_ (.A(_02711_),
    .Y(_02713_));
 sky130_fd_sc_hd__nand2_1 _09801_ (.A(_06261_),
    .B(_01692_),
    .Y(_02714_));
 sky130_fd_sc_hd__nand2_1 _09802_ (.A(_02713_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__inv_2 _09803_ (.A(_02714_),
    .Y(_02716_));
 sky130_fd_sc_hd__nand2_1 _09804_ (.A(_02716_),
    .B(_02711_),
    .Y(_02717_));
 sky130_fd_sc_hd__nand2_1 _09805_ (.A(_00175_),
    .B(_06177_),
    .Y(_02718_));
 sky130_fd_sc_hd__nand3_1 _09806_ (.A(_02715_),
    .B(_02717_),
    .C(_02718_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand2_1 _09807_ (.A(_02716_),
    .B(_02713_),
    .Y(_02720_));
 sky130_fd_sc_hd__inv_2 _09808_ (.A(_02718_),
    .Y(_02721_));
 sky130_fd_sc_hd__nand2_1 _09809_ (.A(_02714_),
    .B(_02711_),
    .Y(_02722_));
 sky130_fd_sc_hd__nand3_1 _09810_ (.A(_02720_),
    .B(_02721_),
    .C(_02722_),
    .Y(_02724_));
 sky130_fd_sc_hd__nand2_1 _09811_ (.A(_02719_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand3_2 _09812_ (.A(_02707_),
    .B(_02710_),
    .C(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__inv_2 _09813_ (.A(_02709_),
    .Y(_02727_));
 sky130_fd_sc_hd__nand2_1 _09814_ (.A(_02727_),
    .B(_02708_),
    .Y(_02728_));
 sky130_fd_sc_hd__inv_2 _09815_ (.A(_02725_),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_1 _09816_ (.A(_02709_),
    .B(_02697_),
    .Y(_02730_));
 sky130_fd_sc_hd__nand3_2 _09817_ (.A(_02728_),
    .B(_02729_),
    .C(_02730_),
    .Y(_02731_));
 sky130_fd_sc_hd__nand3_1 _09818_ (.A(_02695_),
    .B(_02726_),
    .C(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__a21o_1 _09819_ (.A1(_02693_),
    .A2(_02458_),
    .B1(_02694_),
    .X(_02733_));
 sky130_fd_sc_hd__nand2_1 _09820_ (.A(_02731_),
    .B(_02726_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand2_1 _09821_ (.A(_02733_),
    .B(_02735_),
    .Y(_02736_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(_02444_),
    .B(_02446_),
    .Y(_02737_));
 sky130_fd_sc_hd__a21o_1 _09823_ (.A1(_02449_),
    .A2(_02453_),
    .B1(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__nand2_1 _09824_ (.A(_06264_),
    .B(_01278_),
    .Y(_02739_));
 sky130_fd_sc_hd__inv_2 _09825_ (.A(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__nand2_1 _09826_ (.A(_06266_),
    .B(_01280_),
    .Y(_02741_));
 sky130_fd_sc_hd__nand2_1 _09827_ (.A(_02740_),
    .B(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__inv_2 _09828_ (.A(_02741_),
    .Y(_02743_));
 sky130_fd_sc_hd__nand2_1 _09829_ (.A(_02743_),
    .B(_02739_),
    .Y(_02744_));
 sky130_fd_sc_hd__nand2_1 _09830_ (.A(_06290_),
    .B(_00918_),
    .Y(_02746_));
 sky130_fd_sc_hd__nand3_1 _09831_ (.A(_02742_),
    .B(_02744_),
    .C(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__nand2_1 _09832_ (.A(_02740_),
    .B(_02743_),
    .Y(_02748_));
 sky130_fd_sc_hd__inv_2 _09833_ (.A(_02746_),
    .Y(_02749_));
 sky130_fd_sc_hd__nand2_1 _09834_ (.A(_02739_),
    .B(_02741_),
    .Y(_02750_));
 sky130_fd_sc_hd__nand3_1 _09835_ (.A(_02748_),
    .B(_02749_),
    .C(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__nand3_1 _09836_ (.A(_02738_),
    .B(_02747_),
    .C(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__nand2_1 _09837_ (.A(_02747_),
    .B(_02751_),
    .Y(_02753_));
 sky130_fd_sc_hd__a21oi_1 _09838_ (.A1(_02449_),
    .A2(_02453_),
    .B1(_02737_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _09839_ (.A(_02753_),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(_02478_),
    .B(_02475_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand3_1 _09841_ (.A(_02752_),
    .B(_02755_),
    .C(_02757_),
    .Y(_02758_));
 sky130_fd_sc_hd__nand2_1 _09842_ (.A(_02753_),
    .B(_02738_),
    .Y(_02759_));
 sky130_fd_sc_hd__nand3_1 _09843_ (.A(_02754_),
    .B(_02747_),
    .C(_02751_),
    .Y(_02760_));
 sky130_fd_sc_hd__inv_2 _09844_ (.A(_02757_),
    .Y(_02761_));
 sky130_fd_sc_hd__nand3_1 _09845_ (.A(_02759_),
    .B(_02760_),
    .C(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__nand2_2 _09846_ (.A(_02758_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand3_1 _09847_ (.A(_02732_),
    .B(_02736_),
    .C(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__inv_2 _09848_ (.A(_02735_),
    .Y(_02765_));
 sky130_fd_sc_hd__nand2_1 _09849_ (.A(_02765_),
    .B(_02733_),
    .Y(_02766_));
 sky130_fd_sc_hd__inv_2 _09850_ (.A(_02763_),
    .Y(_02768_));
 sky130_fd_sc_hd__nand2_1 _09851_ (.A(_02735_),
    .B(_02695_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand3_1 _09852_ (.A(_02766_),
    .B(_02768_),
    .C(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand3_1 _09853_ (.A(_02692_),
    .B(_02764_),
    .C(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__nand2_1 _09854_ (.A(_02770_),
    .B(_02764_),
    .Y(_02772_));
 sky130_fd_sc_hd__a21o_1 _09855_ (.A1(_02689_),
    .A2(_02491_),
    .B1(_02691_),
    .X(_02773_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(_02772_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2_1 _09857_ (.A(_02479_),
    .B(_02481_),
    .Y(_02775_));
 sky130_fd_sc_hd__nor2_1 _09858_ (.A(_02481_),
    .B(_02479_),
    .Y(_02776_));
 sky130_fd_sc_hd__a21oi_1 _09859_ (.A1(_02775_),
    .A2(_02487_),
    .B1(_02776_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(_06292_),
    .B(_00926_),
    .Y(_02779_));
 sky130_fd_sc_hd__inv_2 _09861_ (.A(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__nand2_2 _09862_ (.A(_06287_),
    .B(_00921_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand2_1 _09863_ (.A(_02780_),
    .B(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__inv_2 _09864_ (.A(_02781_),
    .Y(_02783_));
 sky130_fd_sc_hd__nand2_1 _09865_ (.A(_02783_),
    .B(_02779_),
    .Y(_02784_));
 sky130_fd_sc_hd__nand2_1 _09866_ (.A(_00561_),
    .B(_06220_),
    .Y(_02785_));
 sky130_fd_sc_hd__nand3_1 _09867_ (.A(_02782_),
    .B(_02784_),
    .C(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__nand2_1 _09868_ (.A(_02780_),
    .B(_02783_),
    .Y(_02787_));
 sky130_fd_sc_hd__inv_2 _09869_ (.A(_02785_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _09870_ (.A(_02779_),
    .B(_02781_),
    .Y(_02790_));
 sky130_fd_sc_hd__nand3_1 _09871_ (.A(_02787_),
    .B(_02788_),
    .C(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__nand2_1 _09872_ (.A(_02786_),
    .B(_02791_),
    .Y(_02792_));
 sky130_fd_sc_hd__nor2_1 _09873_ (.A(_02510_),
    .B(_02512_),
    .Y(_02793_));
 sky130_fd_sc_hd__a21o_1 _09874_ (.A1(_02521_),
    .A2(_02520_),
    .B1(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__nand2_1 _09875_ (.A(_02792_),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__a21oi_1 _09876_ (.A1(_02521_),
    .A2(_02520_),
    .B1(_02793_),
    .Y(_02796_));
 sky130_fd_sc_hd__nand3_1 _09877_ (.A(_02796_),
    .B(_02786_),
    .C(_02791_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_1 _09878_ (.A(_00701_),
    .B(_06230_),
    .Y(_02798_));
 sky130_fd_sc_hd__inv_2 _09879_ (.A(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__nand2_1 _09880_ (.A(_00849_),
    .B(_00376_),
    .Y(_02800_));
 sky130_fd_sc_hd__inv_2 _09881_ (.A(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hd__nand2_1 _09882_ (.A(_02799_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _09883_ (.A(_02798_),
    .B(_02800_),
    .Y(_02803_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(_02802_),
    .B(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__nand2_1 _09885_ (.A(_01158_),
    .B(_00780_),
    .Y(_02805_));
 sky130_fd_sc_hd__nand2_1 _09886_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__inv_2 _09887_ (.A(_02805_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand3_1 _09888_ (.A(_02802_),
    .B(_02807_),
    .C(_02803_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _09889_ (.A(_02806_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand3_1 _09890_ (.A(_02795_),
    .B(_02797_),
    .C(_02809_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand3_1 _09891_ (.A(_02794_),
    .B(_02786_),
    .C(_02791_),
    .Y(_02812_));
 sky130_fd_sc_hd__nand2_1 _09892_ (.A(_02792_),
    .B(_02796_),
    .Y(_02813_));
 sky130_fd_sc_hd__inv_2 _09893_ (.A(_02809_),
    .Y(_02814_));
 sky130_fd_sc_hd__nand3_1 _09894_ (.A(_02812_),
    .B(_02813_),
    .C(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__nand3_1 _09895_ (.A(_02777_),
    .B(_02811_),
    .C(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__a21o_1 _09896_ (.A1(_02775_),
    .A2(_02487_),
    .B1(_02776_),
    .X(_02817_));
 sky130_fd_sc_hd__nand2_1 _09897_ (.A(_02815_),
    .B(_02811_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand2_1 _09898_ (.A(_02817_),
    .B(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__nand2_1 _09899_ (.A(_02816_),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__nand2_1 _09900_ (.A(_02541_),
    .B(_02523_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _09901_ (.A(_02820_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand3b_1 _09902_ (.A_N(_02822_),
    .B(_02816_),
    .C(_02819_),
    .Y(_02824_));
 sky130_fd_sc_hd__nand2_2 _09903_ (.A(_02823_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__nand3_1 _09904_ (.A(_02771_),
    .B(_02774_),
    .C(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__nand2_1 _09905_ (.A(_02771_),
    .B(_02774_),
    .Y(_02827_));
 sky130_fd_sc_hd__inv_2 _09906_ (.A(_02825_),
    .Y(_02828_));
 sky130_fd_sc_hd__nand2_1 _09907_ (.A(_02827_),
    .B(_02828_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand3_1 _09908_ (.A(_02688_),
    .B(_02826_),
    .C(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__nand2_1 _09909_ (.A(_02829_),
    .B(_02826_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21o_1 _09910_ (.A1(_02686_),
    .A2(_02557_),
    .B1(_02687_),
    .X(_02833_));
 sky130_fd_sc_hd__nand2_1 _09911_ (.A(_02831_),
    .B(_02833_),
    .Y(_02834_));
 sky130_fd_sc_hd__nand2_1 _09912_ (.A(_02545_),
    .B(_02504_),
    .Y(_02835_));
 sky130_fd_sc_hd__nor2_1 _09913_ (.A(_02504_),
    .B(_02545_),
    .Y(_02836_));
 sky130_fd_sc_hd__a21o_1 _09914_ (.A1(_02835_),
    .A2(_02551_),
    .B1(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__nor2_1 _09915_ (.A(_02586_),
    .B(_02583_),
    .Y(_02838_));
 sky130_fd_sc_hd__a21oi_1 _09916_ (.A1(_02591_),
    .A2(_02588_),
    .B1(_02838_),
    .Y(_02839_));
 sky130_fd_sc_hd__nand2_1 _09917_ (.A(_01211_),
    .B(_06200_),
    .Y(_02840_));
 sky130_fd_sc_hd__inv_2 _09918_ (.A(_02840_),
    .Y(_02841_));
 sky130_fd_sc_hd__nand2_1 _09919_ (.A(_01831_),
    .B(_06226_),
    .Y(_02842_));
 sky130_fd_sc_hd__inv_2 _09920_ (.A(_02842_),
    .Y(_02844_));
 sky130_fd_sc_hd__nand2_1 _09921_ (.A(_02841_),
    .B(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _09922_ (.A(_02840_),
    .B(_02842_),
    .Y(_02846_));
 sky130_fd_sc_hd__nand2_1 _09923_ (.A(_02845_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__nand2_1 _09924_ (.A(_06236_),
    .B(_06202_),
    .Y(_02848_));
 sky130_fd_sc_hd__nand2_1 _09925_ (.A(_02847_),
    .B(_02848_),
    .Y(_02849_));
 sky130_fd_sc_hd__nand3b_2 _09926_ (.A_N(_02848_),
    .B(_02845_),
    .C(_02846_),
    .Y(_02850_));
 sky130_fd_sc_hd__nand2_1 _09927_ (.A(_02849_),
    .B(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__nor2_1 _09928_ (.A(_02526_),
    .B(_02529_),
    .Y(_02852_));
 sky130_fd_sc_hd__a21o_1 _09929_ (.A1(_02532_),
    .A2(_02536_),
    .B1(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__nand2_1 _09930_ (.A(_02851_),
    .B(_02853_),
    .Y(_02855_));
 sky130_fd_sc_hd__a21oi_1 _09931_ (.A1(_02532_),
    .A2(_02536_),
    .B1(_02852_),
    .Y(_02856_));
 sky130_fd_sc_hd__nand3_1 _09932_ (.A(_02849_),
    .B(_02850_),
    .C(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__nand2_1 _09933_ (.A(_02581_),
    .B(_02576_),
    .Y(_02858_));
 sky130_fd_sc_hd__inv_2 _09934_ (.A(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand3_1 _09935_ (.A(_02855_),
    .B(_02857_),
    .C(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__nand2_1 _09936_ (.A(_02851_),
    .B(_02856_),
    .Y(_02861_));
 sky130_fd_sc_hd__nand3_1 _09937_ (.A(_02853_),
    .B(_02850_),
    .C(_02849_),
    .Y(_02862_));
 sky130_fd_sc_hd__nand3_1 _09938_ (.A(_02861_),
    .B(_02862_),
    .C(_02858_),
    .Y(_02863_));
 sky130_fd_sc_hd__nand3_1 _09939_ (.A(_02839_),
    .B(_02860_),
    .C(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__nand2_1 _09940_ (.A(_02594_),
    .B(_02592_),
    .Y(_02866_));
 sky130_fd_sc_hd__nand2_1 _09941_ (.A(_02863_),
    .B(_02860_),
    .Y(_02867_));
 sky130_fd_sc_hd__nand2_1 _09942_ (.A(_02866_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__nand2_1 _09943_ (.A(_06298_),
    .B(_06205_),
    .Y(_02869_));
 sky130_fd_sc_hd__nand3b_1 _09944_ (.A_N(_02869_),
    .B(_06247_),
    .C(_06215_),
    .Y(_02870_));
 sky130_fd_sc_hd__clkinv_4 _09945_ (.A(net14),
    .Y(_02871_));
 sky130_fd_sc_hd__o21ai_1 _09946_ (.A1(_02871_),
    .A2(_06331_),
    .B1(_02869_),
    .Y(_02872_));
 sky130_fd_sc_hd__nand2_1 _09947_ (.A(_02870_),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__nand2_1 _09948_ (.A(_02873_),
    .B(_00331_),
    .Y(_02874_));
 sky130_fd_sc_hd__nand3_1 _09949_ (.A(_02870_),
    .B(_06208_),
    .C(_02872_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _09950_ (.A(_02874_),
    .B(_02875_),
    .Y(_02877_));
 sky130_fd_sc_hd__a21oi_1 _09951_ (.A1(_02600_),
    .A2(_02605_),
    .B1(_02598_),
    .Y(_02878_));
 sky130_fd_sc_hd__inv_2 _09952_ (.A(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_1 _09953_ (.A(_06239_),
    .B(_00176_),
    .Y(_02880_));
 sky130_fd_sc_hd__nand2_1 _09954_ (.A(_06241_),
    .B(_06195_),
    .Y(_02881_));
 sky130_fd_sc_hd__nor2_1 _09955_ (.A(_02880_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__inv_2 _09956_ (.A(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nand2_1 _09957_ (.A(_02880_),
    .B(_02881_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_1 _09958_ (.A(_02883_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__nand2_1 _09959_ (.A(_02095_),
    .B(_06211_),
    .Y(_02886_));
 sky130_fd_sc_hd__nand2_1 _09960_ (.A(_02885_),
    .B(_02886_),
    .Y(_02888_));
 sky130_fd_sc_hd__inv_2 _09961_ (.A(_02886_),
    .Y(_02889_));
 sky130_fd_sc_hd__nand3_1 _09962_ (.A(_02883_),
    .B(_02889_),
    .C(_02884_),
    .Y(_02890_));
 sky130_fd_sc_hd__nand3_1 _09963_ (.A(_02879_),
    .B(_02888_),
    .C(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__nand2_1 _09964_ (.A(_02888_),
    .B(_02890_),
    .Y(_02892_));
 sky130_fd_sc_hd__nand2_1 _09965_ (.A(_02892_),
    .B(_02878_),
    .Y(_02893_));
 sky130_fd_sc_hd__nand3b_1 _09966_ (.A_N(_02877_),
    .B(_02891_),
    .C(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__nand2_1 _09967_ (.A(_02893_),
    .B(_02891_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_1 _09968_ (.A(_02895_),
    .B(_02877_),
    .Y(_02896_));
 sky130_fd_sc_hd__nand2_1 _09969_ (.A(_02894_),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__nand3_1 _09970_ (.A(_02864_),
    .B(_02868_),
    .C(_02897_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _09971_ (.A(_02864_),
    .B(_02868_),
    .Y(_02900_));
 sky130_fd_sc_hd__inv_2 _09972_ (.A(_02897_),
    .Y(_02901_));
 sky130_fd_sc_hd__nand2_1 _09973_ (.A(_02900_),
    .B(_02901_),
    .Y(_02902_));
 sky130_fd_sc_hd__nand3_1 _09974_ (.A(_02837_),
    .B(_02899_),
    .C(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__nand2_1 _09975_ (.A(_02902_),
    .B(_02899_),
    .Y(_02904_));
 sky130_fd_sc_hd__a21oi_1 _09976_ (.A1(_02835_),
    .A2(_02551_),
    .B1(_02836_),
    .Y(_02905_));
 sky130_fd_sc_hd__nand2_1 _09977_ (.A(_02904_),
    .B(_02905_),
    .Y(_02906_));
 sky130_fd_sc_hd__or2_1 _09978_ (.A(_02570_),
    .B(_02621_),
    .X(_02907_));
 sky130_fd_sc_hd__nand2_1 _09979_ (.A(_02626_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__nand3_1 _09980_ (.A(_02903_),
    .B(_02906_),
    .C(_02908_),
    .Y(_02910_));
 sky130_fd_sc_hd__nand2_1 _09981_ (.A(_02904_),
    .B(_02837_),
    .Y(_02911_));
 sky130_fd_sc_hd__nand3_1 _09982_ (.A(_02905_),
    .B(_02902_),
    .C(_02899_),
    .Y(_02912_));
 sky130_fd_sc_hd__inv_2 _09983_ (.A(_02908_),
    .Y(_02913_));
 sky130_fd_sc_hd__nand3_1 _09984_ (.A(_02911_),
    .B(_02912_),
    .C(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__nand2_1 _09985_ (.A(_02910_),
    .B(_02914_),
    .Y(_02915_));
 sky130_fd_sc_hd__nand3_1 _09986_ (.A(_02830_),
    .B(_02834_),
    .C(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__nand2_1 _09987_ (.A(_02830_),
    .B(_02834_),
    .Y(_02917_));
 sky130_fd_sc_hd__inv_2 _09988_ (.A(_02915_),
    .Y(_02918_));
 sky130_fd_sc_hd__nand2_1 _09989_ (.A(_02917_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__nand3_1 _09990_ (.A(_02685_),
    .B(_02916_),
    .C(_02919_),
    .Y(_02921_));
 sky130_fd_sc_hd__a21o_1 _09991_ (.A1(_02638_),
    .A2(_02683_),
    .B1(_02684_),
    .X(_02922_));
 sky130_fd_sc_hd__nand2_1 _09992_ (.A(_02919_),
    .B(_02916_),
    .Y(_02923_));
 sky130_fd_sc_hd__nand2_1 _09993_ (.A(_02922_),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_1 _09994_ (.A(_02921_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand2_1 _09995_ (.A(_02635_),
    .B(_02627_),
    .Y(_02926_));
 sky130_fd_sc_hd__nand2_1 _09996_ (.A(_02618_),
    .B(_02610_),
    .Y(_02927_));
 sky130_fd_sc_hd__nand2_1 _09997_ (.A(_02926_),
    .B(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__inv_2 _09998_ (.A(_02927_),
    .Y(_02929_));
 sky130_fd_sc_hd__nand3_1 _09999_ (.A(_02635_),
    .B(_02627_),
    .C(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__nand2_1 _10000_ (.A(_02928_),
    .B(_02930_),
    .Y(_02932_));
 sky130_fd_sc_hd__nand2_1 _10001_ (.A(_02932_),
    .B(_02613_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand3_1 _10002_ (.A(_02928_),
    .B(_02612_),
    .C(_02930_),
    .Y(_02934_));
 sky130_fd_sc_hd__nand2_1 _10003_ (.A(_02933_),
    .B(_02934_),
    .Y(_02935_));
 sky130_fd_sc_hd__inv_2 _10004_ (.A(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand2_1 _10005_ (.A(_02925_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand3_1 _10006_ (.A(_02921_),
    .B(_02924_),
    .C(_02935_),
    .Y(_02938_));
 sky130_fd_sc_hd__nand2_1 _10007_ (.A(_02937_),
    .B(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__nand2_1 _10008_ (.A(_02641_),
    .B(_02644_),
    .Y(_02940_));
 sky130_fd_sc_hd__nor2_1 _10009_ (.A(_02644_),
    .B(_02641_),
    .Y(_02941_));
 sky130_fd_sc_hd__a21oi_2 _10010_ (.A1(_02940_),
    .A2(_02656_),
    .B1(_02941_),
    .Y(_02943_));
 sky130_fd_sc_hd__inv_2 _10011_ (.A(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_1 _10012_ (.A(_02939_),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__nand3_1 _10013_ (.A(_02943_),
    .B(_02937_),
    .C(_02938_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand2_1 _10014_ (.A(_02945_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__nand2_1 _10015_ (.A(_02947_),
    .B(_02653_),
    .Y(_02948_));
 sky130_fd_sc_hd__nand3_1 _10016_ (.A(_02945_),
    .B(_02946_),
    .C(_02652_),
    .Y(_02949_));
 sky130_fd_sc_hd__nand2_1 _10017_ (.A(_02948_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__nand2_1 _10018_ (.A(_02660_),
    .B(_02663_),
    .Y(_02951_));
 sky130_fd_sc_hd__nor2_1 _10019_ (.A(_02663_),
    .B(_02660_),
    .Y(_02952_));
 sky130_fd_sc_hd__a21o_1 _10020_ (.A1(_02951_),
    .A2(_02172_),
    .B1(_02952_),
    .X(_02954_));
 sky130_fd_sc_hd__nand2_1 _10021_ (.A(_02950_),
    .B(_02954_),
    .Y(_02955_));
 sky130_fd_sc_hd__a21oi_1 _10022_ (.A1(_02951_),
    .A2(_02172_),
    .B1(_02952_),
    .Y(_02956_));
 sky130_fd_sc_hd__nand3_1 _10023_ (.A(_02956_),
    .B(_02948_),
    .C(_02949_),
    .Y(_02957_));
 sky130_fd_sc_hd__nand2_1 _10024_ (.A(_02955_),
    .B(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand2_1 _10025_ (.A(_02681_),
    .B(_02672_),
    .Y(_02959_));
 sky130_fd_sc_hd__xnor2_1 _10026_ (.A(_02958_),
    .B(_02959_),
    .Y(\m1.out[23] ));
 sky130_fd_sc_hd__nand2_1 _10027_ (.A(_01678_),
    .B(_02156_),
    .Y(_02960_));
 sky130_fd_sc_hd__nor2_1 _10028_ (.A(_02673_),
    .B(_02958_),
    .Y(_02961_));
 sky130_fd_sc_hd__nand2_1 _10029_ (.A(_02961_),
    .B(_02675_),
    .Y(_02962_));
 sky130_fd_sc_hd__nor2_2 _10030_ (.A(_02960_),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__nor2_1 _10031_ (.A(_02954_),
    .B(_02950_),
    .Y(_02964_));
 sky130_fd_sc_hd__o21ai_1 _10032_ (.A1(_02672_),
    .A2(_02964_),
    .B1(_02955_),
    .Y(_02965_));
 sky130_fd_sc_hd__a21oi_1 _10033_ (.A1(_02961_),
    .A2(_02677_),
    .B1(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__nand3_1 _10034_ (.A(_02161_),
    .B(_02675_),
    .C(_02961_),
    .Y(_02967_));
 sky130_fd_sc_hd__nand2_2 _10035_ (.A(_02966_),
    .B(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hd__a21oi_4 _10036_ (.A1(_01268_),
    .A2(_02963_),
    .B1(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__inv_2 _10037_ (.A(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__nand2_1 _10038_ (.A(_02939_),
    .B(_02943_),
    .Y(_02971_));
 sky130_fd_sc_hd__nor2_1 _10039_ (.A(_02943_),
    .B(_02939_),
    .Y(_02972_));
 sky130_fd_sc_hd__a21o_1 _10040_ (.A1(_02971_),
    .A2(_02652_),
    .B1(_02972_),
    .X(_02974_));
 sky130_fd_sc_hd__nand2_1 _10041_ (.A(_02923_),
    .B(_02685_),
    .Y(_02975_));
 sky130_fd_sc_hd__nor2_1 _10042_ (.A(_02685_),
    .B(_02923_),
    .Y(_02976_));
 sky130_fd_sc_hd__a21oi_1 _10043_ (.A1(_02975_),
    .A2(_02936_),
    .B1(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__nand2_1 _10044_ (.A(_02831_),
    .B(_02688_),
    .Y(_02978_));
 sky130_fd_sc_hd__nor2_1 _10045_ (.A(_02688_),
    .B(_02831_),
    .Y(_02979_));
 sky130_fd_sc_hd__a21oi_1 _10046_ (.A1(_02978_),
    .A2(_02918_),
    .B1(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hd__nand2_1 _10047_ (.A(_02772_),
    .B(_02692_),
    .Y(_02981_));
 sky130_fd_sc_hd__nor2_1 _10048_ (.A(_02692_),
    .B(_02772_),
    .Y(_02982_));
 sky130_fd_sc_hd__a21oi_1 _10049_ (.A1(_02981_),
    .A2(_02828_),
    .B1(_02982_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2_1 _10050_ (.A(_06276_),
    .B(_06184_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand2_1 _10051_ (.A(_02985_),
    .B(_06328_),
    .Y(_02986_));
 sky130_fd_sc_hd__nand3_1 _10052_ (.A(_06269_),
    .B(_06276_),
    .C(_06184_),
    .Y(_02987_));
 sky130_fd_sc_hd__nand2_1 _10053_ (.A(_02986_),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hd__nand2_1 _10054_ (.A(_06274_),
    .B(_02181_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand2_1 _10055_ (.A(_02988_),
    .B(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__inv_2 _10056_ (.A(_02989_),
    .Y(_02991_));
 sky130_fd_sc_hd__nand3_1 _10057_ (.A(_02986_),
    .B(_02987_),
    .C(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__nand2_1 _10058_ (.A(_02990_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__inv_2 _10059_ (.A(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__a21boi_2 _10060_ (.A1(_02699_),
    .A2(_02705_),
    .B1_N(_02700_),
    .Y(_02996_));
 sky130_fd_sc_hd__inv_2 _10061_ (.A(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__nand2_1 _10062_ (.A(_02994_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand2_1 _10063_ (.A(_06259_),
    .B(_01692_),
    .Y(_02999_));
 sky130_fd_sc_hd__inv_2 _10064_ (.A(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__nand2_1 _10065_ (.A(_06261_),
    .B(_01921_),
    .Y(_03001_));
 sky130_fd_sc_hd__inv_2 _10066_ (.A(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__nand2_1 _10067_ (.A(_03000_),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2_1 _10068_ (.A(_02999_),
    .B(_03001_),
    .Y(_03004_));
 sky130_fd_sc_hd__nand2_1 _10069_ (.A(_03003_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__nand2_1 _10070_ (.A(_06266_),
    .B(_06177_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _10071_ (.A(_03005_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__inv_2 _10072_ (.A(_03007_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand3_1 _10073_ (.A(_03003_),
    .B(_03009_),
    .C(_03004_),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2_1 _10074_ (.A(_03008_),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__inv_2 _10075_ (.A(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__nand2_1 _10076_ (.A(_02993_),
    .B(_02996_),
    .Y(_03013_));
 sky130_fd_sc_hd__nand3_1 _10077_ (.A(_02998_),
    .B(_03012_),
    .C(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_1 _10078_ (.A(_02994_),
    .B(_02996_),
    .Y(_03015_));
 sky130_fd_sc_hd__nand2_1 _10079_ (.A(_02997_),
    .B(_02993_),
    .Y(_03016_));
 sky130_fd_sc_hd__nand3_1 _10080_ (.A(_03015_),
    .B(_03016_),
    .C(_03011_),
    .Y(_03018_));
 sky130_fd_sc_hd__nand2_1 _10081_ (.A(_03014_),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__nor2_1 _10082_ (.A(_02697_),
    .B(_02709_),
    .Y(_03020_));
 sky130_fd_sc_hd__a21oi_2 _10083_ (.A1(_02729_),
    .A2(_02730_),
    .B1(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__inv_2 _10084_ (.A(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__nand2_1 _10085_ (.A(_03019_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__nand3_1 _10086_ (.A(_03021_),
    .B(_03018_),
    .C(_03014_),
    .Y(_03024_));
 sky130_fd_sc_hd__nand2_1 _10087_ (.A(_03023_),
    .B(_03024_),
    .Y(_03025_));
 sky130_fd_sc_hd__nand2_1 _10088_ (.A(_06289_),
    .B(_06173_),
    .Y(_03026_));
 sky130_fd_sc_hd__inv_2 _10089_ (.A(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__nand2_1 _10090_ (.A(_00299_),
    .B(_01280_),
    .Y(_03029_));
 sky130_fd_sc_hd__inv_2 _10091_ (.A(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand2_1 _10092_ (.A(_03027_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__nand2_1 _10093_ (.A(_03026_),
    .B(_03029_),
    .Y(_03032_));
 sky130_fd_sc_hd__nand2_1 _10094_ (.A(_03031_),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__nand2_1 _10095_ (.A(_06288_),
    .B(_00918_),
    .Y(_03034_));
 sky130_fd_sc_hd__nand2_1 _10096_ (.A(_03033_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__nand3b_2 _10097_ (.A_N(_03034_),
    .B(_03031_),
    .C(_03032_),
    .Y(_03036_));
 sky130_fd_sc_hd__nand2_1 _10098_ (.A(_03035_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__nor2_1 _10099_ (.A(_02714_),
    .B(_02711_),
    .Y(_03038_));
 sky130_fd_sc_hd__a21oi_1 _10100_ (.A1(_02722_),
    .A2(_02721_),
    .B1(_03038_),
    .Y(_03040_));
 sky130_fd_sc_hd__nand2_1 _10101_ (.A(_03037_),
    .B(_03040_),
    .Y(_03041_));
 sky130_fd_sc_hd__a21o_1 _10102_ (.A1(_02722_),
    .A2(_02721_),
    .B1(_03038_),
    .X(_03042_));
 sky130_fd_sc_hd__nand3_1 _10103_ (.A(_03042_),
    .B(_03036_),
    .C(_03035_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand2_1 _10104_ (.A(_02751_),
    .B(_02748_),
    .Y(_03044_));
 sky130_fd_sc_hd__nand3_1 _10105_ (.A(_03041_),
    .B(_03043_),
    .C(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__nand2_1 _10106_ (.A(_03037_),
    .B(_03042_),
    .Y(_03046_));
 sky130_fd_sc_hd__nand3_1 _10107_ (.A(_03035_),
    .B(_03036_),
    .C(_03040_),
    .Y(_03047_));
 sky130_fd_sc_hd__inv_2 _10108_ (.A(_03044_),
    .Y(_03048_));
 sky130_fd_sc_hd__nand3_1 _10109_ (.A(_03046_),
    .B(_03047_),
    .C(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__nand2_1 _10110_ (.A(_03045_),
    .B(_03049_),
    .Y(_03051_));
 sky130_fd_sc_hd__inv_2 _10111_ (.A(_03051_),
    .Y(_03052_));
 sky130_fd_sc_hd__nand2_1 _10112_ (.A(_03025_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand3_2 _10113_ (.A(_03023_),
    .B(_03024_),
    .C(_03051_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand2_1 _10114_ (.A(_03053_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__nor2_1 _10115_ (.A(_02695_),
    .B(_02735_),
    .Y(_03056_));
 sky130_fd_sc_hd__a21oi_2 _10116_ (.A1(_02769_),
    .A2(_02768_),
    .B1(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__inv_2 _10117_ (.A(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__nand2_1 _10118_ (.A(_03055_),
    .B(_03058_),
    .Y(_03059_));
 sky130_fd_sc_hd__nand3_1 _10119_ (.A(_03057_),
    .B(_03053_),
    .C(_03054_),
    .Y(_03060_));
 sky130_fd_sc_hd__nor2_1 _10120_ (.A(_02754_),
    .B(_02753_),
    .Y(_03062_));
 sky130_fd_sc_hd__a21oi_1 _10121_ (.A1(_02755_),
    .A2(_02757_),
    .B1(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__nand2_1 _10122_ (.A(_00561_),
    .B(_00926_),
    .Y(_03064_));
 sky130_fd_sc_hd__inv_2 _10123_ (.A(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__nand2_1 _10124_ (.A(_00439_),
    .B(_00921_),
    .Y(_03066_));
 sky130_fd_sc_hd__nand2_1 _10125_ (.A(_03065_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__inv_2 _10126_ (.A(_03066_),
    .Y(_03068_));
 sky130_fd_sc_hd__nand2_1 _10127_ (.A(_03068_),
    .B(_03064_),
    .Y(_03069_));
 sky130_fd_sc_hd__nand2_1 _10128_ (.A(net4),
    .B(_06219_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand3_2 _10129_ (.A(_03067_),
    .B(_03069_),
    .C(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__nand2_1 _10130_ (.A(_03065_),
    .B(_03068_),
    .Y(_03073_));
 sky130_fd_sc_hd__inv_2 _10131_ (.A(_03070_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _10132_ (.A(_03064_),
    .B(_03066_),
    .Y(_03075_));
 sky130_fd_sc_hd__nand3_2 _10133_ (.A(_03073_),
    .B(_03074_),
    .C(_03075_),
    .Y(_03076_));
 sky130_fd_sc_hd__nand2_1 _10134_ (.A(_03071_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__nor2_1 _10135_ (.A(_02779_),
    .B(_02781_),
    .Y(_03078_));
 sky130_fd_sc_hd__a21oi_2 _10136_ (.A1(_02790_),
    .A2(_02788_),
    .B1(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__inv_2 _10137_ (.A(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__nand2_1 _10138_ (.A(_03077_),
    .B(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__nand3_1 _10139_ (.A(_03079_),
    .B(_03071_),
    .C(_03076_),
    .Y(_03082_));
 sky130_fd_sc_hd__nand2_1 _10140_ (.A(_01158_),
    .B(_06230_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2_1 _10141_ (.A(_00701_),
    .B(_00376_),
    .Y(_03085_));
 sky130_fd_sc_hd__nor2_1 _10142_ (.A(_03084_),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__nand2_1 _10143_ (.A(_03084_),
    .B(_03085_),
    .Y(_03087_));
 sky130_fd_sc_hd__inv_2 _10144_ (.A(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__nand2_1 _10145_ (.A(_06281_),
    .B(_00780_),
    .Y(_03089_));
 sky130_fd_sc_hd__o21ai_1 _10146_ (.A1(_03086_),
    .A2(_03088_),
    .B1(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__inv_2 _10147_ (.A(_03089_),
    .Y(_03091_));
 sky130_fd_sc_hd__nand3b_1 _10148_ (.A_N(_03086_),
    .B(_03091_),
    .C(_03087_),
    .Y(_03092_));
 sky130_fd_sc_hd__nand2_1 _10149_ (.A(_03090_),
    .B(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__nand3_1 _10150_ (.A(_03081_),
    .B(_03082_),
    .C(_03093_),
    .Y(_03095_));
 sky130_fd_sc_hd__nand2_1 _10151_ (.A(_03081_),
    .B(_03082_),
    .Y(_03096_));
 sky130_fd_sc_hd__inv_2 _10152_ (.A(_03093_),
    .Y(_03097_));
 sky130_fd_sc_hd__nand2_1 _10153_ (.A(_03096_),
    .B(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__nand3_1 _10154_ (.A(_03063_),
    .B(_03095_),
    .C(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_03098_),
    .B(_03095_),
    .Y(_03100_));
 sky130_fd_sc_hd__nand2_1 _10156_ (.A(_02758_),
    .B(_02752_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _10157_ (.A(_03100_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__nand2_1 _10158_ (.A(_03099_),
    .B(_03102_),
    .Y(_03103_));
 sky130_fd_sc_hd__nand2_1 _10159_ (.A(_02815_),
    .B(_02812_),
    .Y(_03104_));
 sky130_fd_sc_hd__nand2_1 _10160_ (.A(_03103_),
    .B(_03104_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand3b_1 _10161_ (.A_N(_03104_),
    .B(_03099_),
    .C(_03102_),
    .Y(_03107_));
 sky130_fd_sc_hd__nand2_2 _10162_ (.A(_03106_),
    .B(_03107_),
    .Y(_03108_));
 sky130_fd_sc_hd__nand3_2 _10163_ (.A(_03059_),
    .B(_03060_),
    .C(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__nand2_1 _10164_ (.A(_03059_),
    .B(_03060_),
    .Y(_03110_));
 sky130_fd_sc_hd__inv_2 _10165_ (.A(_03108_),
    .Y(_03111_));
 sky130_fd_sc_hd__nand2_1 _10166_ (.A(_03110_),
    .B(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__nand3_1 _10167_ (.A(_02983_),
    .B(_03109_),
    .C(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _10168_ (.A(_03112_),
    .B(_03109_),
    .Y(_03114_));
 sky130_fd_sc_hd__a21o_1 _10169_ (.A1(_02981_),
    .A2(_02828_),
    .B1(_02982_),
    .X(_03115_));
 sky130_fd_sc_hd__nand2_1 _10170_ (.A(_03114_),
    .B(_03115_),
    .Y(_03117_));
 sky130_fd_sc_hd__nand2_1 _10171_ (.A(_02818_),
    .B(_02777_),
    .Y(_03118_));
 sky130_fd_sc_hd__nor2_1 _10172_ (.A(_02777_),
    .B(_02818_),
    .Y(_03119_));
 sky130_fd_sc_hd__a21oi_2 _10173_ (.A1(_03118_),
    .A2(_02822_),
    .B1(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__inv_2 _10174_ (.A(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__inv_2 _10175_ (.A(_02862_),
    .Y(_03122_));
 sky130_fd_sc_hd__a21oi_1 _10176_ (.A1(_02861_),
    .A2(_02858_),
    .B1(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__nand2_1 _10177_ (.A(_02850_),
    .B(_02845_),
    .Y(_03124_));
 sky130_fd_sc_hd__nand2_1 _10178_ (.A(_06235_),
    .B(_06200_),
    .Y(_03125_));
 sky130_fd_sc_hd__inv_2 _10179_ (.A(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__nand2_1 _10180_ (.A(_01211_),
    .B(_06226_),
    .Y(_03128_));
 sky130_fd_sc_hd__inv_2 _10181_ (.A(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_1 _10182_ (.A(_03126_),
    .B(_03129_),
    .Y(_03130_));
 sky130_fd_sc_hd__nand2_1 _10183_ (.A(_03125_),
    .B(_03128_),
    .Y(_03131_));
 sky130_fd_sc_hd__nand2_1 _10184_ (.A(_03130_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__nand2_1 _10185_ (.A(_06243_),
    .B(_06202_),
    .Y(_03133_));
 sky130_fd_sc_hd__nand2_1 _10186_ (.A(_03132_),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hd__nand3b_1 _10187_ (.A_N(_03133_),
    .B(_03130_),
    .C(_03131_),
    .Y(_03135_));
 sky130_fd_sc_hd__nand2_1 _10188_ (.A(_03134_),
    .B(_03135_),
    .Y(_03136_));
 sky130_fd_sc_hd__nor2_1 _10189_ (.A(_02798_),
    .B(_02800_),
    .Y(_03137_));
 sky130_fd_sc_hd__a21oi_2 _10190_ (.A1(_02803_),
    .A2(_02807_),
    .B1(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__inv_2 _10191_ (.A(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__nand2_1 _10192_ (.A(_03136_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hd__nand3_1 _10193_ (.A(_03134_),
    .B(_03135_),
    .C(_03138_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand3b_1 _10194_ (.A_N(_03124_),
    .B(_03140_),
    .C(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2_1 _10195_ (.A(_03140_),
    .B(_03141_),
    .Y(_03143_));
 sky130_fd_sc_hd__nand2_1 _10196_ (.A(_03143_),
    .B(_03124_),
    .Y(_03144_));
 sky130_fd_sc_hd__nand3_1 _10197_ (.A(_03123_),
    .B(_03142_),
    .C(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__nand2_1 _10198_ (.A(_03144_),
    .B(_03142_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand2_1 _10199_ (.A(_02863_),
    .B(_02862_),
    .Y(_03147_));
 sky130_fd_sc_hd__nand2_1 _10200_ (.A(_03146_),
    .B(_03147_),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _10201_ (.A(_02095_),
    .B(_00176_),
    .Y(_03150_));
 sky130_fd_sc_hd__nand2_1 _10202_ (.A(_01858_),
    .B(_06196_),
    .Y(_03151_));
 sky130_fd_sc_hd__or2_1 _10203_ (.A(_03150_),
    .B(_03151_),
    .X(_03152_));
 sky130_fd_sc_hd__nand2_1 _10204_ (.A(_03150_),
    .B(_03151_),
    .Y(_03153_));
 sky130_fd_sc_hd__nand2_1 _10205_ (.A(_03152_),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__nand2_1 _10206_ (.A(_06245_),
    .B(_06211_),
    .Y(_03155_));
 sky130_fd_sc_hd__nand2_1 _10207_ (.A(_03154_),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__nand3b_1 _10208_ (.A_N(_03155_),
    .B(_03152_),
    .C(_03153_),
    .Y(_03157_));
 sky130_fd_sc_hd__nand2_1 _10209_ (.A(_03156_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__nand2_1 _10210_ (.A(_02890_),
    .B(_02883_),
    .Y(_03160_));
 sky130_fd_sc_hd__inv_2 _10211_ (.A(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__nand2_1 _10212_ (.A(_03158_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__nand3_1 _10213_ (.A(_03160_),
    .B(_03156_),
    .C(_03157_),
    .Y(_03163_));
 sky130_fd_sc_hd__nand2_1 _10214_ (.A(_03162_),
    .B(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hd__and3_1 _10215_ (.A(_06298_),
    .B(_06205_),
    .C(_06214_),
    .X(_03165_));
 sky130_fd_sc_hd__inv_2 _10216_ (.A(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__a21o_1 _10217_ (.A1(_06299_),
    .A2(_06215_),
    .B1(_06206_),
    .X(_03167_));
 sky130_fd_sc_hd__nand2_1 _10218_ (.A(_03166_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand2_1 _10219_ (.A(_03164_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__nand3b_1 _10220_ (.A_N(_03168_),
    .B(_03162_),
    .C(_03163_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _10221_ (.A(_03169_),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand3_1 _10222_ (.A(_03145_),
    .B(_03149_),
    .C(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__nand2_1 _10223_ (.A(_03145_),
    .B(_03149_),
    .Y(_03174_));
 sky130_fd_sc_hd__inv_2 _10224_ (.A(_03172_),
    .Y(_03175_));
 sky130_fd_sc_hd__nand2_1 _10225_ (.A(_03174_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand3_2 _10226_ (.A(_03121_),
    .B(_03173_),
    .C(_03176_),
    .Y(_03177_));
 sky130_fd_sc_hd__nand2_1 _10227_ (.A(_03176_),
    .B(_03173_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_1 _10228_ (.A(_03178_),
    .B(_03120_),
    .Y(_03179_));
 sky130_fd_sc_hd__nand2_1 _10229_ (.A(_03177_),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__o21ai_1 _10230_ (.A1(_02839_),
    .A2(_02867_),
    .B1(_02902_),
    .Y(_03182_));
 sky130_fd_sc_hd__inv_2 _10231_ (.A(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2_1 _10232_ (.A(_03180_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__nand3_1 _10233_ (.A(_03177_),
    .B(_03179_),
    .C(_03182_),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_2 _10234_ (.A(_03184_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__nand3_1 _10235_ (.A(_03113_),
    .B(_03117_),
    .C(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_1 _10236_ (.A(_03113_),
    .B(_03117_),
    .Y(_03188_));
 sky130_fd_sc_hd__inv_2 _10237_ (.A(_03186_),
    .Y(_03189_));
 sky130_fd_sc_hd__nand2_1 _10238_ (.A(_03188_),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__nand3_1 _10239_ (.A(_02980_),
    .B(_03187_),
    .C(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__nand2_1 _10240_ (.A(_03190_),
    .B(_03187_),
    .Y(_03193_));
 sky130_fd_sc_hd__a21o_1 _10241_ (.A1(_02978_),
    .A2(_02918_),
    .B1(_02979_),
    .X(_03194_));
 sky130_fd_sc_hd__nand2_1 _10242_ (.A(_03193_),
    .B(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__nand2_1 _10243_ (.A(_02910_),
    .B(_02903_),
    .Y(_03196_));
 sky130_fd_sc_hd__nand2_1 _10244_ (.A(_02894_),
    .B(_02891_),
    .Y(_03197_));
 sky130_fd_sc_hd__nand2_1 _10245_ (.A(_03196_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__inv_2 _10246_ (.A(_03197_),
    .Y(_03199_));
 sky130_fd_sc_hd__nand3_1 _10247_ (.A(_02910_),
    .B(_02903_),
    .C(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__nand2_1 _10248_ (.A(_03198_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__nand2_1 _10249_ (.A(_02875_),
    .B(_02870_),
    .Y(_03202_));
 sky130_fd_sc_hd__inv_2 _10250_ (.A(_03202_),
    .Y(_03204_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(_03201_),
    .B(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand3_1 _10252_ (.A(_03198_),
    .B(_03202_),
    .C(_03200_),
    .Y(_03206_));
 sky130_fd_sc_hd__nand2_1 _10253_ (.A(_03205_),
    .B(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__nand3_1 _10254_ (.A(_03191_),
    .B(_03195_),
    .C(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__nand2_1 _10255_ (.A(_03191_),
    .B(_03195_),
    .Y(_03209_));
 sky130_fd_sc_hd__inv_2 _10256_ (.A(_03207_),
    .Y(_03210_));
 sky130_fd_sc_hd__nand2_1 _10257_ (.A(_03209_),
    .B(_03210_),
    .Y(_03211_));
 sky130_fd_sc_hd__nand3_1 _10258_ (.A(_02977_),
    .B(_03208_),
    .C(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _10259_ (.A(_03211_),
    .B(_03208_),
    .Y(_03213_));
 sky130_fd_sc_hd__a21o_1 _10260_ (.A1(_02975_),
    .A2(_02936_),
    .B1(_02976_),
    .X(_03215_));
 sky130_fd_sc_hd__nand2_1 _10261_ (.A(_03213_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__nand2_2 _10262_ (.A(_02934_),
    .B(_02928_),
    .Y(_03217_));
 sky130_fd_sc_hd__inv_2 _10263_ (.A(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__nand3_1 _10264_ (.A(_03212_),
    .B(_03216_),
    .C(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__nand2_1 _10265_ (.A(_03212_),
    .B(_03216_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand2_1 _10266_ (.A(_03220_),
    .B(_03217_),
    .Y(_03221_));
 sky130_fd_sc_hd__nand3_1 _10267_ (.A(_02974_),
    .B(_03219_),
    .C(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__nand2_1 _10268_ (.A(_03221_),
    .B(_03219_),
    .Y(_03223_));
 sky130_fd_sc_hd__a21oi_1 _10269_ (.A1(_02971_),
    .A2(_02652_),
    .B1(_02972_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand2_1 _10270_ (.A(_03223_),
    .B(_03224_),
    .Y(_03226_));
 sky130_fd_sc_hd__nand2_1 _10271_ (.A(_03222_),
    .B(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__inv_2 _10272_ (.A(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_1 _10273_ (.A(_02970_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand2_1 _10274_ (.A(_02969_),
    .B(_03227_),
    .Y(_03230_));
 sky130_fd_sc_hd__and2_1 _10275_ (.A(_03229_),
    .B(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__clkbuf_1 _10276_ (.A(_03231_),
    .X(\m1.out[24] ));
 sky130_fd_sc_hd__nand2_1 _10277_ (.A(_03213_),
    .B(_02977_),
    .Y(_03232_));
 sky130_fd_sc_hd__nor2_1 _10278_ (.A(_02977_),
    .B(_03213_),
    .Y(_03233_));
 sky130_fd_sc_hd__a21oi_1 _10279_ (.A1(_03232_),
    .A2(_03217_),
    .B1(_03233_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_1 _10280_ (.A(_03114_),
    .B(_02983_),
    .Y(_03236_));
 sky130_fd_sc_hd__inv_2 _10281_ (.A(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__nor2_1 _10282_ (.A(_02983_),
    .B(_03114_),
    .Y(_03238_));
 sky130_fd_sc_hd__o21bai_1 _10283_ (.A1(_03186_),
    .A2(_03237_),
    .B1_N(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__nand2_1 _10284_ (.A(_03055_),
    .B(_03057_),
    .Y(_03240_));
 sky130_fd_sc_hd__nor2_1 _10285_ (.A(_03057_),
    .B(_03055_),
    .Y(_03241_));
 sky130_fd_sc_hd__a21oi_1 _10286_ (.A1(_03240_),
    .A2(_03111_),
    .B1(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__nand2_1 _10287_ (.A(_03019_),
    .B(_03021_),
    .Y(_03243_));
 sky130_fd_sc_hd__nor2_1 _10288_ (.A(_03021_),
    .B(_03019_),
    .Y(_03244_));
 sky130_fd_sc_hd__a21oi_1 _10289_ (.A1(_03243_),
    .A2(_03052_),
    .B1(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__nor2_1 _10290_ (.A(_02996_),
    .B(_02993_),
    .Y(_03247_));
 sky130_fd_sc_hd__a21oi_1 _10291_ (.A1(_03012_),
    .A2(_03013_),
    .B1(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__nand2_1 _10292_ (.A(_06274_),
    .B(_02423_),
    .Y(_03249_));
 sky130_fd_sc_hd__inv_2 _10293_ (.A(_06392_),
    .Y(_03250_));
 sky130_fd_sc_hd__nand2_1 _10294_ (.A(_03249_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand3_2 _10295_ (.A(_06273_),
    .B(_06392_),
    .C(_06183_),
    .Y(_03252_));
 sky130_fd_sc_hd__nand2_1 _10296_ (.A(_03251_),
    .B(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__nand2_1 _10297_ (.A(_06261_),
    .B(_02180_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand2_1 _10298_ (.A(_03253_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__inv_2 _10299_ (.A(_03254_),
    .Y(_03256_));
 sky130_fd_sc_hd__nand3_1 _10300_ (.A(_03251_),
    .B(_03252_),
    .C(_03256_),
    .Y(_03258_));
 sky130_fd_sc_hd__nand2_2 _10301_ (.A(_03255_),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__inv_4 _10302_ (.A(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__a21boi_1 _10303_ (.A1(_02986_),
    .A2(_02991_),
    .B1_N(_02987_),
    .Y(_03261_));
 sky130_fd_sc_hd__nand2_1 _10304_ (.A(_03260_),
    .B(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _10305_ (.A(_06265_),
    .B(_06175_),
    .Y(_03263_));
 sky130_fd_sc_hd__inv_2 _10306_ (.A(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__nand2_1 _10307_ (.A(_00175_),
    .B(_06187_),
    .Y(_03265_));
 sky130_fd_sc_hd__inv_2 _10308_ (.A(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__nand2_1 _10309_ (.A(_03264_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand2_1 _10310_ (.A(_03263_),
    .B(_03265_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(_03267_),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hd__nand2_1 _10312_ (.A(_00299_),
    .B(_06177_),
    .Y(_03271_));
 sky130_fd_sc_hd__nand2_1 _10313_ (.A(_03270_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__inv_2 _10314_ (.A(_03271_),
    .Y(_03273_));
 sky130_fd_sc_hd__nand3_1 _10315_ (.A(_03267_),
    .B(_03273_),
    .C(_03269_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_1 _10316_ (.A(_03272_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__nand2_1 _10317_ (.A(_02992_),
    .B(_02987_),
    .Y(_03276_));
 sky130_fd_sc_hd__nand2_1 _10318_ (.A(_03259_),
    .B(_03276_),
    .Y(_03277_));
 sky130_fd_sc_hd__nand3_1 _10319_ (.A(_03262_),
    .B(_03275_),
    .C(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__nand2_1 _10320_ (.A(_03260_),
    .B(_03276_),
    .Y(_03280_));
 sky130_fd_sc_hd__inv_2 _10321_ (.A(_03275_),
    .Y(_03281_));
 sky130_fd_sc_hd__nand2_1 _10322_ (.A(_03259_),
    .B(_03261_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand3_2 _10323_ (.A(_03280_),
    .B(_03281_),
    .C(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__nand3_1 _10324_ (.A(_03248_),
    .B(_03278_),
    .C(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__nand2_1 _10325_ (.A(_03283_),
    .B(_03278_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _10326_ (.A(_03014_),
    .B(_02998_),
    .Y(_03286_));
 sky130_fd_sc_hd__nand2_1 _10327_ (.A(_03285_),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2_1 _10328_ (.A(_06287_),
    .B(_06173_),
    .Y(_03288_));
 sky130_fd_sc_hd__inv_2 _10329_ (.A(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__nand2_1 _10330_ (.A(_00193_),
    .B(_01280_),
    .Y(_03291_));
 sky130_fd_sc_hd__inv_2 _10331_ (.A(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__nand2_1 _10332_ (.A(_03289_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__nand2_1 _10333_ (.A(_03288_),
    .B(_03291_),
    .Y(_03294_));
 sky130_fd_sc_hd__nand2_1 _10334_ (.A(_03293_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__nand2_1 _10335_ (.A(_06292_),
    .B(_06222_),
    .Y(_03296_));
 sky130_fd_sc_hd__nand2_1 _10336_ (.A(_03295_),
    .B(_03296_),
    .Y(_03297_));
 sky130_fd_sc_hd__nand3b_2 _10337_ (.A_N(_03296_),
    .B(_03293_),
    .C(_03294_),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2_1 _10338_ (.A(_03297_),
    .B(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__nor2_1 _10339_ (.A(_02999_),
    .B(_03001_),
    .Y(_03300_));
 sky130_fd_sc_hd__a21oi_2 _10340_ (.A1(_03004_),
    .A2(_03009_),
    .B1(_03300_),
    .Y(_03302_));
 sky130_fd_sc_hd__inv_2 _10341_ (.A(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__nand2_1 _10342_ (.A(_03299_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__nand3_1 _10343_ (.A(_03297_),
    .B(_03298_),
    .C(_03302_),
    .Y(_03305_));
 sky130_fd_sc_hd__nand2_1 _10344_ (.A(_03304_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__nand2_1 _10345_ (.A(_03036_),
    .B(_03031_),
    .Y(_03307_));
 sky130_fd_sc_hd__nand2_1 _10346_ (.A(_03306_),
    .B(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__nand3b_1 _10347_ (.A_N(_03307_),
    .B(_03304_),
    .C(_03305_),
    .Y(_03309_));
 sky130_fd_sc_hd__nand2_1 _10348_ (.A(_03308_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__nand3_1 _10349_ (.A(_03284_),
    .B(_03287_),
    .C(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__nand3_1 _10350_ (.A(_03286_),
    .B(_03278_),
    .C(_03283_),
    .Y(_03312_));
 sky130_fd_sc_hd__inv_2 _10351_ (.A(_03310_),
    .Y(_03313_));
 sky130_fd_sc_hd__nand2_1 _10352_ (.A(_03285_),
    .B(_03248_),
    .Y(_03314_));
 sky130_fd_sc_hd__nand3_1 _10353_ (.A(_03312_),
    .B(_03313_),
    .C(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__nand3_1 _10354_ (.A(_03245_),
    .B(_03311_),
    .C(_03315_),
    .Y(_03316_));
 sky130_fd_sc_hd__nand2_1 _10355_ (.A(_03315_),
    .B(_03311_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21o_1 _10356_ (.A1(_03243_),
    .A2(_03052_),
    .B1(_03244_),
    .X(_03318_));
 sky130_fd_sc_hd__nand2_1 _10357_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__inv_2 _10358_ (.A(_03043_),
    .Y(_03320_));
 sky130_fd_sc_hd__a21oi_2 _10359_ (.A1(_03041_),
    .A2(_03044_),
    .B1(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__nor2_1 _10360_ (.A(_03064_),
    .B(_03066_),
    .Y(_03323_));
 sky130_fd_sc_hd__a21oi_2 _10361_ (.A1(_03075_),
    .A2(_03074_),
    .B1(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__inv_2 _10362_ (.A(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__nand2_1 _10363_ (.A(_00849_),
    .B(_00926_),
    .Y(_03326_));
 sky130_fd_sc_hd__inv_2 _10364_ (.A(_03326_),
    .Y(_03327_));
 sky130_fd_sc_hd__nand2_1 _10365_ (.A(_00561_),
    .B(_00921_),
    .Y(_03328_));
 sky130_fd_sc_hd__inv_2 _10366_ (.A(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _10367_ (.A(_03327_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand2_1 _10368_ (.A(_06278_),
    .B(_06219_),
    .Y(_03331_));
 sky130_fd_sc_hd__inv_2 _10369_ (.A(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand2_1 _10370_ (.A(_03326_),
    .B(_03328_),
    .Y(_03334_));
 sky130_fd_sc_hd__nand3_1 _10371_ (.A(_03330_),
    .B(_03332_),
    .C(_03334_),
    .Y(_03335_));
 sky130_fd_sc_hd__nand2_1 _10372_ (.A(_03330_),
    .B(_03334_),
    .Y(_03336_));
 sky130_fd_sc_hd__nand2_1 _10373_ (.A(_03336_),
    .B(_03331_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand3_1 _10374_ (.A(_03325_),
    .B(_03335_),
    .C(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _10375_ (.A(_03337_),
    .B(_03335_),
    .Y(_03339_));
 sky130_fd_sc_hd__nand2_1 _10376_ (.A(_03339_),
    .B(_03324_),
    .Y(_03340_));
 sky130_fd_sc_hd__nand2_1 _10377_ (.A(_03338_),
    .B(_03340_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand2_1 _10378_ (.A(_06281_),
    .B(_06230_),
    .Y(_03342_));
 sky130_fd_sc_hd__inv_2 _10379_ (.A(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2_1 _10380_ (.A(_06283_),
    .B(_06227_),
    .Y(_03345_));
 sky130_fd_sc_hd__inv_2 _10381_ (.A(_03345_),
    .Y(_03346_));
 sky130_fd_sc_hd__nand2_1 _10382_ (.A(_03343_),
    .B(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hd__nand2_1 _10383_ (.A(_03342_),
    .B(_03345_),
    .Y(_03348_));
 sky130_fd_sc_hd__nand2_1 _10384_ (.A(_03347_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_1 _10385_ (.A(_01211_),
    .B(_00780_),
    .Y(_03350_));
 sky130_fd_sc_hd__nand2_1 _10386_ (.A(_03349_),
    .B(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hd__inv_2 _10387_ (.A(_03350_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand3_1 _10388_ (.A(_03347_),
    .B(_03352_),
    .C(_03348_),
    .Y(_03353_));
 sky130_fd_sc_hd__nand2_1 _10389_ (.A(_03351_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__nand2_1 _10390_ (.A(_03341_),
    .B(_03354_),
    .Y(_03356_));
 sky130_fd_sc_hd__nand3b_2 _10391_ (.A_N(_03354_),
    .B(_03338_),
    .C(_03340_),
    .Y(_03357_));
 sky130_fd_sc_hd__nand3_1 _10392_ (.A(_03321_),
    .B(_03356_),
    .C(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__inv_2 _10393_ (.A(_03321_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand2_1 _10394_ (.A(_03356_),
    .B(_03357_),
    .Y(_03360_));
 sky130_fd_sc_hd__nand2_1 _10395_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__nand2_1 _10396_ (.A(_03358_),
    .B(_03361_),
    .Y(_03362_));
 sky130_fd_sc_hd__o21ai_2 _10397_ (.A1(_03079_),
    .A2(_03077_),
    .B1(_03098_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand2_1 _10398_ (.A(_03362_),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand3b_1 _10399_ (.A_N(_03363_),
    .B(_03358_),
    .C(_03361_),
    .Y(_03365_));
 sky130_fd_sc_hd__nand2_1 _10400_ (.A(_03364_),
    .B(_03365_),
    .Y(_03367_));
 sky130_fd_sc_hd__nand3_2 _10401_ (.A(_03316_),
    .B(_03319_),
    .C(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _10402_ (.A(_03316_),
    .B(_03319_),
    .Y(_03369_));
 sky130_fd_sc_hd__inv_2 _10403_ (.A(_03367_),
    .Y(_03370_));
 sky130_fd_sc_hd__nand2_2 _10404_ (.A(_03369_),
    .B(_03370_),
    .Y(_03371_));
 sky130_fd_sc_hd__nand3_1 _10405_ (.A(_03242_),
    .B(_03368_),
    .C(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand2_1 _10406_ (.A(_03371_),
    .B(_03368_),
    .Y(_03373_));
 sky130_fd_sc_hd__a21o_1 _10407_ (.A1(_03240_),
    .A2(_03111_),
    .B1(_03241_),
    .X(_03374_));
 sky130_fd_sc_hd__nand2_1 _10408_ (.A(_03373_),
    .B(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__nand2_1 _10409_ (.A(_06241_),
    .B(_06200_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _10410_ (.A(_06235_),
    .B(_06226_),
    .Y(_03378_));
 sky130_fd_sc_hd__nor2_1 _10411_ (.A(_03376_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__nand2_1 _10412_ (.A(_03376_),
    .B(_03378_),
    .Y(_03380_));
 sky130_fd_sc_hd__inv_2 _10413_ (.A(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__nand2_1 _10414_ (.A(_06240_),
    .B(_06202_),
    .Y(_03382_));
 sky130_fd_sc_hd__o21ai_1 _10415_ (.A1(_03379_),
    .A2(_03381_),
    .B1(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__nor2_1 _10416_ (.A(_03379_),
    .B(_03381_),
    .Y(_03384_));
 sky130_fd_sc_hd__inv_2 _10417_ (.A(_03382_),
    .Y(_03385_));
 sky130_fd_sc_hd__nand2_1 _10418_ (.A(_03384_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__nand2_1 _10419_ (.A(_03383_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__a21oi_1 _10420_ (.A1(_03087_),
    .A2(_03091_),
    .B1(_03086_),
    .Y(_03389_));
 sky130_fd_sc_hd__nand2_1 _10421_ (.A(_03387_),
    .B(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__inv_2 _10422_ (.A(_03389_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand3_2 _10423_ (.A(_03383_),
    .B(_03391_),
    .C(_03386_),
    .Y(_03392_));
 sky130_fd_sc_hd__nand2_1 _10424_ (.A(_03390_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__nand2_1 _10425_ (.A(_03135_),
    .B(_03130_),
    .Y(_03394_));
 sky130_fd_sc_hd__inv_2 _10426_ (.A(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__nand2_1 _10427_ (.A(_03393_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__nand3_1 _10428_ (.A(_03390_),
    .B(_03392_),
    .C(_03394_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _10429_ (.A(_03396_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__nand2_1 _10430_ (.A(_03136_),
    .B(_03138_),
    .Y(_03400_));
 sky130_fd_sc_hd__nor2_1 _10431_ (.A(_03138_),
    .B(_03136_),
    .Y(_03401_));
 sky130_fd_sc_hd__a21oi_2 _10432_ (.A1(_03400_),
    .A2(_03124_),
    .B1(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__inv_2 _10433_ (.A(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__nand2_1 _10434_ (.A(_03398_),
    .B(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand3_1 _10435_ (.A(_03396_),
    .B(_03402_),
    .C(_03397_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _10436_ (.A(_03404_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__nand2_1 _10437_ (.A(_03157_),
    .B(_03152_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _10438_ (.A(_06245_),
    .B(_00176_),
    .Y(_03408_));
 sky130_fd_sc_hd__nand3b_1 _10439_ (.A_N(_03408_),
    .B(_06248_),
    .C(_06196_),
    .Y(_03409_));
 sky130_fd_sc_hd__inv_2 _10440_ (.A(net13),
    .Y(_03411_));
 sky130_fd_sc_hd__o21ai_1 _10441_ (.A1(_03411_),
    .A2(_06387_),
    .B1(_03408_),
    .Y(_03412_));
 sky130_fd_sc_hd__nand2_1 _10442_ (.A(_03409_),
    .B(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__nand2_1 _10443_ (.A(_06298_),
    .B(_06211_),
    .Y(_03414_));
 sky130_fd_sc_hd__nand2_1 _10444_ (.A(_03413_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand3b_1 _10445_ (.A_N(_03414_),
    .B(_03409_),
    .C(_03412_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand3_1 _10446_ (.A(_03407_),
    .B(_03415_),
    .C(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__inv_2 _10447_ (.A(_03407_),
    .Y(_03418_));
 sky130_fd_sc_hd__nand2_1 _10448_ (.A(_03415_),
    .B(_03416_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_1 _10449_ (.A(_03418_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand2_1 _10450_ (.A(_03417_),
    .B(_03420_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand2_1 _10451_ (.A(_03422_),
    .B(_06331_),
    .Y(_03423_));
 sky130_fd_sc_hd__nand3_1 _10452_ (.A(_03417_),
    .B(_03420_),
    .C(_06215_),
    .Y(_03424_));
 sky130_fd_sc_hd__nand2_1 _10453_ (.A(_03423_),
    .B(_03424_),
    .Y(_03425_));
 sky130_fd_sc_hd__inv_2 _10454_ (.A(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _10455_ (.A(_03406_),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__nand3_1 _10456_ (.A(_03404_),
    .B(_03405_),
    .C(_03425_),
    .Y(_03428_));
 sky130_fd_sc_hd__nand2_1 _10457_ (.A(_03427_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__nand2_1 _10458_ (.A(_03100_),
    .B(_03063_),
    .Y(_03430_));
 sky130_fd_sc_hd__nor2_1 _10459_ (.A(_03063_),
    .B(_03100_),
    .Y(_03431_));
 sky130_fd_sc_hd__a21oi_2 _10460_ (.A1(_03430_),
    .A2(_03104_),
    .B1(_03431_),
    .Y(_03433_));
 sky130_fd_sc_hd__inv_2 _10461_ (.A(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand2_1 _10462_ (.A(_03429_),
    .B(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__nand3_1 _10463_ (.A(_03427_),
    .B(_03428_),
    .C(_03433_),
    .Y(_03436_));
 sky130_fd_sc_hd__nand2_1 _10464_ (.A(_03435_),
    .B(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__o21a_1 _10465_ (.A1(_03123_),
    .A2(_03146_),
    .B1(_03176_),
    .X(_03438_));
 sky130_fd_sc_hd__inv_2 _10466_ (.A(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand2_1 _10467_ (.A(_03437_),
    .B(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__nand3_1 _10468_ (.A(_03438_),
    .B(_03435_),
    .C(_03436_),
    .Y(_03441_));
 sky130_fd_sc_hd__nand2_1 _10469_ (.A(_03440_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__nand3_2 _10470_ (.A(_03372_),
    .B(_03375_),
    .C(_03442_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _10471_ (.A(_03372_),
    .B(_03375_),
    .Y(_03445_));
 sky130_fd_sc_hd__inv_2 _10472_ (.A(_03442_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand2_2 _10473_ (.A(_03445_),
    .B(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand3_1 _10474_ (.A(_03239_),
    .B(_03444_),
    .C(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__nand2_1 _10475_ (.A(_03185_),
    .B(_03177_),
    .Y(_03449_));
 sky130_fd_sc_hd__nand2_1 _10476_ (.A(_03171_),
    .B(_03163_),
    .Y(_03450_));
 sky130_fd_sc_hd__nand2_1 _10477_ (.A(_03449_),
    .B(_03450_),
    .Y(_03451_));
 sky130_fd_sc_hd__inv_2 _10478_ (.A(_03450_),
    .Y(_03452_));
 sky130_fd_sc_hd__nand3_1 _10479_ (.A(_03185_),
    .B(_03177_),
    .C(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand2_1 _10480_ (.A(_03451_),
    .B(_03453_),
    .Y(_03455_));
 sky130_fd_sc_hd__nand2_1 _10481_ (.A(_03455_),
    .B(_03166_),
    .Y(_03456_));
 sky130_fd_sc_hd__nand3_1 _10482_ (.A(_03451_),
    .B(_03165_),
    .C(_03453_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_1 _10483_ (.A(_03456_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__inv_2 _10484_ (.A(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__nand2_1 _10485_ (.A(_03447_),
    .B(_03444_),
    .Y(_03460_));
 sky130_fd_sc_hd__a21oi_1 _10486_ (.A1(_03189_),
    .A2(_03236_),
    .B1(_03238_),
    .Y(_03461_));
 sky130_fd_sc_hd__nand2_1 _10487_ (.A(_03460_),
    .B(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__nand3_1 _10488_ (.A(_03448_),
    .B(_03459_),
    .C(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__nand3_1 _10489_ (.A(_03461_),
    .B(_03444_),
    .C(_03447_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_1 _10490_ (.A(_03460_),
    .B(_03239_),
    .Y(_03466_));
 sky130_fd_sc_hd__nand3_1 _10491_ (.A(_03464_),
    .B(_03466_),
    .C(_03458_),
    .Y(_03467_));
 sky130_fd_sc_hd__nand2_1 _10492_ (.A(_03463_),
    .B(_03467_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand2_1 _10493_ (.A(_03193_),
    .B(_02980_),
    .Y(_03469_));
 sky130_fd_sc_hd__nor2_1 _10494_ (.A(_02980_),
    .B(_03193_),
    .Y(_03470_));
 sky130_fd_sc_hd__a21oi_2 _10495_ (.A1(_03469_),
    .A2(_03210_),
    .B1(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__inv_2 _10496_ (.A(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand2_1 _10497_ (.A(_03468_),
    .B(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__nand3_1 _10498_ (.A(_03471_),
    .B(_03467_),
    .C(_03463_),
    .Y(_03474_));
 sky130_fd_sc_hd__nand2_1 _10499_ (.A(_03473_),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hd__nand2_1 _10500_ (.A(_03206_),
    .B(_03198_),
    .Y(_03477_));
 sky130_fd_sc_hd__inv_2 _10501_ (.A(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__nand2_1 _10502_ (.A(_03475_),
    .B(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__nand3_1 _10503_ (.A(_03473_),
    .B(_03474_),
    .C(_03477_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand3_1 _10504_ (.A(_03234_),
    .B(_03479_),
    .C(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand2_1 _10505_ (.A(_03479_),
    .B(_03480_),
    .Y(_03482_));
 sky130_fd_sc_hd__a21o_1 _10506_ (.A1(_03232_),
    .A2(_03217_),
    .B1(_03233_),
    .X(_03483_));
 sky130_fd_sc_hd__nand2_1 _10507_ (.A(_03482_),
    .B(_03483_),
    .Y(_03484_));
 sky130_fd_sc_hd__nand2_1 _10508_ (.A(_03481_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand2_1 _10509_ (.A(_03229_),
    .B(_03222_),
    .Y(_03486_));
 sky130_fd_sc_hd__xnor2_1 _10510_ (.A(_03485_),
    .B(_03486_),
    .Y(\m1.out[25] ));
 sky130_fd_sc_hd__nand2_1 _10511_ (.A(_03468_),
    .B(_03471_),
    .Y(_03487_));
 sky130_fd_sc_hd__nor2_1 _10512_ (.A(_03471_),
    .B(_03468_),
    .Y(_03488_));
 sky130_fd_sc_hd__a21o_1 _10513_ (.A1(_03487_),
    .A2(_03477_),
    .B1(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__nand2_2 _10514_ (.A(_03457_),
    .B(_03451_),
    .Y(_03490_));
 sky130_fd_sc_hd__nand2_1 _10515_ (.A(_03373_),
    .B(_03242_),
    .Y(_03491_));
 sky130_fd_sc_hd__nor2_1 _10516_ (.A(_03242_),
    .B(_03373_),
    .Y(_03492_));
 sky130_fd_sc_hd__a21oi_1 _10517_ (.A1(_03446_),
    .A2(_03491_),
    .B1(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__nand2_1 _10518_ (.A(_03317_),
    .B(_03245_),
    .Y(_03494_));
 sky130_fd_sc_hd__nor2_1 _10519_ (.A(_03245_),
    .B(_03317_),
    .Y(_03495_));
 sky130_fd_sc_hd__a21oi_2 _10520_ (.A1(_03370_),
    .A2(_03494_),
    .B1(_03495_),
    .Y(_03497_));
 sky130_fd_sc_hd__nor2_1 _10521_ (.A(_03248_),
    .B(_03285_),
    .Y(_03498_));
 sky130_fd_sc_hd__a21oi_1 _10522_ (.A1(_03313_),
    .A2(_03314_),
    .B1(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__inv_2 _10523_ (.A(_03252_),
    .Y(_03500_));
 sky130_fd_sc_hd__a21oi_1 _10524_ (.A1(_03251_),
    .A2(_03256_),
    .B1(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__nand2_1 _10525_ (.A(_06262_),
    .B(_02423_),
    .Y(_03502_));
 sky130_fd_sc_hd__nand2_1 _10526_ (.A(_03502_),
    .B(_06378_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand3_1 _10527_ (.A(_06274_),
    .B(_06262_),
    .C(_02423_),
    .Y(_03504_));
 sky130_fd_sc_hd__nand2_1 _10528_ (.A(_03503_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand2_1 _10529_ (.A(_00175_),
    .B(_02180_),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2_1 _10530_ (.A(_03505_),
    .B(_03506_),
    .Y(_03508_));
 sky130_fd_sc_hd__inv_2 _10531_ (.A(_03506_),
    .Y(_03509_));
 sky130_fd_sc_hd__nand3_1 _10532_ (.A(_03503_),
    .B(_03504_),
    .C(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__nand3_1 _10533_ (.A(_03501_),
    .B(_03508_),
    .C(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2_1 _10534_ (.A(_03508_),
    .B(_03510_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_1 _10535_ (.A(_03258_),
    .B(_03252_),
    .Y(_03513_));
 sky130_fd_sc_hd__nand2_1 _10536_ (.A(_03512_),
    .B(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2_1 _10537_ (.A(_03511_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _10538_ (.A(_06263_),
    .B(net43),
    .Y(_03516_));
 sky130_fd_sc_hd__inv_2 _10539_ (.A(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__nand2_1 _10540_ (.A(net29),
    .B(net45),
    .Y(_03519_));
 sky130_fd_sc_hd__inv_2 _10541_ (.A(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_03517_),
    .B(_03520_),
    .Y(_03521_));
 sky130_fd_sc_hd__nand2_1 _10543_ (.A(_03516_),
    .B(_03519_),
    .Y(_03522_));
 sky130_fd_sc_hd__nand2_1 _10544_ (.A(_03521_),
    .B(_03522_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _10545_ (.A(_06289_),
    .B(_06177_),
    .Y(_03524_));
 sky130_fd_sc_hd__nand2_1 _10546_ (.A(_03523_),
    .B(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__inv_2 _10547_ (.A(_03524_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand3_1 _10548_ (.A(_03521_),
    .B(_03526_),
    .C(_03522_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_2 _10549_ (.A(_03525_),
    .B(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__inv_2 _10550_ (.A(_03528_),
    .Y(_03530_));
 sky130_fd_sc_hd__nand2_1 _10551_ (.A(_03515_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__nand3_1 _10552_ (.A(_03511_),
    .B(_03514_),
    .C(_03528_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand2_2 _10553_ (.A(_03531_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__inv_2 _10554_ (.A(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__a21boi_2 _10555_ (.A1(_03281_),
    .A2(_03282_),
    .B1_N(_03280_),
    .Y(_03535_));
 sky130_fd_sc_hd__nand2_1 _10556_ (.A(_03534_),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__nor2_1 _10557_ (.A(_03263_),
    .B(_03265_),
    .Y(_03537_));
 sky130_fd_sc_hd__a21oi_1 _10558_ (.A1(_03269_),
    .A2(_03273_),
    .B1(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__inv_2 _10559_ (.A(_03538_),
    .Y(_03539_));
 sky130_fd_sc_hd__nand2_1 _10560_ (.A(_00561_),
    .B(net39),
    .Y(_03541_));
 sky130_fd_sc_hd__nand2_1 _10561_ (.A(net2),
    .B(net40),
    .Y(_03542_));
 sky130_fd_sc_hd__inv_2 _10562_ (.A(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__nand2_1 _10563_ (.A(_06286_),
    .B(net41),
    .Y(_03544_));
 sky130_fd_sc_hd__inv_2 _10564_ (.A(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__nand2_1 _10565_ (.A(_03543_),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand2_1 _10566_ (.A(_03542_),
    .B(_03544_),
    .Y(_03547_));
 sky130_fd_sc_hd__nand3b_1 _10567_ (.A_N(_03541_),
    .B(_03546_),
    .C(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__nand2_1 _10568_ (.A(_03546_),
    .B(_03547_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _10569_ (.A(_03549_),
    .B(_03541_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand3_1 _10570_ (.A(_03539_),
    .B(_03548_),
    .C(_03550_),
    .Y(_03552_));
 sky130_fd_sc_hd__nand2_1 _10571_ (.A(_03550_),
    .B(_03548_),
    .Y(_03553_));
 sky130_fd_sc_hd__nand2_1 _10572_ (.A(_03553_),
    .B(_03538_),
    .Y(_03554_));
 sky130_fd_sc_hd__nand2_1 _10573_ (.A(_03552_),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__nand2_2 _10574_ (.A(_03298_),
    .B(_03293_),
    .Y(_03556_));
 sky130_fd_sc_hd__inv_2 _10575_ (.A(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__nand2_1 _10576_ (.A(_03555_),
    .B(_03557_),
    .Y(_03558_));
 sky130_fd_sc_hd__nand3_1 _10577_ (.A(_03552_),
    .B(_03554_),
    .C(_03556_),
    .Y(_03559_));
 sky130_fd_sc_hd__nand2_2 _10578_ (.A(_03558_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__nand2_1 _10579_ (.A(_03283_),
    .B(_03280_),
    .Y(_03561_));
 sky130_fd_sc_hd__nand2_1 _10580_ (.A(_03561_),
    .B(_03533_),
    .Y(_03563_));
 sky130_fd_sc_hd__nand3_1 _10581_ (.A(_03536_),
    .B(_03560_),
    .C(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand2_1 _10582_ (.A(_03534_),
    .B(_03561_),
    .Y(_03565_));
 sky130_fd_sc_hd__inv_2 _10583_ (.A(_03560_),
    .Y(_03566_));
 sky130_fd_sc_hd__nand2_1 _10584_ (.A(_03535_),
    .B(_03533_),
    .Y(_03567_));
 sky130_fd_sc_hd__nand3_2 _10585_ (.A(_03565_),
    .B(_03566_),
    .C(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__nand3_1 _10586_ (.A(_03499_),
    .B(_03564_),
    .C(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__nand2_1 _10587_ (.A(_03568_),
    .B(_03564_),
    .Y(_03570_));
 sky130_fd_sc_hd__inv_2 _10588_ (.A(_03314_),
    .Y(_03571_));
 sky130_fd_sc_hd__o21ai_1 _10589_ (.A1(_03310_),
    .A2(_03571_),
    .B1(_03312_),
    .Y(_03572_));
 sky130_fd_sc_hd__nand2_1 _10590_ (.A(_03570_),
    .B(_03572_),
    .Y(_03574_));
 sky130_fd_sc_hd__nand2_1 _10591_ (.A(_03299_),
    .B(_03302_),
    .Y(_03575_));
 sky130_fd_sc_hd__nor2_1 _10592_ (.A(_03302_),
    .B(_03299_),
    .Y(_03576_));
 sky130_fd_sc_hd__a21oi_2 _10593_ (.A1(_03575_),
    .A2(_03307_),
    .B1(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__nand2_1 _10594_ (.A(_00701_),
    .B(_00926_),
    .Y(_03578_));
 sky130_fd_sc_hd__inv_2 _10595_ (.A(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand2_1 _10596_ (.A(_00849_),
    .B(_00921_),
    .Y(_03580_));
 sky130_fd_sc_hd__inv_2 _10597_ (.A(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__nand2_1 _10598_ (.A(_03579_),
    .B(_03581_),
    .Y(_03582_));
 sky130_fd_sc_hd__nand2_1 _10599_ (.A(_03578_),
    .B(_03580_),
    .Y(_03583_));
 sky130_fd_sc_hd__nand2_1 _10600_ (.A(_03582_),
    .B(_03583_),
    .Y(_03585_));
 sky130_fd_sc_hd__nand2_1 _10601_ (.A(_06283_),
    .B(_06219_),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(_03585_),
    .B(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__inv_2 _10603_ (.A(_03586_),
    .Y(_03588_));
 sky130_fd_sc_hd__nand3_1 _10604_ (.A(_03582_),
    .B(_03588_),
    .C(_03583_),
    .Y(_03589_));
 sky130_fd_sc_hd__nand2_1 _10605_ (.A(_03587_),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__nor2_1 _10606_ (.A(_03326_),
    .B(_03328_),
    .Y(_03591_));
 sky130_fd_sc_hd__a21oi_2 _10607_ (.A1(_03334_),
    .A2(_03332_),
    .B1(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__inv_2 _10608_ (.A(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_1 _10609_ (.A(_03590_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__nand3_1 _10610_ (.A(_03587_),
    .B(_03592_),
    .C(_03589_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_1 _10611_ (.A(_03594_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__nand2_1 _10612_ (.A(_06237_),
    .B(_06230_),
    .Y(_03598_));
 sky130_fd_sc_hd__inv_2 _10613_ (.A(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _10614_ (.A(_06281_),
    .B(_06227_),
    .Y(_03600_));
 sky130_fd_sc_hd__inv_2 _10615_ (.A(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_1 _10616_ (.A(_03599_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__nand2_1 _10617_ (.A(_03598_),
    .B(_03600_),
    .Y(_03603_));
 sky130_fd_sc_hd__nand2_1 _10618_ (.A(_06235_),
    .B(_00780_),
    .Y(_03604_));
 sky130_fd_sc_hd__inv_2 _10619_ (.A(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__a21o_1 _10620_ (.A1(_03602_),
    .A2(_03603_),
    .B1(_03605_),
    .X(_03607_));
 sky130_fd_sc_hd__nand3_1 _10621_ (.A(_03602_),
    .B(_03605_),
    .C(_03603_),
    .Y(_03608_));
 sky130_fd_sc_hd__nand2_1 _10622_ (.A(_03607_),
    .B(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__inv_2 _10623_ (.A(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand2_1 _10624_ (.A(_03597_),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand3_1 _10625_ (.A(_03594_),
    .B(_03609_),
    .C(_03596_),
    .Y(_03612_));
 sky130_fd_sc_hd__nand3_1 _10626_ (.A(_03577_),
    .B(_03611_),
    .C(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__inv_2 _10627_ (.A(_03577_),
    .Y(_03614_));
 sky130_fd_sc_hd__nand2_1 _10628_ (.A(_03611_),
    .B(_03612_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _10629_ (.A(_03614_),
    .B(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_1 _10630_ (.A(_03613_),
    .B(_03616_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _10631_ (.A(_03357_),
    .B(_03338_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand2_1 _10632_ (.A(_03618_),
    .B(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand3b_1 _10633_ (.A_N(_03619_),
    .B(_03613_),
    .C(_03616_),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2_1 _10634_ (.A(_03620_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand3_1 _10635_ (.A(_03569_),
    .B(_03574_),
    .C(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand3_1 _10636_ (.A(_03572_),
    .B(_03564_),
    .C(_03568_),
    .Y(_03624_));
 sky130_fd_sc_hd__inv_2 _10637_ (.A(_03622_),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_1 _10638_ (.A(_03570_),
    .B(_03499_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand3_1 _10639_ (.A(_03624_),
    .B(_03625_),
    .C(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand3_1 _10640_ (.A(_03497_),
    .B(_03623_),
    .C(_03627_),
    .Y(_03629_));
 sky130_fd_sc_hd__nand2_1 _10641_ (.A(_03627_),
    .B(_03623_),
    .Y(_03630_));
 sky130_fd_sc_hd__inv_2 _10642_ (.A(_03495_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_1 _10643_ (.A(_03371_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__nand2_1 _10644_ (.A(_03630_),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__inv_2 _10645_ (.A(_03392_),
    .Y(_03634_));
 sky130_fd_sc_hd__a21oi_1 _10646_ (.A1(_03390_),
    .A2(_03394_),
    .B1(_03634_),
    .Y(_03635_));
 sky130_fd_sc_hd__nand2_1 _10647_ (.A(_01858_),
    .B(_06200_),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2_1 _10648_ (.A(_06242_),
    .B(_06226_),
    .Y(_03637_));
 sky130_fd_sc_hd__nor2_1 _10649_ (.A(_03636_),
    .B(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__nand2_1 _10650_ (.A(_03636_),
    .B(_03637_),
    .Y(_03640_));
 sky130_fd_sc_hd__inv_2 _10651_ (.A(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__nand2_1 _10652_ (.A(_02095_),
    .B(_06202_),
    .Y(_03642_));
 sky130_fd_sc_hd__o21ai_1 _10653_ (.A1(_03638_),
    .A2(_03641_),
    .B1(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__nor2_1 _10654_ (.A(_03638_),
    .B(_03641_),
    .Y(_03644_));
 sky130_fd_sc_hd__inv_2 _10655_ (.A(_03642_),
    .Y(_03645_));
 sky130_fd_sc_hd__nand2_1 _10656_ (.A(_03644_),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__nand2_1 _10657_ (.A(_03643_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__nand2_2 _10658_ (.A(_03353_),
    .B(_03347_),
    .Y(_03648_));
 sky130_fd_sc_hd__inv_2 _10659_ (.A(_03648_),
    .Y(_03649_));
 sky130_fd_sc_hd__nand2_1 _10660_ (.A(_03647_),
    .B(_03649_),
    .Y(_03651_));
 sky130_fd_sc_hd__nand3_1 _10661_ (.A(_03648_),
    .B(_03643_),
    .C(_03646_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_1 _10662_ (.A(_03651_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__a21oi_1 _10663_ (.A1(_03380_),
    .A2(_03385_),
    .B1(_03379_),
    .Y(_03654_));
 sky130_fd_sc_hd__nand2_1 _10664_ (.A(_03653_),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__inv_2 _10665_ (.A(_03654_),
    .Y(_03656_));
 sky130_fd_sc_hd__nand3_1 _10666_ (.A(_03651_),
    .B(_03652_),
    .C(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand3_1 _10667_ (.A(_03635_),
    .B(_03655_),
    .C(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__nand2_1 _10668_ (.A(_03655_),
    .B(_03657_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand2_1 _10669_ (.A(_03397_),
    .B(_03392_),
    .Y(_03660_));
 sky130_fd_sc_hd__nand2_1 _10670_ (.A(_03659_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__nand2_1 _10671_ (.A(_03658_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__and2_1 _10672_ (.A(_03416_),
    .B(_03409_),
    .X(_03663_));
 sky130_fd_sc_hd__nand2_1 _10673_ (.A(net15),
    .B(_00176_),
    .Y(_03664_));
 sky130_fd_sc_hd__nor3_1 _10674_ (.A(_02871_),
    .B(_06387_),
    .C(_03664_),
    .Y(_03665_));
 sky130_fd_sc_hd__o21ai_1 _10675_ (.A1(_02871_),
    .A2(_06387_),
    .B1(_03664_),
    .Y(_03666_));
 sky130_fd_sc_hd__nor2b_1 _10676_ (.A(_03665_),
    .B_N(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__nand2_1 _10677_ (.A(_03667_),
    .B(_06212_),
    .Y(_03668_));
 sky130_fd_sc_hd__or2_1 _10678_ (.A(_06212_),
    .B(_03667_),
    .X(_03669_));
 sky130_fd_sc_hd__nand3b_2 _10679_ (.A_N(_03663_),
    .B(_03668_),
    .C(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_1 _10680_ (.A(_03669_),
    .B(_03668_),
    .Y(_03672_));
 sky130_fd_sc_hd__nand2_1 _10681_ (.A(_03672_),
    .B(_03663_),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2_1 _10682_ (.A(_03670_),
    .B(_03673_),
    .Y(_03674_));
 sky130_fd_sc_hd__inv_2 _10683_ (.A(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__nand2_1 _10684_ (.A(_03662_),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__nand3_1 _10685_ (.A(_03658_),
    .B(_03661_),
    .C(_03674_),
    .Y(_03677_));
 sky130_fd_sc_hd__nand2_1 _10686_ (.A(_03676_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__nand2_1 _10687_ (.A(_03360_),
    .B(_03321_),
    .Y(_03679_));
 sky130_fd_sc_hd__nor2_1 _10688_ (.A(_03321_),
    .B(_03360_),
    .Y(_03680_));
 sky130_fd_sc_hd__a21oi_2 _10689_ (.A1(_03679_),
    .A2(_03363_),
    .B1(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__inv_2 _10690_ (.A(_03681_),
    .Y(_03683_));
 sky130_fd_sc_hd__nand2_1 _10691_ (.A(_03678_),
    .B(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__nand3_1 _10692_ (.A(_03676_),
    .B(_03681_),
    .C(_03677_),
    .Y(_03685_));
 sky130_fd_sc_hd__nand2_1 _10693_ (.A(_03684_),
    .B(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__or2_1 _10694_ (.A(_03402_),
    .B(_03398_),
    .X(_03687_));
 sky130_fd_sc_hd__nand2_1 _10695_ (.A(_03427_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__nand2_1 _10696_ (.A(_03686_),
    .B(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand3b_1 _10697_ (.A_N(_03688_),
    .B(_03684_),
    .C(_03685_),
    .Y(_03690_));
 sky130_fd_sc_hd__nand2_1 _10698_ (.A(_03689_),
    .B(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__nand3_2 _10699_ (.A(_03629_),
    .B(_03633_),
    .C(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__nand2_1 _10700_ (.A(_03629_),
    .B(_03633_),
    .Y(_03694_));
 sky130_fd_sc_hd__inv_2 _10701_ (.A(_03691_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_1 _10702_ (.A(_03694_),
    .B(_03695_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand3_1 _10703_ (.A(_03493_),
    .B(_03692_),
    .C(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand2_1 _10704_ (.A(_03696_),
    .B(_03692_),
    .Y(_03698_));
 sky130_fd_sc_hd__a21o_1 _10705_ (.A1(_03446_),
    .A2(_03491_),
    .B1(_03492_),
    .X(_03699_));
 sky130_fd_sc_hd__nand2_1 _10706_ (.A(_03698_),
    .B(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand2_1 _10707_ (.A(_03697_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__and2_1 _10708_ (.A(_03424_),
    .B(_03417_),
    .X(_03702_));
 sky130_fd_sc_hd__o21ai_2 _10709_ (.A1(_03429_),
    .A2(_03433_),
    .B1(_03440_),
    .Y(_03703_));
 sky130_fd_sc_hd__xnor2_2 _10710_ (.A(_03702_),
    .B(_03703_),
    .Y(_03705_));
 sky130_fd_sc_hd__nand2_1 _10711_ (.A(_03701_),
    .B(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__nand3b_2 _10712_ (.A_N(_03705_),
    .B(_03697_),
    .C(_03700_),
    .Y(_03707_));
 sky130_fd_sc_hd__nand2_1 _10713_ (.A(_03706_),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__nor2_1 _10714_ (.A(_03461_),
    .B(_03460_),
    .Y(_03709_));
 sky130_fd_sc_hd__a21oi_2 _10715_ (.A1(_03462_),
    .A2(_03459_),
    .B1(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__inv_2 _10716_ (.A(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__nand2_1 _10717_ (.A(_03708_),
    .B(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand3_1 _10718_ (.A(_03710_),
    .B(_03706_),
    .C(_03707_),
    .Y(_03713_));
 sky130_fd_sc_hd__nand3b_1 _10719_ (.A_N(_03490_),
    .B(_03712_),
    .C(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__nand2_1 _10720_ (.A(_03712_),
    .B(_03713_),
    .Y(_03716_));
 sky130_fd_sc_hd__nand2_1 _10721_ (.A(_03716_),
    .B(_03490_),
    .Y(_03717_));
 sky130_fd_sc_hd__nand3_1 _10722_ (.A(_03489_),
    .B(_03714_),
    .C(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand2_1 _10723_ (.A(_03717_),
    .B(_03714_),
    .Y(_03719_));
 sky130_fd_sc_hd__a21oi_1 _10724_ (.A1(_03487_),
    .A2(_03477_),
    .B1(_03488_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand2_1 _10725_ (.A(_03719_),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__nand2_1 _10726_ (.A(_03718_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__inv_2 _10727_ (.A(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__nor2_1 _10728_ (.A(_03485_),
    .B(_03227_),
    .Y(_03724_));
 sky130_fd_sc_hd__nor2_1 _10729_ (.A(_03224_),
    .B(_03223_),
    .Y(_03725_));
 sky130_fd_sc_hd__nand3_1 _10730_ (.A(_03725_),
    .B(_03481_),
    .C(_03484_),
    .Y(_03727_));
 sky130_fd_sc_hd__nand2_1 _10731_ (.A(_03727_),
    .B(_03484_),
    .Y(_03728_));
 sky130_fd_sc_hd__a21o_1 _10732_ (.A1(_02970_),
    .A2(_03724_),
    .B1(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__or2_1 _10733_ (.A(_03723_),
    .B(_03729_),
    .X(_03730_));
 sky130_fd_sc_hd__nand2_1 _10734_ (.A(_03729_),
    .B(_03723_),
    .Y(_03731_));
 sky130_fd_sc_hd__and2_1 _10735_ (.A(_03730_),
    .B(_03731_),
    .X(_03732_));
 sky130_fd_sc_hd__clkbuf_1 _10736_ (.A(_03732_),
    .X(\m1.out[26] ));
 sky130_fd_sc_hd__nand2_1 _10737_ (.A(_03698_),
    .B(_03493_),
    .Y(_03733_));
 sky130_fd_sc_hd__nor2_1 _10738_ (.A(_03493_),
    .B(_03698_),
    .Y(_03734_));
 sky130_fd_sc_hd__a21oi_2 _10739_ (.A1(_03733_),
    .A2(_03705_),
    .B1(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand2_1 _10740_ (.A(_03630_),
    .B(_03497_),
    .Y(_03737_));
 sky130_fd_sc_hd__nor2_1 _10741_ (.A(_03497_),
    .B(_03630_),
    .Y(_03738_));
 sky130_fd_sc_hd__a21oi_1 _10742_ (.A1(_03695_),
    .A2(_03737_),
    .B1(_03738_),
    .Y(_03739_));
 sky130_fd_sc_hd__nor2_1 _10743_ (.A(_03499_),
    .B(_03570_),
    .Y(_03740_));
 sky130_fd_sc_hd__a21oi_1 _10744_ (.A1(_03625_),
    .A2(_03626_),
    .B1(_03740_),
    .Y(_03741_));
 sky130_fd_sc_hd__nor2_1 _10745_ (.A(_03533_),
    .B(_03535_),
    .Y(_03742_));
 sky130_fd_sc_hd__a21oi_1 _10746_ (.A1(_03566_),
    .A2(_03567_),
    .B1(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__nor2_1 _10747_ (.A(_06378_),
    .B(_03502_),
    .Y(_03744_));
 sky130_fd_sc_hd__a21oi_2 _10748_ (.A1(_03503_),
    .A2(_03509_),
    .B1(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__nand2_1 _10749_ (.A(_06259_),
    .B(_06183_),
    .Y(_03746_));
 sky130_fd_sc_hd__inv_2 _10750_ (.A(_06261_),
    .Y(_03748_));
 sky130_fd_sc_hd__nand2_1 _10751_ (.A(_03746_),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__nand3_2 _10752_ (.A(_06259_),
    .B(_06261_),
    .C(_06183_),
    .Y(_03750_));
 sky130_fd_sc_hd__nand2_1 _10753_ (.A(_06265_),
    .B(_02180_),
    .Y(_03751_));
 sky130_fd_sc_hd__inv_2 _10754_ (.A(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__nand3_1 _10755_ (.A(_03749_),
    .B(_03750_),
    .C(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__nand2_1 _10756_ (.A(_03749_),
    .B(_03750_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2_1 _10757_ (.A(_03754_),
    .B(_03751_),
    .Y(_03755_));
 sky130_fd_sc_hd__nand3_1 _10758_ (.A(_03745_),
    .B(_03753_),
    .C(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_1 _10759_ (.A(_03755_),
    .B(_03753_),
    .Y(_03757_));
 sky130_fd_sc_hd__nand2_1 _10760_ (.A(_03510_),
    .B(_03504_),
    .Y(_03759_));
 sky130_fd_sc_hd__nand2_1 _10761_ (.A(_03757_),
    .B(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__nand2_1 _10762_ (.A(_03756_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__nand2_1 _10763_ (.A(_06289_),
    .B(net43),
    .Y(_03762_));
 sky130_fd_sc_hd__inv_2 _10764_ (.A(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__nand2_1 _10765_ (.A(_06263_),
    .B(_06187_),
    .Y(_03764_));
 sky130_fd_sc_hd__inv_2 _10766_ (.A(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__nand2_1 _10767_ (.A(_03763_),
    .B(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__nand2_1 _10768_ (.A(_03762_),
    .B(_03764_),
    .Y(_03767_));
 sky130_fd_sc_hd__nand2_1 _10769_ (.A(_03766_),
    .B(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__nand2_1 _10770_ (.A(_06286_),
    .B(_06177_),
    .Y(_03770_));
 sky130_fd_sc_hd__nand2_1 _10771_ (.A(_03768_),
    .B(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__inv_2 _10772_ (.A(_03770_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand3_1 _10773_ (.A(_03766_),
    .B(_03772_),
    .C(_03767_),
    .Y(_03773_));
 sky130_fd_sc_hd__nand2_1 _10774_ (.A(_03771_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__inv_2 _10775_ (.A(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_1 _10776_ (.A(_03761_),
    .B(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand3_1 _10777_ (.A(_03756_),
    .B(_03760_),
    .C(_03774_),
    .Y(_03777_));
 sky130_fd_sc_hd__nand2_1 _10778_ (.A(_03776_),
    .B(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__inv_2 _10779_ (.A(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__nand2_1 _10780_ (.A(_03512_),
    .B(_03501_),
    .Y(_03781_));
 sky130_fd_sc_hd__nor2_1 _10781_ (.A(_03501_),
    .B(_03512_),
    .Y(_03782_));
 sky130_fd_sc_hd__a21oi_2 _10782_ (.A1(_03530_),
    .A2(_03781_),
    .B1(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__inv_2 _10783_ (.A(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2_1 _10784_ (.A(_03779_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__nand2_1 _10785_ (.A(_03778_),
    .B(_03783_),
    .Y(_03786_));
 sky130_fd_sc_hd__nand2_1 _10786_ (.A(_03785_),
    .B(_03786_),
    .Y(_03787_));
 sky130_fd_sc_hd__nand2_1 _10787_ (.A(net3),
    .B(net40),
    .Y(_03788_));
 sky130_fd_sc_hd__inv_2 _10788_ (.A(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__nand2_1 _10789_ (.A(net2),
    .B(net41),
    .Y(_03790_));
 sky130_fd_sc_hd__inv_2 _10790_ (.A(_03790_),
    .Y(_03792_));
 sky130_fd_sc_hd__nand2_1 _10791_ (.A(_03789_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_1 _10792_ (.A(_03788_),
    .B(_03790_),
    .Y(_03794_));
 sky130_fd_sc_hd__nand2_1 _10793_ (.A(_03793_),
    .B(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _10794_ (.A(_00849_),
    .B(net39),
    .Y(_03796_));
 sky130_fd_sc_hd__nand2_1 _10795_ (.A(_03795_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__nand3b_1 _10796_ (.A_N(_03796_),
    .B(_03793_),
    .C(_03794_),
    .Y(_03798_));
 sky130_fd_sc_hd__nand2_1 _10797_ (.A(_03797_),
    .B(_03798_),
    .Y(_03799_));
 sky130_fd_sc_hd__nor2_1 _10798_ (.A(_03516_),
    .B(_03519_),
    .Y(_03800_));
 sky130_fd_sc_hd__a21oi_2 _10799_ (.A1(_03522_),
    .A2(_03526_),
    .B1(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__inv_2 _10800_ (.A(_03801_),
    .Y(_03803_));
 sky130_fd_sc_hd__nand2_1 _10801_ (.A(_03799_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__nand3_1 _10802_ (.A(_03797_),
    .B(_03798_),
    .C(_03801_),
    .Y(_03805_));
 sky130_fd_sc_hd__nand2_1 _10803_ (.A(_03804_),
    .B(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__nand2_1 _10804_ (.A(_03548_),
    .B(_03546_),
    .Y(_03807_));
 sky130_fd_sc_hd__nand2_1 _10805_ (.A(_03806_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand3b_1 _10806_ (.A_N(_03807_),
    .B(_03804_),
    .C(_03805_),
    .Y(_03809_));
 sky130_fd_sc_hd__nand2_1 _10807_ (.A(_03808_),
    .B(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__nand2_1 _10808_ (.A(_03787_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__inv_2 _10809_ (.A(_03810_),
    .Y(_03812_));
 sky130_fd_sc_hd__nand3_1 _10810_ (.A(_03785_),
    .B(_03812_),
    .C(_03786_),
    .Y(_03814_));
 sky130_fd_sc_hd__nand3_1 _10811_ (.A(_03743_),
    .B(_03811_),
    .C(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__nand2_1 _10812_ (.A(_03811_),
    .B(_03814_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _10813_ (.A(_03568_),
    .B(_03565_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand2_1 _10814_ (.A(_03816_),
    .B(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__a21boi_2 _10815_ (.A1(_03556_),
    .A2(_03554_),
    .B1_N(_03552_),
    .Y(_03819_));
 sky130_fd_sc_hd__nor2_1 _10816_ (.A(_03578_),
    .B(_03580_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21oi_2 _10817_ (.A1(_03583_),
    .A2(_03588_),
    .B1(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__inv_2 _10818_ (.A(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__nand2_1 _10819_ (.A(_06283_),
    .B(_06217_),
    .Y(_03823_));
 sky130_fd_sc_hd__inv_2 _10820_ (.A(_03823_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2_1 _10821_ (.A(_06278_),
    .B(net38),
    .Y(_03826_));
 sky130_fd_sc_hd__inv_2 _10822_ (.A(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_1 _10823_ (.A(_03825_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__nand2_1 _10824_ (.A(_06281_),
    .B(_06219_),
    .Y(_03829_));
 sky130_fd_sc_hd__inv_2 _10825_ (.A(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_1 _10826_ (.A(_03823_),
    .B(_03826_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand3_1 _10827_ (.A(_03828_),
    .B(_03830_),
    .C(_03831_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _10828_ (.A(_03828_),
    .B(_03831_),
    .Y(_03833_));
 sky130_fd_sc_hd__nand2_1 _10829_ (.A(_03833_),
    .B(_03829_),
    .Y(_03834_));
 sky130_fd_sc_hd__nand3_1 _10830_ (.A(_03822_),
    .B(_03832_),
    .C(_03834_),
    .Y(_03836_));
 sky130_fd_sc_hd__nand2_1 _10831_ (.A(_03834_),
    .B(_03832_),
    .Y(_03837_));
 sky130_fd_sc_hd__nand2_1 _10832_ (.A(_03837_),
    .B(_03821_),
    .Y(_03838_));
 sky130_fd_sc_hd__nand2_1 _10833_ (.A(_03836_),
    .B(_03838_),
    .Y(_03839_));
 sky130_fd_sc_hd__nand2_1 _10834_ (.A(_06234_),
    .B(_06230_),
    .Y(_03840_));
 sky130_fd_sc_hd__inv_2 _10835_ (.A(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__nand2_1 _10836_ (.A(_06237_),
    .B(_00376_),
    .Y(_03842_));
 sky130_fd_sc_hd__inv_2 _10837_ (.A(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _10838_ (.A(_03841_),
    .B(_03843_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _10839_ (.A(_03840_),
    .B(_03842_),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2_1 _10840_ (.A(_03844_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_1 _10841_ (.A(_06242_),
    .B(_06225_),
    .Y(_03847_));
 sky130_fd_sc_hd__nand2_1 _10842_ (.A(_03846_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__inv_2 _10843_ (.A(_03847_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand3_1 _10844_ (.A(_03844_),
    .B(_03849_),
    .C(_03845_),
    .Y(_03850_));
 sky130_fd_sc_hd__nand2_1 _10845_ (.A(_03848_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__nand2_1 _10846_ (.A(_03839_),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__nand3b_1 _10847_ (.A_N(_03851_),
    .B(_03836_),
    .C(_03838_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand3_1 _10848_ (.A(_03819_),
    .B(_03852_),
    .C(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand2_1 _10849_ (.A(_03852_),
    .B(_03853_),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2_1 _10850_ (.A(_03559_),
    .B(_03552_),
    .Y(_03857_));
 sky130_fd_sc_hd__nand2_1 _10851_ (.A(_03855_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__nand2_1 _10852_ (.A(_03854_),
    .B(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__o21ai_2 _10853_ (.A1(_03592_),
    .A2(_03590_),
    .B1(_03611_),
    .Y(_03860_));
 sky130_fd_sc_hd__nand2_1 _10854_ (.A(_03859_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__nand3b_1 _10855_ (.A_N(_03860_),
    .B(_03854_),
    .C(_03858_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _10856_ (.A(_03861_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__nand3_1 _10857_ (.A(_03815_),
    .B(_03818_),
    .C(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__nand2_1 _10858_ (.A(_03815_),
    .B(_03818_),
    .Y(_03865_));
 sky130_fd_sc_hd__inv_2 _10859_ (.A(_03863_),
    .Y(_03866_));
 sky130_fd_sc_hd__nand2_1 _10860_ (.A(_03865_),
    .B(_03866_),
    .Y(_03868_));
 sky130_fd_sc_hd__nand3_1 _10861_ (.A(_03741_),
    .B(_03864_),
    .C(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__nand2_1 _10862_ (.A(_03868_),
    .B(_03864_),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _10863_ (.A(_03627_),
    .B(_03624_),
    .Y(_03871_));
 sky130_fd_sc_hd__nand2_1 _10864_ (.A(_03870_),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__nor2_1 _10865_ (.A(_03649_),
    .B(_03647_),
    .Y(_03873_));
 sky130_fd_sc_hd__a21oi_1 _10866_ (.A1(_03651_),
    .A2(_03656_),
    .B1(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nand2_1 _10867_ (.A(_03608_),
    .B(_03602_),
    .Y(_03875_));
 sky130_fd_sc_hd__nand2_1 _10868_ (.A(_06246_),
    .B(_06202_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _10869_ (.A(net13),
    .B(_06199_),
    .Y(_03877_));
 sky130_fd_sc_hd__inv_2 _10870_ (.A(_03877_),
    .Y(_03879_));
 sky130_fd_sc_hd__nand2_1 _10871_ (.A(_06239_),
    .B(_00270_),
    .Y(_03880_));
 sky130_fd_sc_hd__inv_2 _10872_ (.A(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__nand2_1 _10873_ (.A(_03879_),
    .B(_03881_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _10874_ (.A(_03877_),
    .B(_03880_),
    .Y(_03883_));
 sky130_fd_sc_hd__nand3b_1 _10875_ (.A_N(_03876_),
    .B(_03882_),
    .C(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hd__nand2_1 _10876_ (.A(_03882_),
    .B(_03883_),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _10877_ (.A(_03885_),
    .B(_03876_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand3_1 _10878_ (.A(_03875_),
    .B(_03884_),
    .C(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__nand2_1 _10879_ (.A(_03886_),
    .B(_03884_),
    .Y(_03888_));
 sky130_fd_sc_hd__a21boi_1 _10880_ (.A1(_03605_),
    .A2(_03603_),
    .B1_N(_03602_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _10881_ (.A(_03888_),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__nand2_1 _10882_ (.A(_03887_),
    .B(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__a21oi_1 _10883_ (.A1(_03640_),
    .A2(_03645_),
    .B1(_03638_),
    .Y(_03893_));
 sky130_fd_sc_hd__nand2_1 _10884_ (.A(_03892_),
    .B(_03893_),
    .Y(_03894_));
 sky130_fd_sc_hd__inv_2 _10885_ (.A(_03893_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand3_1 _10886_ (.A(_03887_),
    .B(_03891_),
    .C(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__nand3_1 _10887_ (.A(_03874_),
    .B(_03894_),
    .C(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_1 _10888_ (.A(_03657_),
    .B(_03652_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _10889_ (.A(_03894_),
    .B(_03896_),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _10890_ (.A(_03898_),
    .B(_03899_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _10891_ (.A(_03897_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__and3_1 _10892_ (.A(net15),
    .B(_06196_),
    .C(_00176_),
    .X(_03903_));
 sky130_fd_sc_hd__inv_2 _10893_ (.A(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__clkbuf_4 _10894_ (.A(_06298_),
    .X(_03905_));
 sky130_fd_sc_hd__a21o_1 _10895_ (.A1(_03905_),
    .A2(_06196_),
    .B1(_06198_),
    .X(_03906_));
 sky130_fd_sc_hd__nand2_1 _10896_ (.A(_03904_),
    .B(_03906_),
    .Y(_03907_));
 sky130_fd_sc_hd__a21oi_1 _10897_ (.A1(_03666_),
    .A2(_06212_),
    .B1(_03665_),
    .Y(_03908_));
 sky130_fd_sc_hd__nor2_1 _10898_ (.A(_03907_),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__inv_2 _10899_ (.A(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _10900_ (.A(_03908_),
    .B(_03907_),
    .Y(_03912_));
 sky130_fd_sc_hd__and2_1 _10901_ (.A(_03910_),
    .B(_03912_),
    .X(_03913_));
 sky130_fd_sc_hd__nand2_1 _10902_ (.A(_03902_),
    .B(_03913_),
    .Y(_03914_));
 sky130_fd_sc_hd__nand3b_1 _10903_ (.A_N(_03913_),
    .B(_03897_),
    .C(_03901_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand2_1 _10904_ (.A(_03914_),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2_1 _10905_ (.A(_03615_),
    .B(_03577_),
    .Y(_03917_));
 sky130_fd_sc_hd__nor2_1 _10906_ (.A(_03577_),
    .B(_03615_),
    .Y(_03918_));
 sky130_fd_sc_hd__a21oi_2 _10907_ (.A1(_03917_),
    .A2(_03619_),
    .B1(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__inv_2 _10908_ (.A(_03919_),
    .Y(_03920_));
 sky130_fd_sc_hd__nand2_1 _10909_ (.A(_03916_),
    .B(_03920_),
    .Y(_03921_));
 sky130_fd_sc_hd__nand3_1 _10910_ (.A(_03914_),
    .B(_03915_),
    .C(_03919_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand2_1 _10911_ (.A(_03921_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__or2_1 _10912_ (.A(_03635_),
    .B(_03659_),
    .X(_03925_));
 sky130_fd_sc_hd__nand2_1 _10913_ (.A(_03676_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__nand2_1 _10914_ (.A(_03924_),
    .B(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand3b_1 _10915_ (.A_N(_03926_),
    .B(_03921_),
    .C(_03923_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand2_1 _10916_ (.A(_03927_),
    .B(_03928_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand3_1 _10917_ (.A(_03869_),
    .B(_03872_),
    .C(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__nand2_1 _10918_ (.A(_03869_),
    .B(_03872_),
    .Y(_03931_));
 sky130_fd_sc_hd__inv_2 _10919_ (.A(_03929_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _10920_ (.A(_03931_),
    .B(_03932_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand3_1 _10921_ (.A(_03739_),
    .B(_03930_),
    .C(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__nand2_1 _10922_ (.A(_03934_),
    .B(_03930_),
    .Y(_03936_));
 sky130_fd_sc_hd__inv_2 _10923_ (.A(_03737_),
    .Y(_03937_));
 sky130_fd_sc_hd__o21bai_1 _10924_ (.A1(_03691_),
    .A2(_03937_),
    .B1_N(_03738_),
    .Y(_03938_));
 sky130_fd_sc_hd__nand2_1 _10925_ (.A(_03936_),
    .B(_03938_),
    .Y(_03939_));
 sky130_fd_sc_hd__or2_1 _10926_ (.A(_03681_),
    .B(_03678_),
    .X(_03940_));
 sky130_fd_sc_hd__and2_1 _10927_ (.A(_03689_),
    .B(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__nor2_2 _10928_ (.A(_03670_),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__inv_2 _10929_ (.A(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _10930_ (.A(_03941_),
    .B(_03670_),
    .Y(_03945_));
 sky130_fd_sc_hd__nand2_1 _10931_ (.A(_03943_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__nand3_2 _10932_ (.A(_03935_),
    .B(_03939_),
    .C(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand3_1 _10933_ (.A(_03938_),
    .B(_03930_),
    .C(_03934_),
    .Y(_03948_));
 sky130_fd_sc_hd__nor2b_1 _10934_ (.A(_03942_),
    .B_N(_03945_),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_1 _10935_ (.A(_03936_),
    .B(_03739_),
    .Y(_03950_));
 sky130_fd_sc_hd__nand3_2 _10936_ (.A(_03948_),
    .B(_03949_),
    .C(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__nand3_2 _10937_ (.A(_03735_),
    .B(_03947_),
    .C(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__nand2_1 _10938_ (.A(_03951_),
    .B(_03947_),
    .Y(_03953_));
 sky130_fd_sc_hd__a21o_1 _10939_ (.A1(_03733_),
    .A2(_03705_),
    .B1(_03734_),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_2 _10940_ (.A(_03953_),
    .B(_03954_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand2_1 _10941_ (.A(_03952_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__inv_2 _10942_ (.A(_03703_),
    .Y(_03958_));
 sky130_fd_sc_hd__nor2_2 _10943_ (.A(_03702_),
    .B(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__inv_2 _10944_ (.A(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_1 _10945_ (.A(_03957_),
    .B(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand3_1 _10946_ (.A(_03952_),
    .B(_03956_),
    .C(_03959_),
    .Y(_03962_));
 sky130_fd_sc_hd__nand2_1 _10947_ (.A(_03961_),
    .B(_03962_),
    .Y(_03963_));
 sky130_fd_sc_hd__nand2_1 _10948_ (.A(_03708_),
    .B(_03710_),
    .Y(_03964_));
 sky130_fd_sc_hd__nor2_1 _10949_ (.A(_03710_),
    .B(_03708_),
    .Y(_03965_));
 sky130_fd_sc_hd__a21o_1 _10950_ (.A1(_03964_),
    .A2(_03490_),
    .B1(_03965_),
    .X(_03967_));
 sky130_fd_sc_hd__nand2_1 _10951_ (.A(_03963_),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__nand2_1 _10952_ (.A(_03957_),
    .B(_03959_),
    .Y(_03969_));
 sky130_fd_sc_hd__nand3_1 _10953_ (.A(_03952_),
    .B(_03956_),
    .C(_03960_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _10954_ (.A(_03969_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__a21oi_1 _10955_ (.A1(_03964_),
    .A2(_03490_),
    .B1(_03965_),
    .Y(_03972_));
 sky130_fd_sc_hd__nand2_1 _10956_ (.A(_03971_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand2_1 _10957_ (.A(_03968_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _10958_ (.A(_03731_),
    .B(_03718_),
    .Y(_03975_));
 sky130_fd_sc_hd__xnor2_1 _10959_ (.A(_03974_),
    .B(_03975_),
    .Y(\m1.out[27] ));
 sky130_fd_sc_hd__nand2_1 _10960_ (.A(_03953_),
    .B(_03735_),
    .Y(_03977_));
 sky130_fd_sc_hd__nor2_1 _10961_ (.A(_03735_),
    .B(_03953_),
    .Y(_03978_));
 sky130_fd_sc_hd__a21oi_2 _10962_ (.A1(_03977_),
    .A2(_03959_),
    .B1(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_1 _10963_ (.A(_03870_),
    .B(_03741_),
    .Y(_03980_));
 sky130_fd_sc_hd__inv_2 _10964_ (.A(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__nor2_1 _10965_ (.A(_03741_),
    .B(_03870_),
    .Y(_03982_));
 sky130_fd_sc_hd__o21bai_1 _10966_ (.A1(_03929_),
    .A2(_03981_),
    .B1_N(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _10967_ (.A(_03816_),
    .B(_03743_),
    .Y(_03984_));
 sky130_fd_sc_hd__nor2_1 _10968_ (.A(_03743_),
    .B(_03816_),
    .Y(_03985_));
 sky130_fd_sc_hd__a21oi_1 _10969_ (.A1(_03866_),
    .A2(_03984_),
    .B1(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__nand2_1 _10970_ (.A(_03757_),
    .B(_03745_),
    .Y(_03988_));
 sky130_fd_sc_hd__nor2_1 _10971_ (.A(_03745_),
    .B(_03757_),
    .Y(_03989_));
 sky130_fd_sc_hd__a21o_1 _10972_ (.A1(_03775_),
    .A2(_03988_),
    .B1(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__nand2_1 _10973_ (.A(_03753_),
    .B(_03750_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _10974_ (.A(_06264_),
    .B(_02180_),
    .Y(_03992_));
 sky130_fd_sc_hd__nand2_1 _10975_ (.A(_06266_),
    .B(_06183_),
    .Y(_03993_));
 sky130_fd_sc_hd__inv_2 _10976_ (.A(_06258_),
    .Y(_03994_));
 sky130_fd_sc_hd__nand2_1 _10977_ (.A(_03993_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand3_2 _10978_ (.A(_00175_),
    .B(_06266_),
    .C(_06183_),
    .Y(_03996_));
 sky130_fd_sc_hd__nand3b_2 _10979_ (.A_N(_03992_),
    .B(_03995_),
    .C(_03996_),
    .Y(_03997_));
 sky130_fd_sc_hd__nand2_1 _10980_ (.A(_03995_),
    .B(_03996_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_1 _10981_ (.A(_03999_),
    .B(_03992_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand3_2 _10982_ (.A(_03991_),
    .B(_03997_),
    .C(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__nand2_1 _10983_ (.A(_04000_),
    .B(_03997_),
    .Y(_04002_));
 sky130_fd_sc_hd__a21boi_1 _10984_ (.A1(_03749_),
    .A2(_03752_),
    .B1_N(_03750_),
    .Y(_04003_));
 sky130_fd_sc_hd__nand2_1 _10985_ (.A(_04002_),
    .B(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2_1 _10986_ (.A(_04001_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__nand2_1 _10987_ (.A(_06286_),
    .B(_06175_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_1 _10988_ (.A(_06289_),
    .B(_06187_),
    .Y(_04007_));
 sky130_fd_sc_hd__nor2_1 _10989_ (.A(_04006_),
    .B(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__inv_2 _10990_ (.A(_04008_),
    .Y(_04010_));
 sky130_fd_sc_hd__nand2_1 _10991_ (.A(_04006_),
    .B(_04007_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand2_1 _10992_ (.A(_04010_),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__nand2_1 _10993_ (.A(_00439_),
    .B(_06177_),
    .Y(_04013_));
 sky130_fd_sc_hd__nand2_1 _10994_ (.A(_04012_),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__inv_2 _10995_ (.A(_04013_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand3_1 _10996_ (.A(_04010_),
    .B(_04015_),
    .C(_04011_),
    .Y(_04016_));
 sky130_fd_sc_hd__nand2_2 _10997_ (.A(_04014_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__nand2_1 _10998_ (.A(_04005_),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__inv_2 _10999_ (.A(_04017_),
    .Y(_04019_));
 sky130_fd_sc_hd__nand3_1 _11000_ (.A(_04019_),
    .B(_04001_),
    .C(_04004_),
    .Y(_04020_));
 sky130_fd_sc_hd__nand3_1 _11001_ (.A(_03990_),
    .B(_04018_),
    .C(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__nand2_1 _11002_ (.A(_04020_),
    .B(_04018_),
    .Y(_04022_));
 sky130_fd_sc_hd__a21oi_1 _11003_ (.A1(_03775_),
    .A2(_03988_),
    .B1(_03989_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2_1 _11004_ (.A(_04022_),
    .B(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hd__nand2_1 _11005_ (.A(net4),
    .B(_06173_),
    .Y(_04025_));
 sky130_fd_sc_hd__inv_2 _11006_ (.A(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__nand2_1 _11007_ (.A(_00561_),
    .B(_01280_),
    .Y(_04027_));
 sky130_fd_sc_hd__inv_2 _11008_ (.A(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__nand2_1 _11009_ (.A(_04026_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _11010_ (.A(_04025_),
    .B(_04027_),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_1 _11011_ (.A(_04029_),
    .B(_04031_),
    .Y(_04032_));
 sky130_fd_sc_hd__nand2_1 _11012_ (.A(_06279_),
    .B(_00918_),
    .Y(_04033_));
 sky130_fd_sc_hd__nand2_1 _11013_ (.A(_04032_),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__nand3b_1 _11014_ (.A_N(_04033_),
    .B(_04029_),
    .C(_04031_),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_1 _11015_ (.A(_04034_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__nor2_1 _11016_ (.A(_03762_),
    .B(_03764_),
    .Y(_04037_));
 sky130_fd_sc_hd__a21oi_2 _11017_ (.A1(_03767_),
    .A2(_03772_),
    .B1(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__inv_2 _11018_ (.A(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__nand2_1 _11019_ (.A(_04036_),
    .B(_04039_),
    .Y(_04040_));
 sky130_fd_sc_hd__nand3_1 _11020_ (.A(_04034_),
    .B(_04035_),
    .C(_04038_),
    .Y(_04042_));
 sky130_fd_sc_hd__nand2_1 _11021_ (.A(_04040_),
    .B(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__nand2_1 _11022_ (.A(_03798_),
    .B(_03793_),
    .Y(_04044_));
 sky130_fd_sc_hd__nand2_1 _11023_ (.A(_04043_),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand3b_1 _11024_ (.A_N(_04044_),
    .B(_04040_),
    .C(_04042_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_1 _11025_ (.A(_04045_),
    .B(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__inv_2 _11026_ (.A(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hd__nand3_1 _11027_ (.A(_04021_),
    .B(_04024_),
    .C(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__nand2_1 _11028_ (.A(_04022_),
    .B(_03990_),
    .Y(_04050_));
 sky130_fd_sc_hd__nand3_1 _11029_ (.A(_04023_),
    .B(_04018_),
    .C(_04020_),
    .Y(_04051_));
 sky130_fd_sc_hd__nand3_1 _11030_ (.A(_04050_),
    .B(_04051_),
    .C(_04047_),
    .Y(_04053_));
 sky130_fd_sc_hd__nand2_1 _11031_ (.A(_04049_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__nor2_1 _11032_ (.A(_03783_),
    .B(_03778_),
    .Y(_04055_));
 sky130_fd_sc_hd__a21oi_2 _11033_ (.A1(_03812_),
    .A2(_03786_),
    .B1(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hd__inv_2 _11034_ (.A(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__nand2_1 _11035_ (.A(_04054_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__nand3_1 _11036_ (.A(_04056_),
    .B(_04049_),
    .C(_04053_),
    .Y(_04059_));
 sky130_fd_sc_hd__nand2_1 _11037_ (.A(_03832_),
    .B(_03828_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _11038_ (.A(_01831_),
    .B(_00926_),
    .Y(_04061_));
 sky130_fd_sc_hd__inv_2 _11039_ (.A(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__nand2_1 _11040_ (.A(_01158_),
    .B(_00921_),
    .Y(_04064_));
 sky130_fd_sc_hd__inv_2 _11041_ (.A(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand2_1 _11042_ (.A(_04062_),
    .B(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__nand2_1 _11043_ (.A(_01211_),
    .B(_06220_),
    .Y(_04067_));
 sky130_fd_sc_hd__inv_2 _11044_ (.A(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__nand2_1 _11045_ (.A(_04061_),
    .B(_04064_),
    .Y(_04069_));
 sky130_fd_sc_hd__nand3_1 _11046_ (.A(_04066_),
    .B(_04068_),
    .C(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_1 _11047_ (.A(_04066_),
    .B(_04069_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_1 _11048_ (.A(_04071_),
    .B(_04067_),
    .Y(_04072_));
 sky130_fd_sc_hd__nand3_1 _11049_ (.A(_04060_),
    .B(_04070_),
    .C(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__inv_2 _11050_ (.A(_04060_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_1 _11051_ (.A(_04072_),
    .B(_04070_),
    .Y(_04076_));
 sky130_fd_sc_hd__nand2_1 _11052_ (.A(_04075_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__nand2_1 _11053_ (.A(_04073_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__nand2_1 _11054_ (.A(_06241_),
    .B(_06230_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2_1 _11055_ (.A(_06234_),
    .B(_00376_),
    .Y(_04080_));
 sky130_fd_sc_hd__or2_1 _11056_ (.A(_04079_),
    .B(_04080_),
    .X(_04081_));
 sky130_fd_sc_hd__nand2_1 _11057_ (.A(_04079_),
    .B(_04080_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _11058_ (.A(_04081_),
    .B(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__nand2_1 _11059_ (.A(_06239_),
    .B(_00780_),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _11060_ (.A(_04083_),
    .B(_04084_),
    .Y(_04086_));
 sky130_fd_sc_hd__inv_2 _11061_ (.A(_04084_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand3_1 _11062_ (.A(_04081_),
    .B(_04082_),
    .C(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand2_1 _11063_ (.A(_04086_),
    .B(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__nand2_1 _11064_ (.A(_04078_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__inv_2 _11065_ (.A(_04089_),
    .Y(_04091_));
 sky130_fd_sc_hd__nand3_1 _11066_ (.A(_04091_),
    .B(_04073_),
    .C(_04077_),
    .Y(_04092_));
 sky130_fd_sc_hd__nand2_1 _11067_ (.A(_04090_),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__nand2_1 _11068_ (.A(_03799_),
    .B(_03801_),
    .Y(_04094_));
 sky130_fd_sc_hd__nor2_1 _11069_ (.A(_03801_),
    .B(_03799_),
    .Y(_04095_));
 sky130_fd_sc_hd__a21oi_2 _11070_ (.A1(_04094_),
    .A2(_03807_),
    .B1(_04095_),
    .Y(_04097_));
 sky130_fd_sc_hd__inv_2 _11071_ (.A(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__nand2_1 _11072_ (.A(_04093_),
    .B(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__nand3_1 _11073_ (.A(_04097_),
    .B(_04090_),
    .C(_04092_),
    .Y(_04100_));
 sky130_fd_sc_hd__nand2_1 _11074_ (.A(_04099_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_1 _11075_ (.A(_03853_),
    .B(_03836_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand2_1 _11076_ (.A(_04101_),
    .B(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__nand3b_1 _11077_ (.A_N(_04102_),
    .B(_04099_),
    .C(_04100_),
    .Y(_04104_));
 sky130_fd_sc_hd__nand2_1 _11078_ (.A(_04103_),
    .B(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hd__nand3_1 _11079_ (.A(_04058_),
    .B(_04059_),
    .C(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__nand2_1 _11080_ (.A(_04058_),
    .B(_04059_),
    .Y(_04108_));
 sky130_fd_sc_hd__inv_2 _11081_ (.A(_04105_),
    .Y(_04109_));
 sky130_fd_sc_hd__nand2_1 _11082_ (.A(_04108_),
    .B(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__nand3_1 _11083_ (.A(_03986_),
    .B(_04106_),
    .C(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__a21o_1 _11084_ (.A1(_03866_),
    .A2(_03984_),
    .B1(_03985_),
    .X(_04112_));
 sky130_fd_sc_hd__nand2_1 _11085_ (.A(_04110_),
    .B(_04106_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand2_1 _11086_ (.A(_04112_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand2_1 _11087_ (.A(_03850_),
    .B(_03844_),
    .Y(_04115_));
 sky130_fd_sc_hd__nand2_1 _11088_ (.A(_06298_),
    .B(_06202_),
    .Y(_04116_));
 sky130_fd_sc_hd__nand2_1 _11089_ (.A(_06245_),
    .B(_06199_),
    .Y(_04117_));
 sky130_fd_sc_hd__inv_2 _11090_ (.A(_04117_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _11091_ (.A(net13),
    .B(_00270_),
    .Y(_04120_));
 sky130_fd_sc_hd__inv_2 _11092_ (.A(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _11093_ (.A(_04119_),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand2_1 _11094_ (.A(_04117_),
    .B(_04120_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand3b_1 _11095_ (.A_N(_04116_),
    .B(_04122_),
    .C(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_1 _11096_ (.A(_04122_),
    .B(_04123_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _11097_ (.A(_04125_),
    .B(_04116_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand3_1 _11098_ (.A(_04115_),
    .B(_04124_),
    .C(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__nand2_1 _11099_ (.A(_04126_),
    .B(_04124_),
    .Y(_04128_));
 sky130_fd_sc_hd__a21boi_1 _11100_ (.A1(_03849_),
    .A2(_03845_),
    .B1_N(_03844_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _11101_ (.A(_04128_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__nand2_1 _11102_ (.A(_04127_),
    .B(_04131_),
    .Y(_04132_));
 sky130_fd_sc_hd__nand2_1 _11103_ (.A(_03884_),
    .B(_03882_),
    .Y(_04133_));
 sky130_fd_sc_hd__inv_2 _11104_ (.A(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2_1 _11105_ (.A(_04132_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__nand3_1 _11106_ (.A(_04127_),
    .B(_04131_),
    .C(_04133_),
    .Y(_04136_));
 sky130_fd_sc_hd__nand2_1 _11107_ (.A(_04135_),
    .B(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hd__nor2_1 _11108_ (.A(_03890_),
    .B(_03888_),
    .Y(_04138_));
 sky130_fd_sc_hd__a21oi_2 _11109_ (.A1(_03891_),
    .A2(_03895_),
    .B1(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__inv_2 _11110_ (.A(_04139_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_1 _11111_ (.A(_04137_),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand3_1 _11112_ (.A(_04139_),
    .B(_04135_),
    .C(_04136_),
    .Y(_04143_));
 sky130_fd_sc_hd__nand2_1 _11113_ (.A(_04142_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__nor2_1 _11114_ (.A(_06387_),
    .B(_03903_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2_1 _11115_ (.A(_04144_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand3b_1 _11116_ (.A_N(_04145_),
    .B(_04142_),
    .C(_04143_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand2_1 _11117_ (.A(_04146_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__nand2_1 _11118_ (.A(_03855_),
    .B(_03819_),
    .Y(_04149_));
 sky130_fd_sc_hd__nor2_1 _11119_ (.A(_03819_),
    .B(_03855_),
    .Y(_04150_));
 sky130_fd_sc_hd__a21oi_4 _11120_ (.A1(_04149_),
    .A2(_03860_),
    .B1(_04150_),
    .Y(_04152_));
 sky130_fd_sc_hd__inv_2 _11121_ (.A(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__nand2_1 _11122_ (.A(_04148_),
    .B(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__nand3_1 _11123_ (.A(_04152_),
    .B(_04146_),
    .C(_04147_),
    .Y(_04155_));
 sky130_fd_sc_hd__nand2_1 _11124_ (.A(_04154_),
    .B(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__or2_1 _11125_ (.A(_03874_),
    .B(_03899_),
    .X(_04157_));
 sky130_fd_sc_hd__nand2_1 _11126_ (.A(_03914_),
    .B(_04157_),
    .Y(_04158_));
 sky130_fd_sc_hd__nand2_1 _11127_ (.A(_04156_),
    .B(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__nand3b_1 _11128_ (.A_N(_04158_),
    .B(_04154_),
    .C(_04155_),
    .Y(_04160_));
 sky130_fd_sc_hd__nand2_1 _11129_ (.A(_04159_),
    .B(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__nand3_2 _11130_ (.A(_04111_),
    .B(_04114_),
    .C(_04161_),
    .Y(_04163_));
 sky130_fd_sc_hd__inv_2 _11131_ (.A(_04113_),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2_1 _11132_ (.A(_04164_),
    .B(_04112_),
    .Y(_04165_));
 sky130_fd_sc_hd__inv_2 _11133_ (.A(_04161_),
    .Y(_04166_));
 sky130_fd_sc_hd__nand2_1 _11134_ (.A(_04113_),
    .B(_03986_),
    .Y(_04167_));
 sky130_fd_sc_hd__nand3_2 _11135_ (.A(_04165_),
    .B(_04166_),
    .C(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__nand3_1 _11136_ (.A(_03983_),
    .B(_04163_),
    .C(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__o21a_1 _11137_ (.A1(_03916_),
    .A2(_03919_),
    .B1(_03927_),
    .X(_04170_));
 sky130_fd_sc_hd__xor2_1 _11138_ (.A(_03910_),
    .B(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__nand2_1 _11139_ (.A(_04168_),
    .B(_04163_),
    .Y(_04172_));
 sky130_fd_sc_hd__a21oi_2 _11140_ (.A1(_03932_),
    .A2(_03980_),
    .B1(_03982_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand2_1 _11141_ (.A(_04172_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nand3_1 _11142_ (.A(_04169_),
    .B(_04171_),
    .C(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__nand3_1 _11143_ (.A(_04174_),
    .B(_04163_),
    .C(_04168_),
    .Y(_04177_));
 sky130_fd_sc_hd__nand2_1 _11144_ (.A(_04172_),
    .B(_03983_),
    .Y(_04178_));
 sky130_fd_sc_hd__nor2_1 _11145_ (.A(_03910_),
    .B(_04170_),
    .Y(_04179_));
 sky130_fd_sc_hd__inv_2 _11146_ (.A(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__nand2_1 _11147_ (.A(_04170_),
    .B(_03910_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand2_1 _11148_ (.A(_04180_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__nand3_1 _11149_ (.A(_04177_),
    .B(_04178_),
    .C(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_1 _11150_ (.A(_04176_),
    .B(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__nor2_1 _11151_ (.A(_03739_),
    .B(_03936_),
    .Y(_04185_));
 sky130_fd_sc_hd__a21oi_2 _11152_ (.A1(_03950_),
    .A2(_03949_),
    .B1(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__inv_2 _11153_ (.A(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand2_1 _11154_ (.A(_04184_),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand3_1 _11155_ (.A(_04186_),
    .B(_04176_),
    .C(_04183_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand2_1 _11156_ (.A(_04188_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__nand2_1 _11157_ (.A(_04190_),
    .B(_03942_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand3_1 _11158_ (.A(_04188_),
    .B(_04189_),
    .C(_03943_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand2_1 _11159_ (.A(_04191_),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__nor2_1 _11160_ (.A(_03979_),
    .B(_04193_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _11161_ (.A(_04193_),
    .B(_03979_),
    .Y(_04196_));
 sky130_fd_sc_hd__inv_2 _11162_ (.A(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hd__nor2_1 _11163_ (.A(_04195_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__nor2_1 _11164_ (.A(_03974_),
    .B(_03722_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_2 _11165_ (.A(_03724_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _11166_ (.A(_03728_),
    .B(_04199_),
    .Y(_04201_));
 sky130_fd_sc_hd__nor2_1 _11167_ (.A(_03967_),
    .B(_03963_),
    .Y(_04202_));
 sky130_fd_sc_hd__o21a_1 _11168_ (.A1(_03718_),
    .A2(_04202_),
    .B1(_03968_),
    .X(_04203_));
 sky130_fd_sc_hd__nand2_2 _11169_ (.A(_04201_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o21bai_2 _11170_ (.A1(_04200_),
    .A2(_02969_),
    .B1_N(_04204_),
    .Y(_04206_));
 sky130_fd_sc_hd__or2_1 _11171_ (.A(_04198_),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__nand2_1 _11172_ (.A(_04206_),
    .B(_04198_),
    .Y(_04208_));
 sky130_fd_sc_hd__and2_1 _11173_ (.A(_04207_),
    .B(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__buf_1 _11174_ (.A(_04209_),
    .X(\m1.out[28] ));
 sky130_fd_sc_hd__nor2_1 _11175_ (.A(_03986_),
    .B(_04113_),
    .Y(_04210_));
 sky130_fd_sc_hd__a21oi_1 _11176_ (.A1(_04166_),
    .A2(_04167_),
    .B1(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__nand2_1 _11177_ (.A(_04054_),
    .B(_04056_),
    .Y(_04212_));
 sky130_fd_sc_hd__nor2_1 _11178_ (.A(_04056_),
    .B(_04054_),
    .Y(_04213_));
 sky130_fd_sc_hd__a21oi_1 _11179_ (.A1(_04109_),
    .A2(_04212_),
    .B1(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__inv_2 _11180_ (.A(_04004_),
    .Y(_04216_));
 sky130_fd_sc_hd__o21ai_2 _11181_ (.A1(_04017_),
    .A2(_04216_),
    .B1(_04001_),
    .Y(_04217_));
 sky130_fd_sc_hd__inv_2 _11182_ (.A(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__nand2_1 _11183_ (.A(_06264_),
    .B(_02423_),
    .Y(_04219_));
 sky130_fd_sc_hd__nand2_1 _11184_ (.A(_04219_),
    .B(_00069_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand3_2 _11185_ (.A(_06264_),
    .B(_06266_),
    .C(_06184_),
    .Y(_04221_));
 sky130_fd_sc_hd__nand2_1 _11186_ (.A(_04220_),
    .B(_04221_),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_1 _11187_ (.A(_06290_),
    .B(_02181_),
    .Y(_04223_));
 sky130_fd_sc_hd__nand2_1 _11188_ (.A(_04222_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hd__nand3b_2 _11189_ (.A_N(_04223_),
    .B(_04220_),
    .C(_04221_),
    .Y(_04225_));
 sky130_fd_sc_hd__nand2_1 _11190_ (.A(_04224_),
    .B(_04225_),
    .Y(_04227_));
 sky130_fd_sc_hd__nand3_1 _11191_ (.A(_04227_),
    .B(_03996_),
    .C(_03997_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand2_1 _11192_ (.A(_03997_),
    .B(_03996_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand3_2 _11193_ (.A(_04229_),
    .B(_04224_),
    .C(_04225_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_1 _11194_ (.A(_04228_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__nand2_1 _11195_ (.A(_00439_),
    .B(_06175_),
    .Y(_04232_));
 sky130_fd_sc_hd__inv_2 _11196_ (.A(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__nand2_1 _11197_ (.A(_06286_),
    .B(_06187_),
    .Y(_04234_));
 sky130_fd_sc_hd__inv_2 _11198_ (.A(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hd__nand2_1 _11199_ (.A(_04233_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__nand2_1 _11200_ (.A(_04232_),
    .B(_04234_),
    .Y(_04238_));
 sky130_fd_sc_hd__nand2_1 _11201_ (.A(_04236_),
    .B(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_1 _11202_ (.A(_00561_),
    .B(_06177_),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2_1 _11203_ (.A(_04239_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__inv_2 _11204_ (.A(_04240_),
    .Y(_04242_));
 sky130_fd_sc_hd__nand3_1 _11205_ (.A(_04236_),
    .B(_04242_),
    .C(_04238_),
    .Y(_04243_));
 sky130_fd_sc_hd__nand2_1 _11206_ (.A(_04241_),
    .B(_04243_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_1 _11207_ (.A(_04231_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__inv_2 _11208_ (.A(_04244_),
    .Y(_04246_));
 sky130_fd_sc_hd__nand3_2 _11209_ (.A(_04228_),
    .B(_04230_),
    .C(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__nand2_1 _11210_ (.A(_04245_),
    .B(_04247_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_1 _11211_ (.A(_04218_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__nand3_2 _11212_ (.A(_04217_),
    .B(_04245_),
    .C(_04247_),
    .Y(_04251_));
 sky130_fd_sc_hd__nand2_1 _11213_ (.A(_04250_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _11214_ (.A(_06278_),
    .B(_06173_),
    .Y(_04253_));
 sky130_fd_sc_hd__nand2_1 _11215_ (.A(_00849_),
    .B(_01280_),
    .Y(_04254_));
 sky130_fd_sc_hd__or2_1 _11216_ (.A(_04253_),
    .B(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__nand2_1 _11217_ (.A(_04253_),
    .B(_04254_),
    .Y(_04256_));
 sky130_fd_sc_hd__nand2_1 _11218_ (.A(_04255_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__nand2_1 _11219_ (.A(_01158_),
    .B(net39),
    .Y(_04258_));
 sky130_fd_sc_hd__nand2_1 _11220_ (.A(_04257_),
    .B(_04258_),
    .Y(_04260_));
 sky130_fd_sc_hd__inv_2 _11221_ (.A(_04258_),
    .Y(_04261_));
 sky130_fd_sc_hd__nand3_2 _11222_ (.A(_04255_),
    .B(_04261_),
    .C(_04256_),
    .Y(_04262_));
 sky130_fd_sc_hd__nand2_1 _11223_ (.A(_04260_),
    .B(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__a21oi_2 _11224_ (.A1(_04011_),
    .A2(_04015_),
    .B1(_04008_),
    .Y(_04264_));
 sky130_fd_sc_hd__inv_2 _11225_ (.A(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_1 _11226_ (.A(_04263_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__nand3_1 _11227_ (.A(_04260_),
    .B(_04262_),
    .C(_04264_),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _11228_ (.A(_04266_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_1 _11229_ (.A(_04035_),
    .B(_04029_),
    .Y(_04269_));
 sky130_fd_sc_hd__nand2_1 _11230_ (.A(_04268_),
    .B(_04269_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand3b_1 _11231_ (.A_N(_04269_),
    .B(_04266_),
    .C(_04267_),
    .Y(_04272_));
 sky130_fd_sc_hd__nand2_1 _11232_ (.A(_04271_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__nand2_1 _11233_ (.A(_04252_),
    .B(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__inv_2 _11234_ (.A(_04273_),
    .Y(_04275_));
 sky130_fd_sc_hd__nand3_2 _11235_ (.A(_04275_),
    .B(_04250_),
    .C(_04251_),
    .Y(_04276_));
 sky130_fd_sc_hd__nand2_1 _11236_ (.A(_04274_),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(_04049_),
    .B(_04021_),
    .Y(_04278_));
 sky130_fd_sc_hd__nand2_1 _11238_ (.A(_04277_),
    .B(_04278_),
    .Y(_04279_));
 sky130_fd_sc_hd__nor2_1 _11239_ (.A(_04023_),
    .B(_04022_),
    .Y(_04280_));
 sky130_fd_sc_hd__a21oi_1 _11240_ (.A1(_04048_),
    .A2(_04024_),
    .B1(_04280_),
    .Y(_04282_));
 sky130_fd_sc_hd__nand3_1 _11241_ (.A(_04282_),
    .B(_04274_),
    .C(_04276_),
    .Y(_04283_));
 sky130_fd_sc_hd__nand2_1 _11242_ (.A(_01858_),
    .B(_06231_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_1 _11243_ (.A(_06242_),
    .B(_06228_),
    .Y(_04285_));
 sky130_fd_sc_hd__or2_1 _11244_ (.A(_04284_),
    .B(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__nand2_1 _11245_ (.A(_04284_),
    .B(_04285_),
    .Y(_04287_));
 sky130_fd_sc_hd__nand2_1 _11246_ (.A(_04286_),
    .B(_04287_),
    .Y(_04288_));
 sky130_fd_sc_hd__nand2_1 _11247_ (.A(_06248_),
    .B(_06225_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_1 _11248_ (.A(_04288_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__inv_2 _11249_ (.A(_04289_),
    .Y(_04291_));
 sky130_fd_sc_hd__nand3_1 _11250_ (.A(_04286_),
    .B(_04291_),
    .C(_04287_),
    .Y(_04293_));
 sky130_fd_sc_hd__nand2_2 _11251_ (.A(_04290_),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand2_1 _11252_ (.A(_04070_),
    .B(_04066_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_1 _11253_ (.A(_06237_),
    .B(_06217_),
    .Y(_04296_));
 sky130_fd_sc_hd__inv_2 _11254_ (.A(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__nand2_1 _11255_ (.A(_06281_),
    .B(net38),
    .Y(_04298_));
 sky130_fd_sc_hd__inv_2 _11256_ (.A(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__nand2_1 _11257_ (.A(_04297_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__nand2_1 _11258_ (.A(_06234_),
    .B(_06220_),
    .Y(_04301_));
 sky130_fd_sc_hd__inv_2 _11259_ (.A(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__nand2_1 _11260_ (.A(_04296_),
    .B(_04298_),
    .Y(_04304_));
 sky130_fd_sc_hd__nand3_2 _11261_ (.A(_04300_),
    .B(_04302_),
    .C(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__nand2_1 _11262_ (.A(_04300_),
    .B(_04304_),
    .Y(_04306_));
 sky130_fd_sc_hd__nand2_1 _11263_ (.A(_04306_),
    .B(_04301_),
    .Y(_04307_));
 sky130_fd_sc_hd__nand3_1 _11264_ (.A(_04295_),
    .B(_04305_),
    .C(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__nand2_1 _11265_ (.A(_04307_),
    .B(_04305_),
    .Y(_04309_));
 sky130_fd_sc_hd__a21boi_1 _11266_ (.A1(_04068_),
    .A2(_04069_),
    .B1_N(_04066_),
    .Y(_04310_));
 sky130_fd_sc_hd__nand2_1 _11267_ (.A(_04309_),
    .B(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand3b_1 _11268_ (.A_N(_04294_),
    .B(_04308_),
    .C(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand2_1 _11269_ (.A(_04308_),
    .B(_04311_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _11270_ (.A(_04313_),
    .B(_04294_),
    .Y(_04315_));
 sky130_fd_sc_hd__nand2_1 _11271_ (.A(_04312_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_1 _11272_ (.A(_04036_),
    .B(_04038_),
    .Y(_04317_));
 sky130_fd_sc_hd__nor2_1 _11273_ (.A(_04038_),
    .B(_04036_),
    .Y(_04318_));
 sky130_fd_sc_hd__a21oi_2 _11274_ (.A1(_04317_),
    .A2(_04044_),
    .B1(_04318_),
    .Y(_04319_));
 sky130_fd_sc_hd__inv_2 _11275_ (.A(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand2_1 _11276_ (.A(_04316_),
    .B(_04320_),
    .Y(_04321_));
 sky130_fd_sc_hd__nand3_1 _11277_ (.A(_04319_),
    .B(_04312_),
    .C(_04315_),
    .Y(_04322_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(_04321_),
    .B(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__nand2_1 _11279_ (.A(_04092_),
    .B(_04073_),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _11280_ (.A(_04323_),
    .B(_04324_),
    .Y(_04326_));
 sky130_fd_sc_hd__nand3b_1 _11281_ (.A_N(_04324_),
    .B(_04321_),
    .C(_04322_),
    .Y(_04327_));
 sky130_fd_sc_hd__nand2_1 _11282_ (.A(_04326_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__nand3_1 _11283_ (.A(_04279_),
    .B(_04283_),
    .C(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__nand3_1 _11284_ (.A(_04278_),
    .B(_04274_),
    .C(_04276_),
    .Y(_04330_));
 sky130_fd_sc_hd__inv_2 _11285_ (.A(_04328_),
    .Y(_04331_));
 sky130_fd_sc_hd__nand2_1 _11286_ (.A(_04277_),
    .B(_04282_),
    .Y(_04332_));
 sky130_fd_sc_hd__nand3_1 _11287_ (.A(_04330_),
    .B(_04331_),
    .C(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__nand3_1 _11288_ (.A(_04214_),
    .B(_04329_),
    .C(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__nand2_1 _11289_ (.A(_04333_),
    .B(_04329_),
    .Y(_04335_));
 sky130_fd_sc_hd__a21o_1 _11290_ (.A1(_04109_),
    .A2(_04212_),
    .B1(_04213_),
    .X(_04337_));
 sky130_fd_sc_hd__nand2_1 _11291_ (.A(_04335_),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__or2_1 _11292_ (.A(_04139_),
    .B(_04137_),
    .X(_04339_));
 sky130_fd_sc_hd__nand2_1 _11293_ (.A(_04146_),
    .B(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hd__and2_1 _11294_ (.A(_04136_),
    .B(_04127_),
    .X(_04341_));
 sky130_fd_sc_hd__nand2_1 _11295_ (.A(net15),
    .B(_06199_),
    .Y(_04342_));
 sky130_fd_sc_hd__nand3b_2 _11296_ (.A_N(_04342_),
    .B(_06245_),
    .C(_06226_),
    .Y(_04343_));
 sky130_fd_sc_hd__inv_2 _11297_ (.A(_00270_),
    .Y(_04344_));
 sky130_fd_sc_hd__o21ai_1 _11298_ (.A1(_02871_),
    .A2(_04344_),
    .B1(_04342_),
    .Y(_04345_));
 sky130_fd_sc_hd__nand2_1 _11299_ (.A(_04343_),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__nand2_1 _11300_ (.A(_04346_),
    .B(_06413_),
    .Y(_04348_));
 sky130_fd_sc_hd__nand3_2 _11301_ (.A(_04343_),
    .B(_04345_),
    .C(_06202_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_1 _11302_ (.A(_04348_),
    .B(_04349_),
    .Y(_04350_));
 sky130_fd_sc_hd__a21boi_1 _11303_ (.A1(_04087_),
    .A2(_04082_),
    .B1_N(_04081_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2_1 _11304_ (.A(_04350_),
    .B(_04351_),
    .Y(_04352_));
 sky130_fd_sc_hd__nand2_1 _11305_ (.A(_04088_),
    .B(_04081_),
    .Y(_04353_));
 sky130_fd_sc_hd__nand3_1 _11306_ (.A(_04353_),
    .B(_04348_),
    .C(_04349_),
    .Y(_04354_));
 sky130_fd_sc_hd__nand2_1 _11307_ (.A(_04352_),
    .B(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__nand2_1 _11308_ (.A(_04124_),
    .B(_04122_),
    .Y(_04356_));
 sky130_fd_sc_hd__inv_2 _11309_ (.A(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__nand2_1 _11310_ (.A(_04355_),
    .B(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hd__nand3_1 _11311_ (.A(_04352_),
    .B(_04354_),
    .C(_04356_),
    .Y(_04359_));
 sky130_fd_sc_hd__nand2_1 _11312_ (.A(_04358_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__nor2_1 _11313_ (.A(_04341_),
    .B(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__nand2_1 _11314_ (.A(_04360_),
    .B(_04341_),
    .Y(_04362_));
 sky130_fd_sc_hd__nor2b_1 _11315_ (.A(_04361_),
    .B_N(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _11316_ (.A(_04093_),
    .B(_04097_),
    .Y(_04364_));
 sky130_fd_sc_hd__nor2_1 _11317_ (.A(_04097_),
    .B(_04093_),
    .Y(_04365_));
 sky130_fd_sc_hd__a21oi_1 _11318_ (.A1(_04364_),
    .A2(_04102_),
    .B1(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand2_1 _11319_ (.A(_04363_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__a21o_1 _11320_ (.A1(_04364_),
    .A2(_04102_),
    .B1(_04365_),
    .X(_04368_));
 sky130_fd_sc_hd__inv_2 _11321_ (.A(_04361_),
    .Y(_04369_));
 sky130_fd_sc_hd__nand2_1 _11322_ (.A(_04369_),
    .B(_04362_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_1 _11323_ (.A(_04368_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__nand3b_1 _11324_ (.A_N(_04340_),
    .B(_04367_),
    .C(_04371_),
    .Y(_04372_));
 sky130_fd_sc_hd__nand2_1 _11325_ (.A(_04363_),
    .B(_04368_),
    .Y(_04373_));
 sky130_fd_sc_hd__nand2_1 _11326_ (.A(_04370_),
    .B(_04366_),
    .Y(_04374_));
 sky130_fd_sc_hd__nand3_1 _11327_ (.A(_04373_),
    .B(_04374_),
    .C(_04340_),
    .Y(_04375_));
 sky130_fd_sc_hd__nand2_1 _11328_ (.A(_04372_),
    .B(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand3_1 _11329_ (.A(_04334_),
    .B(_04338_),
    .C(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand2_1 _11330_ (.A(_04334_),
    .B(_04338_),
    .Y(_04379_));
 sky130_fd_sc_hd__inv_2 _11331_ (.A(_04376_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2_1 _11332_ (.A(_04379_),
    .B(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__nand3_1 _11333_ (.A(_04211_),
    .B(_04377_),
    .C(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_1 _11334_ (.A(_04381_),
    .B(_04377_),
    .Y(_04383_));
 sky130_fd_sc_hd__a21o_1 _11335_ (.A1(_04166_),
    .A2(_04167_),
    .B1(_04210_),
    .X(_04384_));
 sky130_fd_sc_hd__nand2_1 _11336_ (.A(_04383_),
    .B(_04384_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _11337_ (.A(_04382_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__o21a_1 _11338_ (.A1(_04148_),
    .A2(_04152_),
    .B1(_04159_),
    .X(_04387_));
 sky130_fd_sc_hd__nor2_1 _11339_ (.A(_03904_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__nand2_1 _11340_ (.A(_04387_),
    .B(_03904_),
    .Y(_04389_));
 sky130_fd_sc_hd__and2b_1 _11341_ (.A_N(_04388_),
    .B(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__nand2_1 _11342_ (.A(_04386_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hd__or2b_1 _11343_ (.A(_04388_),
    .B_N(_04389_),
    .X(_04392_));
 sky130_fd_sc_hd__nand3_1 _11344_ (.A(_04382_),
    .B(_04385_),
    .C(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__nand2_1 _11345_ (.A(_04391_),
    .B(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hd__nor2_1 _11346_ (.A(_04174_),
    .B(_04172_),
    .Y(_04395_));
 sky130_fd_sc_hd__a21oi_2 _11347_ (.A1(_04175_),
    .A2(_04171_),
    .B1(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__inv_2 _11348_ (.A(_04396_),
    .Y(_04397_));
 sky130_fd_sc_hd__nand2_1 _11349_ (.A(_04394_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand3_1 _11350_ (.A(_04396_),
    .B(_04391_),
    .C(_04393_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_1 _11351_ (.A(_04398_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _11352_ (.A(_04401_),
    .B(_04180_),
    .Y(_04402_));
 sky130_fd_sc_hd__nand3_1 _11353_ (.A(_04398_),
    .B(_04400_),
    .C(_04179_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_1 _11354_ (.A(_04402_),
    .B(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hd__nand2_1 _11355_ (.A(_04184_),
    .B(_04186_),
    .Y(_04405_));
 sky130_fd_sc_hd__nor2_1 _11356_ (.A(_04186_),
    .B(_04184_),
    .Y(_04406_));
 sky130_fd_sc_hd__a21oi_1 _11357_ (.A1(_04405_),
    .A2(_03942_),
    .B1(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__inv_2 _11358_ (.A(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hd__nand2_1 _11359_ (.A(_04404_),
    .B(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__nand3_1 _11360_ (.A(_04407_),
    .B(_04403_),
    .C(_04402_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand2_1 _11361_ (.A(_04409_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hd__inv_2 _11362_ (.A(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__inv_2 _11363_ (.A(_03979_),
    .Y(_04414_));
 sky130_fd_sc_hd__nand3_1 _11364_ (.A(_04414_),
    .B(_04192_),
    .C(_04191_),
    .Y(_04415_));
 sky130_fd_sc_hd__nand2_2 _11365_ (.A(_04208_),
    .B(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__xor2_4 _11366_ (.A(_04413_),
    .B(_04416_),
    .X(\m1.out[29] ));
 sky130_fd_sc_hd__nand2_1 _11367_ (.A(_04394_),
    .B(_04396_),
    .Y(_04417_));
 sky130_fd_sc_hd__nor2_1 _11368_ (.A(_04396_),
    .B(_04394_),
    .Y(_04418_));
 sky130_fd_sc_hd__a21oi_2 _11369_ (.A1(_04417_),
    .A2(_04179_),
    .B1(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__nand2_1 _11370_ (.A(_04335_),
    .B(_04214_),
    .Y(_04421_));
 sky130_fd_sc_hd__nor2_1 _11371_ (.A(_04214_),
    .B(_04335_),
    .Y(_04422_));
 sky130_fd_sc_hd__a21o_1 _11372_ (.A1(_04421_),
    .A2(_04380_),
    .B1(_04422_),
    .X(_04423_));
 sky130_fd_sc_hd__nand2_1 _11373_ (.A(_04276_),
    .B(_04251_),
    .Y(_04424_));
 sky130_fd_sc_hd__nand2_1 _11374_ (.A(_04247_),
    .B(_04230_),
    .Y(_04425_));
 sky130_fd_sc_hd__inv_2 _11375_ (.A(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__a21o_1 _11376_ (.A1(_06290_),
    .A2(_06184_),
    .B1(_06264_),
    .X(_04427_));
 sky130_fd_sc_hd__nand3_1 _11377_ (.A(_06264_),
    .B(_06290_),
    .C(_06184_),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_1 _11378_ (.A(_04427_),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__nand2_1 _11379_ (.A(_06288_),
    .B(_02181_),
    .Y(_04430_));
 sky130_fd_sc_hd__nand2_1 _11380_ (.A(_04429_),
    .B(_04430_),
    .Y(_04432_));
 sky130_fd_sc_hd__inv_2 _11381_ (.A(_04430_),
    .Y(_04433_));
 sky130_fd_sc_hd__nand3_1 _11382_ (.A(_04427_),
    .B(_04433_),
    .C(_04428_),
    .Y(_04434_));
 sky130_fd_sc_hd__nand2_1 _11383_ (.A(_04432_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__nand2_1 _11384_ (.A(_04225_),
    .B(_04221_),
    .Y(_04436_));
 sky130_fd_sc_hd__inv_2 _11385_ (.A(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand2_1 _11386_ (.A(_04435_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__nand3_1 _11387_ (.A(_04432_),
    .B(_04436_),
    .C(_04434_),
    .Y(_04439_));
 sky130_fd_sc_hd__nand2_1 _11388_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__nand2_1 _11389_ (.A(_06291_),
    .B(_01692_),
    .Y(_04441_));
 sky130_fd_sc_hd__inv_2 _11390_ (.A(_04441_),
    .Y(_04443_));
 sky130_fd_sc_hd__nand2_1 _11391_ (.A(_06292_),
    .B(_01921_),
    .Y(_04444_));
 sky130_fd_sc_hd__inv_2 _11392_ (.A(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__nand2_1 _11393_ (.A(_04443_),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__nand2_1 _11394_ (.A(_04441_),
    .B(_04444_),
    .Y(_04447_));
 sky130_fd_sc_hd__nand2_1 _11395_ (.A(_06280_),
    .B(_06178_),
    .Y(_04448_));
 sky130_fd_sc_hd__inv_2 _11396_ (.A(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hd__a21o_1 _11397_ (.A1(_04446_),
    .A2(_04447_),
    .B1(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__nand3_1 _11398_ (.A(_04446_),
    .B(_04449_),
    .C(_04447_),
    .Y(_04451_));
 sky130_fd_sc_hd__nand2_1 _11399_ (.A(_04450_),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(_04440_),
    .B(_04452_),
    .Y(_04454_));
 sky130_fd_sc_hd__inv_2 _11401_ (.A(_04452_),
    .Y(_04455_));
 sky130_fd_sc_hd__nand3_2 _11402_ (.A(_04455_),
    .B(_04438_),
    .C(_04439_),
    .Y(_04456_));
 sky130_fd_sc_hd__nand2_1 _11403_ (.A(_04454_),
    .B(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__nand2_1 _11404_ (.A(_04426_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand3_2 _11405_ (.A(_04425_),
    .B(_04454_),
    .C(_04456_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2_1 _11406_ (.A(_04458_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_2 _11407_ (.A(_04262_),
    .B(_04255_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand2_1 _11408_ (.A(_01158_),
    .B(_01278_),
    .Y(_04462_));
 sky130_fd_sc_hd__inv_2 _11409_ (.A(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__nand2_1 _11410_ (.A(_00701_),
    .B(_06171_),
    .Y(_04465_));
 sky130_fd_sc_hd__inv_2 _11411_ (.A(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hd__nand2_1 _11412_ (.A(_04463_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _11413_ (.A(_04462_),
    .B(_04465_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand2_1 _11414_ (.A(_06282_),
    .B(_06222_),
    .Y(_04469_));
 sky130_fd_sc_hd__inv_2 _11415_ (.A(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__a21o_1 _11416_ (.A1(_04467_),
    .A2(_04468_),
    .B1(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__nand3_2 _11417_ (.A(_04467_),
    .B(_04470_),
    .C(_04468_),
    .Y(_04472_));
 sky130_fd_sc_hd__nand2_1 _11418_ (.A(_04471_),
    .B(_04472_),
    .Y(_04473_));
 sky130_fd_sc_hd__nand2_1 _11419_ (.A(_04243_),
    .B(_04236_),
    .Y(_04474_));
 sky130_fd_sc_hd__nand2_1 _11420_ (.A(_04473_),
    .B(_04474_),
    .Y(_04476_));
 sky130_fd_sc_hd__a21boi_1 _11421_ (.A1(_04242_),
    .A2(_04238_),
    .B1_N(_04236_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand3_1 _11422_ (.A(_04471_),
    .B(_04477_),
    .C(_04472_),
    .Y(_04478_));
 sky130_fd_sc_hd__nand3b_1 _11423_ (.A_N(_04461_),
    .B(_04476_),
    .C(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__nand2_1 _11424_ (.A(_04473_),
    .B(_04477_),
    .Y(_04480_));
 sky130_fd_sc_hd__nand3_1 _11425_ (.A(_04471_),
    .B(_04474_),
    .C(_04472_),
    .Y(_04481_));
 sky130_fd_sc_hd__nand3_1 _11426_ (.A(_04480_),
    .B(_04481_),
    .C(_04461_),
    .Y(_04482_));
 sky130_fd_sc_hd__nand2_1 _11427_ (.A(_04479_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_1 _11428_ (.A(_04460_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__inv_2 _11429_ (.A(_04483_),
    .Y(_04485_));
 sky130_fd_sc_hd__nand3_2 _11430_ (.A(_04485_),
    .B(_04458_),
    .C(_04459_),
    .Y(_04487_));
 sky130_fd_sc_hd__nand3_1 _11431_ (.A(_04424_),
    .B(_04484_),
    .C(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__nand2_1 _11432_ (.A(_04484_),
    .B(_04487_),
    .Y(_04489_));
 sky130_fd_sc_hd__a21boi_1 _11433_ (.A1(_04275_),
    .A2(_04250_),
    .B1_N(_04251_),
    .Y(_04490_));
 sky130_fd_sc_hd__nand2_1 _11434_ (.A(_04489_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand2_1 _11435_ (.A(_04488_),
    .B(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__nand2_1 _11436_ (.A(_02095_),
    .B(_06230_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand3b_1 _11437_ (.A_N(_04493_),
    .B(_06240_),
    .C(_06228_),
    .Y(_04494_));
 sky130_fd_sc_hd__inv_2 _11438_ (.A(_06239_),
    .Y(_04495_));
 sky130_fd_sc_hd__inv_2 _11439_ (.A(_00376_),
    .Y(_04496_));
 sky130_fd_sc_hd__o21ai_1 _11440_ (.A1(_04495_),
    .A2(_04496_),
    .B1(_04493_),
    .Y(_04498_));
 sky130_fd_sc_hd__nand2_1 _11441_ (.A(_04494_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__nand2_1 _11442_ (.A(_06246_),
    .B(_06225_),
    .Y(_04500_));
 sky130_fd_sc_hd__nand2_1 _11443_ (.A(_04499_),
    .B(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand3b_1 _11444_ (.A_N(_04500_),
    .B(_04494_),
    .C(_04498_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand2_1 _11445_ (.A(_04501_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_2 _11446_ (.A(_04305_),
    .B(_04300_),
    .Y(_04504_));
 sky130_fd_sc_hd__nand2_1 _11447_ (.A(_06235_),
    .B(_06218_),
    .Y(_04505_));
 sky130_fd_sc_hd__nand2_1 _11448_ (.A(_01211_),
    .B(_06223_),
    .Y(_04506_));
 sky130_fd_sc_hd__or2_1 _11449_ (.A(_04505_),
    .B(_04506_),
    .X(_04507_));
 sky130_fd_sc_hd__nand2_1 _11450_ (.A(_04505_),
    .B(_04506_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _11451_ (.A(_04507_),
    .B(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand2_1 _11452_ (.A(_06243_),
    .B(_06221_),
    .Y(_04511_));
 sky130_fd_sc_hd__nand2_1 _11453_ (.A(_04510_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__nand3b_1 _11454_ (.A_N(_04511_),
    .B(_04507_),
    .C(_04509_),
    .Y(_04513_));
 sky130_fd_sc_hd__nand3_1 _11455_ (.A(_04504_),
    .B(_04512_),
    .C(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__nand2_1 _11456_ (.A(_04512_),
    .B(_04513_),
    .Y(_04515_));
 sky130_fd_sc_hd__inv_2 _11457_ (.A(_04504_),
    .Y(_04516_));
 sky130_fd_sc_hd__nand2_1 _11458_ (.A(_04515_),
    .B(_04516_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand3b_2 _11459_ (.A_N(_04503_),
    .B(_04514_),
    .C(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__nand2_1 _11460_ (.A(_04517_),
    .B(_04514_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _11461_ (.A(_04520_),
    .B(_04503_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand2_1 _11462_ (.A(_04518_),
    .B(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__nand2_1 _11463_ (.A(_04263_),
    .B(_04264_),
    .Y(_04523_));
 sky130_fd_sc_hd__nor2_1 _11464_ (.A(_04264_),
    .B(_04263_),
    .Y(_04524_));
 sky130_fd_sc_hd__a21oi_2 _11465_ (.A1(_04523_),
    .A2(_04269_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__inv_2 _11466_ (.A(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__nand2_1 _11467_ (.A(_04522_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__nand3_1 _11468_ (.A(_04525_),
    .B(_04521_),
    .C(_04518_),
    .Y(_04528_));
 sky130_fd_sc_hd__nand2_1 _11469_ (.A(_04527_),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__nand2_1 _11470_ (.A(_04312_),
    .B(_04308_),
    .Y(_04531_));
 sky130_fd_sc_hd__nand2_1 _11471_ (.A(_04529_),
    .B(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__nand3b_1 _11472_ (.A_N(_04531_),
    .B(_04527_),
    .C(_04528_),
    .Y(_04533_));
 sky130_fd_sc_hd__nand2_1 _11473_ (.A(_04532_),
    .B(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _11474_ (.A(_04492_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__inv_2 _11475_ (.A(_04534_),
    .Y(_04536_));
 sky130_fd_sc_hd__nand3_2 _11476_ (.A(_04488_),
    .B(_04536_),
    .C(_04491_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_1 _11477_ (.A(_04535_),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_1 _11478_ (.A(_04333_),
    .B(_04330_),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _11479_ (.A(_04538_),
    .B(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__nor2_1 _11480_ (.A(_04282_),
    .B(_04277_),
    .Y(_04542_));
 sky130_fd_sc_hd__a21oi_1 _11481_ (.A1(_04332_),
    .A2(_04331_),
    .B1(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__nand3_1 _11482_ (.A(_04543_),
    .B(_04535_),
    .C(_04537_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand2_1 _11483_ (.A(_04316_),
    .B(_04319_),
    .Y(_04545_));
 sky130_fd_sc_hd__nor2_1 _11484_ (.A(_04319_),
    .B(_04316_),
    .Y(_04546_));
 sky130_fd_sc_hd__a21oi_2 _11485_ (.A1(_04545_),
    .A2(_04324_),
    .B1(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__inv_2 _11486_ (.A(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__and3_1 _11487_ (.A(_06298_),
    .B(_06200_),
    .C(_06226_),
    .X(_04549_));
 sky130_fd_sc_hd__inv_2 _11488_ (.A(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__a21o_1 _11489_ (.A1(_03905_),
    .A2(_06226_),
    .B1(_06200_),
    .X(_04551_));
 sky130_fd_sc_hd__nand2_1 _11490_ (.A(_04550_),
    .B(_04551_),
    .Y(_04553_));
 sky130_fd_sc_hd__a21o_1 _11491_ (.A1(_04293_),
    .A2(_04286_),
    .B1(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__nand3_1 _11492_ (.A(_04293_),
    .B(_04553_),
    .C(_04286_),
    .Y(_04555_));
 sky130_fd_sc_hd__nand2_1 _11493_ (.A(_04554_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__nand3_1 _11494_ (.A(_04556_),
    .B(_04343_),
    .C(_04349_),
    .Y(_04557_));
 sky130_fd_sc_hd__nand2_1 _11495_ (.A(_04349_),
    .B(_04343_),
    .Y(_04558_));
 sky130_fd_sc_hd__nand3_1 _11496_ (.A(_04554_),
    .B(_04555_),
    .C(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__nand2_1 _11497_ (.A(_04557_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_1 _11498_ (.A(_04359_),
    .B(_04354_),
    .Y(_04561_));
 sky130_fd_sc_hd__inv_2 _11499_ (.A(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__nand2_1 _11500_ (.A(_04560_),
    .B(_04562_),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_1 _11501_ (.A(_04562_),
    .B(_04560_),
    .Y(_04565_));
 sky130_fd_sc_hd__inv_2 _11502_ (.A(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hd__nand3_2 _11503_ (.A(_04548_),
    .B(_04564_),
    .C(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__nand2_1 _11504_ (.A(_04566_),
    .B(_04564_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand2_1 _11505_ (.A(_04568_),
    .B(_04547_),
    .Y(_04569_));
 sky130_fd_sc_hd__nand2_1 _11506_ (.A(_04567_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__nand2_1 _11507_ (.A(_04570_),
    .B(_04369_),
    .Y(_04571_));
 sky130_fd_sc_hd__nand3_1 _11508_ (.A(_04567_),
    .B(_04569_),
    .C(_04361_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand2_1 _11509_ (.A(_04571_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__nand3_1 _11510_ (.A(_04540_),
    .B(_04544_),
    .C(_04573_),
    .Y(_04575_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(_04540_),
    .B(_04544_),
    .Y(_04576_));
 sky130_fd_sc_hd__inv_2 _11512_ (.A(_04573_),
    .Y(_04577_));
 sky130_fd_sc_hd__nand2_1 _11513_ (.A(_04576_),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand3_1 _11514_ (.A(_04423_),
    .B(_04575_),
    .C(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__nand2_1 _11515_ (.A(_04578_),
    .B(_04575_),
    .Y(_04580_));
 sky130_fd_sc_hd__a21oi_1 _11516_ (.A1(_04421_),
    .A2(_04380_),
    .B1(_04422_),
    .Y(_04581_));
 sky130_fd_sc_hd__nand2_1 _11517_ (.A(_04580_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_2 _11518_ (.A(_04375_),
    .B(_04373_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand3_1 _11519_ (.A(_04579_),
    .B(_04582_),
    .C(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__nand2_1 _11520_ (.A(_04580_),
    .B(_04423_),
    .Y(_04586_));
 sky130_fd_sc_hd__nand3_1 _11521_ (.A(_04581_),
    .B(_04578_),
    .C(_04575_),
    .Y(_04587_));
 sky130_fd_sc_hd__inv_2 _11522_ (.A(_04583_),
    .Y(_04588_));
 sky130_fd_sc_hd__nand3_1 _11523_ (.A(_04586_),
    .B(_04587_),
    .C(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__nand2_1 _11524_ (.A(_04584_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _11525_ (.A(_04383_),
    .B(_04211_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2_1 _11526_ (.A(_04211_),
    .B(_04383_),
    .Y(_04592_));
 sky130_fd_sc_hd__a21oi_2 _11527_ (.A1(_04591_),
    .A2(_04390_),
    .B1(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__inv_2 _11528_ (.A(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _11529_ (.A(_04590_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand3_1 _11530_ (.A(_04593_),
    .B(_04584_),
    .C(_04589_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _11531_ (.A(_04595_),
    .B(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_1 _11532_ (.A(_04598_),
    .B(_04388_),
    .Y(_04599_));
 sky130_fd_sc_hd__nand3b_1 _11533_ (.A_N(_04388_),
    .B(_04595_),
    .C(_04597_),
    .Y(_04600_));
 sky130_fd_sc_hd__nand2_1 _11534_ (.A(_04599_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__nor2_1 _11535_ (.A(_04419_),
    .B(_04601_),
    .Y(_04602_));
 sky130_fd_sc_hd__nand2_1 _11536_ (.A(_04601_),
    .B(_04419_),
    .Y(_04603_));
 sky130_fd_sc_hd__inv_2 _11537_ (.A(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__nor2_1 _11538_ (.A(_04602_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__nand2_1 _11539_ (.A(_04415_),
    .B(_04196_),
    .Y(_04606_));
 sky130_fd_sc_hd__nor2_1 _11540_ (.A(_04412_),
    .B(_04606_),
    .Y(_04608_));
 sky130_fd_sc_hd__nand3_1 _11541_ (.A(_04195_),
    .B(_04409_),
    .C(_04411_),
    .Y(_04609_));
 sky130_fd_sc_hd__nand2_1 _11542_ (.A(_04609_),
    .B(_04409_),
    .Y(_04610_));
 sky130_fd_sc_hd__a21o_1 _11543_ (.A1(_04206_),
    .A2(_04608_),
    .B1(_04610_),
    .X(_04611_));
 sky130_fd_sc_hd__or2_1 _11544_ (.A(_04605_),
    .B(_04611_),
    .X(_04612_));
 sky130_fd_sc_hd__nand2_1 _11545_ (.A(_04611_),
    .B(_04605_),
    .Y(_04613_));
 sky130_fd_sc_hd__and2_1 _11546_ (.A(_04612_),
    .B(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__buf_6 _11547_ (.A(_04614_),
    .X(\m1.out[30] ));
 sky130_fd_sc_hd__inv_2 _11548_ (.A(_04419_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand3_1 _11549_ (.A(_04615_),
    .B(_04600_),
    .C(_04599_),
    .Y(_04616_));
 sky130_fd_sc_hd__nand2_1 _11550_ (.A(_04613_),
    .B(_04616_),
    .Y(_04618_));
 sky130_fd_sc_hd__nand2_1 _11551_ (.A(_04590_),
    .B(_04593_),
    .Y(_04619_));
 sky130_fd_sc_hd__nor2_1 _11552_ (.A(_04593_),
    .B(_04590_),
    .Y(_04620_));
 sky130_fd_sc_hd__a21oi_1 _11553_ (.A1(_04619_),
    .A2(_04388_),
    .B1(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__inv_2 _11554_ (.A(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__and2_1 _11555_ (.A(_04502_),
    .B(_04494_),
    .X(_04623_));
 sky130_fd_sc_hd__or2_1 _11556_ (.A(_04344_),
    .B(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__nand2_1 _11557_ (.A(_04623_),
    .B(_04344_),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_1 _11558_ (.A(_04624_),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__nand2_1 _11559_ (.A(_04626_),
    .B(_04550_),
    .Y(_04627_));
 sky130_fd_sc_hd__nand3_1 _11560_ (.A(_04624_),
    .B(_04549_),
    .C(_04625_),
    .Y(_04629_));
 sky130_fd_sc_hd__nand2_1 _11561_ (.A(_04627_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _11562_ (.A(_04559_),
    .B(_04554_),
    .Y(_04631_));
 sky130_fd_sc_hd__inv_2 _11563_ (.A(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand2_1 _11564_ (.A(_04630_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__nand3_2 _11565_ (.A(_04627_),
    .B(_04631_),
    .C(_04629_),
    .Y(_04634_));
 sky130_fd_sc_hd__nand2_1 _11566_ (.A(_04633_),
    .B(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__o21ai_1 _11567_ (.A1(_04522_),
    .A2(_04525_),
    .B1(_04532_),
    .Y(_04636_));
 sky130_fd_sc_hd__nand2b_2 _11568_ (.A_N(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__or2_1 _11569_ (.A(_04525_),
    .B(_04522_),
    .X(_04638_));
 sky130_fd_sc_hd__nand3_1 _11570_ (.A(_04635_),
    .B(_04638_),
    .C(_04532_),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2_1 _11571_ (.A(_04637_),
    .B(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand2_1 _11572_ (.A(_04641_),
    .B(_04566_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand3_2 _11573_ (.A(_04637_),
    .B(_04640_),
    .C(_04565_),
    .Y(_04643_));
 sky130_fd_sc_hd__nand2_1 _11574_ (.A(_04642_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__inv_2 _11575_ (.A(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__nand2_1 _11576_ (.A(_06279_),
    .B(_06179_),
    .Y(_04646_));
 sky130_fd_sc_hd__nand2_1 _11577_ (.A(_00849_),
    .B(_06175_),
    .Y(_04647_));
 sky130_fd_sc_hd__nand2_1 _11578_ (.A(_00561_),
    .B(_01921_),
    .Y(_04648_));
 sky130_fd_sc_hd__or2_1 _11579_ (.A(_04647_),
    .B(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__nand2_1 _11580_ (.A(_04647_),
    .B(_04648_),
    .Y(_04651_));
 sky130_fd_sc_hd__nand2_1 _11581_ (.A(_04649_),
    .B(_04651_),
    .Y(_04652_));
 sky130_fd_sc_hd__or2_1 _11582_ (.A(_04646_),
    .B(_04652_),
    .X(_04653_));
 sky130_fd_sc_hd__nand2_1 _11583_ (.A(_04652_),
    .B(_04646_),
    .Y(_04654_));
 sky130_fd_sc_hd__nand2_1 _11584_ (.A(_04653_),
    .B(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__a21o_1 _11585_ (.A1(_06288_),
    .A2(_06184_),
    .B1(_06290_),
    .X(_04656_));
 sky130_fd_sc_hd__nand3_1 _11586_ (.A(_06288_),
    .B(_06290_),
    .C(_06184_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _11587_ (.A(_04656_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__nand2_1 _11588_ (.A(_06292_),
    .B(_02181_),
    .Y(_04659_));
 sky130_fd_sc_hd__nand2_1 _11589_ (.A(_04658_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__nand3b_1 _11590_ (.A_N(_04659_),
    .B(_04656_),
    .C(_04657_),
    .Y(_04662_));
 sky130_fd_sc_hd__nand2_1 _11591_ (.A(_04660_),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__a21boi_2 _11592_ (.A1(_04427_),
    .A2(_04433_),
    .B1_N(_04428_),
    .Y(_04664_));
 sky130_fd_sc_hd__nand2_1 _11593_ (.A(_04663_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__nor2_1 _11594_ (.A(_04664_),
    .B(_04663_),
    .Y(_04666_));
 sky130_fd_sc_hd__inv_2 _11595_ (.A(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__nand3b_1 _11596_ (.A_N(_04655_),
    .B(_04665_),
    .C(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__nand2_1 _11597_ (.A(_04667_),
    .B(_04665_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand2_1 _11598_ (.A(_04669_),
    .B(_04655_),
    .Y(_04670_));
 sky130_fd_sc_hd__nand2_1 _11599_ (.A(_04668_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__nand2_1 _11600_ (.A(_04456_),
    .B(_04439_),
    .Y(_04673_));
 sky130_fd_sc_hd__inv_2 _11601_ (.A(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__nand2_1 _11602_ (.A(_04671_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand3_1 _11603_ (.A(_04668_),
    .B(_04670_),
    .C(_04673_),
    .Y(_04676_));
 sky130_fd_sc_hd__nand2_1 _11604_ (.A(_04675_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2_1 _11605_ (.A(_04472_),
    .B(_04467_),
    .Y(_04678_));
 sky130_fd_sc_hd__nand2_1 _11606_ (.A(_06282_),
    .B(_06174_),
    .Y(_04679_));
 sky130_fd_sc_hd__nand2_1 _11607_ (.A(_06284_),
    .B(_06172_),
    .Y(_04680_));
 sky130_fd_sc_hd__or2_1 _11608_ (.A(_04679_),
    .B(_04680_),
    .X(_04681_));
 sky130_fd_sc_hd__nand2_1 _11609_ (.A(_04679_),
    .B(_04680_),
    .Y(_04682_));
 sky130_fd_sc_hd__nand2_1 _11610_ (.A(_04681_),
    .B(_04682_),
    .Y(_04684_));
 sky130_fd_sc_hd__nand2_1 _11611_ (.A(_06238_),
    .B(_06222_),
    .Y(_04685_));
 sky130_fd_sc_hd__inv_2 _11612_ (.A(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__or2b_1 _11613_ (.A(_04684_),
    .B_N(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__nand2_1 _11614_ (.A(_04684_),
    .B(_04685_),
    .Y(_04688_));
 sky130_fd_sc_hd__nand2_1 _11615_ (.A(_04687_),
    .B(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__nand2_1 _11616_ (.A(_04451_),
    .B(_04446_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand2_1 _11617_ (.A(_04689_),
    .B(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__inv_2 _11618_ (.A(_04690_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand3_1 _11619_ (.A(_04687_),
    .B(_04692_),
    .C(_04688_),
    .Y(_04693_));
 sky130_fd_sc_hd__nand3b_1 _11620_ (.A_N(_04678_),
    .B(_04691_),
    .C(_04693_),
    .Y(_04695_));
 sky130_fd_sc_hd__nand2_1 _11621_ (.A(_04689_),
    .B(_04692_),
    .Y(_04696_));
 sky130_fd_sc_hd__nand3_1 _11622_ (.A(_04687_),
    .B(_04688_),
    .C(_04690_),
    .Y(_04697_));
 sky130_fd_sc_hd__nand3_1 _11623_ (.A(_04696_),
    .B(_04678_),
    .C(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__nand2_1 _11624_ (.A(_04695_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__nand2_1 _11625_ (.A(_04677_),
    .B(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__inv_2 _11626_ (.A(_04699_),
    .Y(_04701_));
 sky130_fd_sc_hd__nand3_1 _11627_ (.A(_04675_),
    .B(_04676_),
    .C(_04701_),
    .Y(_04702_));
 sky130_fd_sc_hd__nand2_1 _11628_ (.A(_04700_),
    .B(_04702_),
    .Y(_04703_));
 sky130_fd_sc_hd__nand2_2 _11629_ (.A(_04487_),
    .B(_04459_),
    .Y(_04704_));
 sky130_fd_sc_hd__inv_2 _11630_ (.A(_04704_),
    .Y(_04706_));
 sky130_fd_sc_hd__nand2_1 _11631_ (.A(_04703_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__nand3_1 _11632_ (.A(_04700_),
    .B(_04704_),
    .C(_04702_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand2_1 _11633_ (.A(_04707_),
    .B(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__nand2_1 _11634_ (.A(_06240_),
    .B(_06221_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_1 _11635_ (.A(_06242_),
    .B(_00926_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand2_1 _11636_ (.A(_06235_),
    .B(_06223_),
    .Y(_04712_));
 sky130_fd_sc_hd__or2_1 _11637_ (.A(_04711_),
    .B(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(_04711_),
    .B(_04712_),
    .Y(_04714_));
 sky130_fd_sc_hd__nand2_1 _11639_ (.A(_04713_),
    .B(_04714_),
    .Y(_04715_));
 sky130_fd_sc_hd__or2_1 _11640_ (.A(_04710_),
    .B(_04715_),
    .X(_04717_));
 sky130_fd_sc_hd__nand2_1 _11641_ (.A(_04715_),
    .B(_04710_),
    .Y(_04718_));
 sky130_fd_sc_hd__nand2_1 _11642_ (.A(_04717_),
    .B(_04718_),
    .Y(_04719_));
 sky130_fd_sc_hd__nand2_1 _11643_ (.A(_04513_),
    .B(_04507_),
    .Y(_04720_));
 sky130_fd_sc_hd__inv_2 _11644_ (.A(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2_1 _11645_ (.A(_04719_),
    .B(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand3_1 _11646_ (.A(_04717_),
    .B(_04720_),
    .C(_04718_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand2_1 _11647_ (.A(_04722_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__nand2_1 _11648_ (.A(_06245_),
    .B(_06231_),
    .Y(_04725_));
 sky130_fd_sc_hd__nand2_1 _11649_ (.A(_06248_),
    .B(_06228_),
    .Y(_04726_));
 sky130_fd_sc_hd__or2_1 _11650_ (.A(_04725_),
    .B(_04726_),
    .X(_04728_));
 sky130_fd_sc_hd__nand2_1 _11651_ (.A(_04725_),
    .B(_04726_),
    .Y(_04729_));
 sky130_fd_sc_hd__nand2_1 _11652_ (.A(_04728_),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand3b_1 _11653_ (.A_N(_04730_),
    .B(_06299_),
    .C(_06225_),
    .Y(_04731_));
 sky130_fd_sc_hd__inv_2 _11654_ (.A(_06225_),
    .Y(_04732_));
 sky130_fd_sc_hd__o21ai_1 _11655_ (.A1(_06250_),
    .A2(_04732_),
    .B1(_04730_),
    .Y(_04733_));
 sky130_fd_sc_hd__nand2_1 _11656_ (.A(_04731_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__nand2_1 _11657_ (.A(_04724_),
    .B(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__inv_2 _11658_ (.A(_04734_),
    .Y(_04736_));
 sky130_fd_sc_hd__nand3_1 _11659_ (.A(_04736_),
    .B(_04722_),
    .C(_04723_),
    .Y(_04737_));
 sky130_fd_sc_hd__nand2_1 _11660_ (.A(_04735_),
    .B(_04737_),
    .Y(_04739_));
 sky130_fd_sc_hd__a21boi_4 _11661_ (.A1(_04480_),
    .A2(_04461_),
    .B1_N(_04481_),
    .Y(_04740_));
 sky130_fd_sc_hd__inv_2 _11662_ (.A(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand2_1 _11663_ (.A(_04739_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand3_1 _11664_ (.A(_04735_),
    .B(_04737_),
    .C(_04740_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _11665_ (.A(_04742_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2_1 _11666_ (.A(_04518_),
    .B(_04514_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_1 _11667_ (.A(_04744_),
    .B(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__nand3b_1 _11668_ (.A_N(_04745_),
    .B(_04742_),
    .C(_04743_),
    .Y(_04747_));
 sky130_fd_sc_hd__nand2_1 _11669_ (.A(_04746_),
    .B(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__nand2_1 _11670_ (.A(_04709_),
    .B(_04748_),
    .Y(_04750_));
 sky130_fd_sc_hd__inv_2 _11671_ (.A(_04748_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand3_2 _11672_ (.A(_04707_),
    .B(_04751_),
    .C(_04708_),
    .Y(_04752_));
 sky130_fd_sc_hd__nand2_1 _11673_ (.A(_04750_),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand2_1 _11674_ (.A(_04537_),
    .B(_04488_),
    .Y(_04754_));
 sky130_fd_sc_hd__inv_2 _11675_ (.A(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _11676_ (.A(_04753_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand3_1 _11677_ (.A(_04750_),
    .B(_04752_),
    .C(_04754_),
    .Y(_04757_));
 sky130_fd_sc_hd__nand3_1 _11678_ (.A(_04645_),
    .B(_04756_),
    .C(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _11679_ (.A(_04756_),
    .B(_04757_),
    .Y(_04759_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(_04759_),
    .B(_04644_),
    .Y(_04761_));
 sky130_fd_sc_hd__nand2_1 _11681_ (.A(_04758_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__nand3_1 _11682_ (.A(_04539_),
    .B(_04535_),
    .C(_04537_),
    .Y(_04763_));
 sky130_fd_sc_hd__nand2_1 _11683_ (.A(_04578_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__inv_2 _11684_ (.A(_04764_),
    .Y(_04765_));
 sky130_fd_sc_hd__nand2_1 _11685_ (.A(_04762_),
    .B(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__nand3_1 _11686_ (.A(_04758_),
    .B(_04761_),
    .C(_04764_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _11687_ (.A(_04766_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__nand3_2 _11688_ (.A(_04768_),
    .B(_04567_),
    .C(_04572_),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_1 _11689_ (.A(_04572_),
    .B(_04567_),
    .Y(_04770_));
 sky130_fd_sc_hd__nand3_2 _11690_ (.A(_04766_),
    .B(_04767_),
    .C(_04770_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand2_1 _11691_ (.A(_04769_),
    .B(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__inv_2 _11692_ (.A(_04579_),
    .Y(_04774_));
 sky130_fd_sc_hd__a21oi_2 _11693_ (.A1(_04582_),
    .A2(_04583_),
    .B1(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__inv_2 _11694_ (.A(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nand2_1 _11695_ (.A(_04773_),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand3_1 _11696_ (.A(_04769_),
    .B(_04772_),
    .C(_04775_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_1 _11697_ (.A(_04777_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__nand2_1 _11698_ (.A(_04622_),
    .B(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _11699_ (.A(_04773_),
    .B(_04775_),
    .Y(_04781_));
 sky130_fd_sc_hd__nand3_4 _11700_ (.A(_04769_),
    .B(_04776_),
    .C(_04772_),
    .Y(_04783_));
 sky130_fd_sc_hd__nand2_1 _11701_ (.A(_04781_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__nand2_1 _11702_ (.A(_04784_),
    .B(_04621_),
    .Y(_04785_));
 sky130_fd_sc_hd__nand2_1 _11703_ (.A(_04780_),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand2_1 _11704_ (.A(_04618_),
    .B(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__inv_2 _11705_ (.A(_04786_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand3_1 _11706_ (.A(_04613_),
    .B(_04616_),
    .C(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__nand2_2 _11707_ (.A(_04787_),
    .B(_04789_),
    .Y(\m1.out[31] ));
 sky130_fd_sc_hd__and2_2 _11708_ (.A(_04758_),
    .B(_04757_),
    .X(_04790_));
 sky130_fd_sc_hd__and2_1 _11709_ (.A(_04752_),
    .B(_04708_),
    .X(_04791_));
 sky130_fd_sc_hd__and2_1 _11710_ (.A(_04702_),
    .B(_04676_),
    .X(_04793_));
 sky130_fd_sc_hd__nand2_1 _11711_ (.A(_06284_),
    .B(_06179_),
    .Y(_04794_));
 sky130_fd_sc_hd__and4_1 _11712_ (.A(_06279_),
    .B(_06280_),
    .C(_06176_),
    .D(_01922_),
    .X(_04795_));
 sky130_fd_sc_hd__a22o_1 _11713_ (.A1(_06279_),
    .A2(_06176_),
    .B1(_06280_),
    .B2(_01922_),
    .X(_04796_));
 sky130_fd_sc_hd__inv_2 _11714_ (.A(_04796_),
    .Y(_04797_));
 sky130_fd_sc_hd__nor2_1 _11715_ (.A(_04795_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__xor2_1 _11716_ (.A(_04794_),
    .B(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__inv_2 _11717_ (.A(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__inv_2 _11718_ (.A(net47),
    .Y(_04801_));
 sky130_fd_sc_hd__or3_2 _11719_ (.A(_00329_),
    .B(_00330_),
    .C(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__a21o_1 _11720_ (.A1(_06292_),
    .A2(_06184_),
    .B1(_06288_),
    .X(_04804_));
 sky130_fd_sc_hd__nand2_1 _11721_ (.A(_04802_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__nand2_1 _11722_ (.A(_06291_),
    .B(_02181_),
    .Y(_04806_));
 sky130_fd_sc_hd__nand2_1 _11723_ (.A(_04805_),
    .B(_04806_),
    .Y(_04807_));
 sky130_fd_sc_hd__nand3b_2 _11724_ (.A_N(_04806_),
    .B(_04802_),
    .C(_04804_),
    .Y(_04808_));
 sky130_fd_sc_hd__nand2_1 _11725_ (.A(_04807_),
    .B(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__nand2_1 _11726_ (.A(_04662_),
    .B(_04657_),
    .Y(_04810_));
 sky130_fd_sc_hd__inv_2 _11727_ (.A(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__nand2_1 _11728_ (.A(_04809_),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__nand3_1 _11729_ (.A(_04807_),
    .B(_04808_),
    .C(_04810_),
    .Y(_04813_));
 sky130_fd_sc_hd__nand3_1 _11730_ (.A(_04800_),
    .B(_04812_),
    .C(_04813_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_1 _11731_ (.A(_04812_),
    .B(_04813_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _11732_ (.A(_04816_),
    .B(_04799_),
    .Y(_04817_));
 sky130_fd_sc_hd__nand2_1 _11733_ (.A(_04815_),
    .B(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__a31oi_2 _11734_ (.A1(_04665_),
    .A2(_04653_),
    .A3(_04654_),
    .B1(_04666_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _11735_ (.A(_04818_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand3b_2 _11736_ (.A_N(_04819_),
    .B(_04815_),
    .C(_04817_),
    .Y(_04821_));
 sky130_fd_sc_hd__nand2_1 _11737_ (.A(_04820_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand2_1 _11738_ (.A(_04687_),
    .B(_04681_),
    .Y(_04823_));
 sky130_fd_sc_hd__and4_1 _11739_ (.A(_06282_),
    .B(_06238_),
    .C(_06171_),
    .D(_06174_),
    .X(_04824_));
 sky130_fd_sc_hd__a22o_1 _11740_ (.A1(_01831_),
    .A2(_01280_),
    .B1(_01211_),
    .B2(_01278_),
    .X(_04826_));
 sky130_fd_sc_hd__inv_2 _11741_ (.A(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__nand2_1 _11742_ (.A(_06236_),
    .B(_06222_),
    .Y(_04828_));
 sky130_fd_sc_hd__o21ai_1 _11743_ (.A1(_04824_),
    .A2(_04827_),
    .B1(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__nor2_1 _11744_ (.A(_04824_),
    .B(_04827_),
    .Y(_04830_));
 sky130_fd_sc_hd__inv_2 _11745_ (.A(_04828_),
    .Y(_04831_));
 sky130_fd_sc_hd__nand2_1 _11746_ (.A(_04830_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__nand2_1 _11747_ (.A(_04829_),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__and2_1 _11748_ (.A(_04653_),
    .B(_04649_),
    .X(_04834_));
 sky130_fd_sc_hd__nand2b_1 _11749_ (.A_N(_04833_),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__or2b_1 _11750_ (.A(_04834_),
    .B_N(_04833_),
    .X(_04837_));
 sky130_fd_sc_hd__nand3b_1 _11751_ (.A_N(_04823_),
    .B(_04835_),
    .C(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__nor2_1 _11752_ (.A(_04834_),
    .B(_04833_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand2_1 _11753_ (.A(_04833_),
    .B(_04834_),
    .Y(_04840_));
 sky130_fd_sc_hd__nand3b_1 _11754_ (.A_N(_04839_),
    .B(_04823_),
    .C(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__nand2_1 _11755_ (.A(_04838_),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__nand2_1 _11756_ (.A(_04822_),
    .B(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__inv_2 _11757_ (.A(_04842_),
    .Y(_04844_));
 sky130_fd_sc_hd__nand3_2 _11758_ (.A(_04844_),
    .B(_04820_),
    .C(_04821_),
    .Y(_04845_));
 sky130_fd_sc_hd__nand3b_2 _11759_ (.A_N(_04793_),
    .B(_04843_),
    .C(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_1 _11760_ (.A(_04845_),
    .B(_04843_),
    .Y(_04848_));
 sky130_fd_sc_hd__nand2_1 _11761_ (.A(_04848_),
    .B(_04793_),
    .Y(_04849_));
 sky130_fd_sc_hd__nand2_1 _11762_ (.A(_04846_),
    .B(_04849_),
    .Y(_04850_));
 sky130_fd_sc_hd__and2_1 _11763_ (.A(_04717_),
    .B(_04713_),
    .X(_04851_));
 sky130_fd_sc_hd__nand2_1 _11764_ (.A(_06248_),
    .B(_06221_),
    .Y(_04852_));
 sky130_fd_sc_hd__inv_2 _11765_ (.A(net10),
    .Y(_04853_));
 sky130_fd_sc_hd__inv_2 _11766_ (.A(_06223_),
    .Y(_04854_));
 sky130_fd_sc_hd__nand2_1 _11767_ (.A(_06240_),
    .B(_06218_),
    .Y(_04855_));
 sky130_fd_sc_hd__nor3_1 _11768_ (.A(_04853_),
    .B(_04854_),
    .C(_04855_),
    .Y(_04856_));
 sky130_fd_sc_hd__inv_2 _11769_ (.A(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__o21ai_1 _11770_ (.A1(_04853_),
    .A2(_04854_),
    .B1(_04855_),
    .Y(_04859_));
 sky130_fd_sc_hd__nand2_1 _11771_ (.A(_04857_),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__or2_1 _11772_ (.A(_04852_),
    .B(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__nand2_1 _11773_ (.A(_04860_),
    .B(_04852_),
    .Y(_04862_));
 sky130_fd_sc_hd__nand2_1 _11774_ (.A(_04861_),
    .B(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hd__nor2_1 _11775_ (.A(_04851_),
    .B(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__and4_1 _11776_ (.A(_06246_),
    .B(_03905_),
    .C(_06228_),
    .D(_06231_),
    .X(_04865_));
 sky130_fd_sc_hd__a22o_1 _11777_ (.A1(_06247_),
    .A2(_06228_),
    .B1(_06299_),
    .B2(_06231_),
    .X(_04866_));
 sky130_fd_sc_hd__nor2b_1 _11778_ (.A(_04865_),
    .B_N(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__xor2_1 _11779_ (.A(_04732_),
    .B(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__inv_2 _11780_ (.A(_04868_),
    .Y(_04870_));
 sky130_fd_sc_hd__nand2_1 _11781_ (.A(_04863_),
    .B(_04851_),
    .Y(_04871_));
 sky130_fd_sc_hd__nand3b_1 _11782_ (.A_N(_04864_),
    .B(_04870_),
    .C(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hd__nand2b_1 _11783_ (.A_N(_04863_),
    .B(_04851_),
    .Y(_04873_));
 sky130_fd_sc_hd__nand2b_1 _11784_ (.A_N(_04851_),
    .B(_04863_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand3_1 _11785_ (.A(_04873_),
    .B(_04874_),
    .C(_04868_),
    .Y(_04875_));
 sky130_fd_sc_hd__nand2_1 _11786_ (.A(_04872_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__nand2_1 _11787_ (.A(_04698_),
    .B(_04697_),
    .Y(_04877_));
 sky130_fd_sc_hd__nand2_1 _11788_ (.A(_04876_),
    .B(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__inv_2 _11789_ (.A(_04877_),
    .Y(_04879_));
 sky130_fd_sc_hd__nand3_1 _11790_ (.A(_04872_),
    .B(_04875_),
    .C(_04879_),
    .Y(_04881_));
 sky130_fd_sc_hd__nand2_1 _11791_ (.A(_04878_),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__nand2_1 _11792_ (.A(_04737_),
    .B(_04723_),
    .Y(_04883_));
 sky130_fd_sc_hd__nand2_1 _11793_ (.A(_04882_),
    .B(_04883_),
    .Y(_04884_));
 sky130_fd_sc_hd__nand3b_1 _11794_ (.A_N(_04883_),
    .B(_04878_),
    .C(_04881_),
    .Y(_04885_));
 sky130_fd_sc_hd__nand2_1 _11795_ (.A(_04884_),
    .B(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__nand2_1 _11796_ (.A(_04850_),
    .B(_04886_),
    .Y(_04887_));
 sky130_fd_sc_hd__inv_2 _11797_ (.A(_04886_),
    .Y(_04888_));
 sky130_fd_sc_hd__nand3_1 _11798_ (.A(_04846_),
    .B(_04888_),
    .C(_04849_),
    .Y(_04889_));
 sky130_fd_sc_hd__nand3b_2 _11799_ (.A_N(_04791_),
    .B(_04887_),
    .C(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand2_1 _11800_ (.A(_04887_),
    .B(_04889_),
    .Y(_04892_));
 sky130_fd_sc_hd__nand2_1 _11801_ (.A(_04892_),
    .B(_04791_),
    .Y(_04893_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(_04890_),
    .B(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hd__and2_1 _11803_ (.A(_04731_),
    .B(_04728_),
    .X(_04895_));
 sky130_fd_sc_hd__and2_1 _11804_ (.A(_04629_),
    .B(_04624_),
    .X(_04896_));
 sky130_fd_sc_hd__nor2_1 _11805_ (.A(_04895_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__inv_2 _11806_ (.A(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand2_1 _11807_ (.A(_04896_),
    .B(_04895_),
    .Y(_04899_));
 sky130_fd_sc_hd__nand2_1 _11808_ (.A(_04898_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__or2_1 _11809_ (.A(_04740_),
    .B(_04739_),
    .X(_04901_));
 sky130_fd_sc_hd__and2_1 _11810_ (.A(_04746_),
    .B(_04901_),
    .X(_04903_));
 sky130_fd_sc_hd__nor2_1 _11811_ (.A(_04900_),
    .B(_04903_),
    .Y(_04904_));
 sky130_fd_sc_hd__inv_2 _11812_ (.A(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__nand2_1 _11813_ (.A(_04903_),
    .B(_04900_),
    .Y(_04906_));
 sky130_fd_sc_hd__nand2_1 _11814_ (.A(_04905_),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hd__nand2_1 _11815_ (.A(_04907_),
    .B(_04634_),
    .Y(_04908_));
 sky130_fd_sc_hd__inv_2 _11816_ (.A(_04634_),
    .Y(_04909_));
 sky130_fd_sc_hd__nand3_1 _11817_ (.A(_04905_),
    .B(_04909_),
    .C(_04906_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand2_1 _11818_ (.A(_04908_),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__nand2_1 _11819_ (.A(_04894_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__inv_2 _11820_ (.A(_04911_),
    .Y(_04914_));
 sky130_fd_sc_hd__nand3_1 _11821_ (.A(_04890_),
    .B(_04893_),
    .C(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__nand3b_2 _11822_ (.A_N(_04790_),
    .B(_04912_),
    .C(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__nand2_1 _11823_ (.A(_04912_),
    .B(_04915_),
    .Y(_04917_));
 sky130_fd_sc_hd__nand2_1 _11824_ (.A(_04917_),
    .B(_04790_),
    .Y(_04918_));
 sky130_fd_sc_hd__nand2_1 _11825_ (.A(_04916_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__nand2_4 _11826_ (.A(_04643_),
    .B(_04637_),
    .Y(_04920_));
 sky130_fd_sc_hd__inv_2 _11827_ (.A(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_1 _11828_ (.A(_04919_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__nand3_1 _11829_ (.A(_04916_),
    .B(_04918_),
    .C(_04920_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand2_1 _11830_ (.A(_04922_),
    .B(_04923_),
    .Y(_04925_));
 sky130_fd_sc_hd__and2_2 _11831_ (.A(_04772_),
    .B(_04767_),
    .X(_04926_));
 sky130_fd_sc_hd__nand2_1 _11832_ (.A(_04925_),
    .B(_04926_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand3b_2 _11833_ (.A_N(_04926_),
    .B(_04922_),
    .C(_04923_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _11834_ (.A(_04927_),
    .B(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _11835_ (.A(_04929_),
    .B(_04783_),
    .Y(_04930_));
 sky130_fd_sc_hd__inv_2 _11836_ (.A(_04783_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand3_1 _11837_ (.A(_04927_),
    .B(_04928_),
    .C(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__nand2_1 _11838_ (.A(_04930_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__inv_2 _11839_ (.A(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__nand2_1 _11840_ (.A(_04198_),
    .B(_04413_),
    .Y(_04936_));
 sky130_fd_sc_hd__nand2_1 _11841_ (.A(_04605_),
    .B(_04788_),
    .Y(_04937_));
 sky130_fd_sc_hd__nor2_1 _11842_ (.A(_04936_),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_1 _11843_ (.A(_04616_),
    .B(_04603_),
    .Y(_04939_));
 sky130_fd_sc_hd__nor2_1 _11844_ (.A(_04786_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__nand2_1 _11845_ (.A(_04610_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__a21boi_1 _11846_ (.A1(_04602_),
    .A2(_04785_),
    .B1_N(_04780_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_1 _11847_ (.A(_04941_),
    .B(_04942_),
    .Y(_04943_));
 sky130_fd_sc_hd__a21oi_2 _11848_ (.A1(_04204_),
    .A2(_04938_),
    .B1(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand2_1 _11849_ (.A(_04940_),
    .B(_04608_),
    .Y(_04945_));
 sky130_fd_sc_hd__nor2_1 _11850_ (.A(_04200_),
    .B(_04945_),
    .Y(_04947_));
 sky130_fd_sc_hd__nand3_2 _11851_ (.A(_04947_),
    .B(_01268_),
    .C(_02963_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_1 _11852_ (.A(_02968_),
    .B(_04947_),
    .Y(_04949_));
 sky130_fd_sc_hd__nand3_4 _11853_ (.A(_04944_),
    .B(_04948_),
    .C(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__or2_1 _11854_ (.A(_04934_),
    .B(_04950_),
    .X(_04951_));
 sky130_fd_sc_hd__nand2_1 _11855_ (.A(_04950_),
    .B(_04934_),
    .Y(_04952_));
 sky130_fd_sc_hd__and2_1 _11856_ (.A(_04951_),
    .B(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__clkbuf_1 _11857_ (.A(_04953_),
    .X(\m1.out[32] ));
 sky130_fd_sc_hd__nand2_1 _11858_ (.A(_04923_),
    .B(_04916_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _11859_ (.A(_04915_),
    .B(_04890_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _11860_ (.A(_04889_),
    .B(_04846_),
    .Y(_04957_));
 sky130_fd_sc_hd__nand2_1 _11861_ (.A(_04845_),
    .B(_04821_),
    .Y(_04958_));
 sky130_fd_sc_hd__inv_2 _11862_ (.A(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__nand2_1 _11863_ (.A(_04815_),
    .B(_04813_),
    .Y(_04960_));
 sky130_fd_sc_hd__inv_2 _11864_ (.A(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__inv_2 _11865_ (.A(net3),
    .Y(_04962_));
 sky130_fd_sc_hd__or3_2 _11866_ (.A(_04962_),
    .B(_00330_),
    .C(_04801_),
    .X(_04963_));
 sky130_fd_sc_hd__a21o_1 _11867_ (.A1(_06291_),
    .A2(_02423_),
    .B1(_06292_),
    .X(_04964_));
 sky130_fd_sc_hd__nand2_1 _11868_ (.A(_04963_),
    .B(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__nand2_1 _11869_ (.A(_06280_),
    .B(_02180_),
    .Y(_04966_));
 sky130_fd_sc_hd__nand2_1 _11870_ (.A(_04965_),
    .B(_04966_),
    .Y(_04968_));
 sky130_fd_sc_hd__inv_2 _11871_ (.A(_04966_),
    .Y(_04969_));
 sky130_fd_sc_hd__nand3_1 _11872_ (.A(_04963_),
    .B(_04969_),
    .C(_04964_),
    .Y(_04970_));
 sky130_fd_sc_hd__nand2_1 _11873_ (.A(_04968_),
    .B(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand2_1 _11874_ (.A(_04808_),
    .B(_04802_),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2b_2 _11875_ (.A_N(_04971_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__nand3_2 _11876_ (.A(_04971_),
    .B(_04802_),
    .C(_04808_),
    .Y(_04974_));
 sky130_fd_sc_hd__nand2_1 _11877_ (.A(_04973_),
    .B(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hd__nand2_1 _11878_ (.A(_06282_),
    .B(_06178_),
    .Y(_04976_));
 sky130_fd_sc_hd__and4_1 _11879_ (.A(_06279_),
    .B(_06284_),
    .C(_06176_),
    .D(_01922_),
    .X(_04977_));
 sky130_fd_sc_hd__a22o_1 _11880_ (.A1(_06279_),
    .A2(_01921_),
    .B1(_06284_),
    .B2(_01692_),
    .X(_04979_));
 sky130_fd_sc_hd__inv_2 _11881_ (.A(_04979_),
    .Y(_04980_));
 sky130_fd_sc_hd__nor2_1 _11882_ (.A(_04977_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__xor2_1 _11883_ (.A(_04976_),
    .B(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__nand2_1 _11884_ (.A(_04975_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__inv_2 _11885_ (.A(_04982_),
    .Y(_04984_));
 sky130_fd_sc_hd__nand3_2 _11886_ (.A(_04973_),
    .B(_04984_),
    .C(_04974_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_1 _11887_ (.A(_04983_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_1 _11888_ (.A(_04961_),
    .B(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand3_2 _11889_ (.A(_04960_),
    .B(_04983_),
    .C(_04985_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand2_1 _11890_ (.A(_04987_),
    .B(_04988_),
    .Y(_04990_));
 sky130_fd_sc_hd__inv_2 _11891_ (.A(_04794_),
    .Y(_04991_));
 sky130_fd_sc_hd__a21oi_1 _11892_ (.A1(_04796_),
    .A2(_04991_),
    .B1(_04795_),
    .Y(_04992_));
 sky130_fd_sc_hd__nand2_1 _11893_ (.A(_06243_),
    .B(_06222_),
    .Y(_04993_));
 sky130_fd_sc_hd__inv_2 _11894_ (.A(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nand2_1 _11895_ (.A(_06235_),
    .B(_06174_),
    .Y(_04995_));
 sky130_fd_sc_hd__nand2_1 _11896_ (.A(_06238_),
    .B(_06172_),
    .Y(_04996_));
 sky130_fd_sc_hd__xor2_1 _11897_ (.A(_04995_),
    .B(_04996_),
    .X(_04997_));
 sky130_fd_sc_hd__or2_1 _11898_ (.A(_04994_),
    .B(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__nand2_1 _11899_ (.A(_04997_),
    .B(_04994_),
    .Y(_04999_));
 sky130_fd_sc_hd__nand2_1 _11900_ (.A(_04998_),
    .B(_04999_),
    .Y(_05001_));
 sky130_fd_sc_hd__or2_1 _11901_ (.A(_04992_),
    .B(_05001_),
    .X(_05002_));
 sky130_fd_sc_hd__nand2_1 _11902_ (.A(_05001_),
    .B(_04992_),
    .Y(_05003_));
 sky130_fd_sc_hd__nand2_1 _11903_ (.A(_05002_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__inv_2 _11904_ (.A(_04832_),
    .Y(_05005_));
 sky130_fd_sc_hd__nor2_1 _11905_ (.A(_04824_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__nand2_1 _11906_ (.A(_05004_),
    .B(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__inv_2 _11907_ (.A(_05006_),
    .Y(_05008_));
 sky130_fd_sc_hd__nand3_1 _11908_ (.A(_05008_),
    .B(_05002_),
    .C(_05003_),
    .Y(_05009_));
 sky130_fd_sc_hd__nand2_1 _11909_ (.A(_05007_),
    .B(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__nand2_1 _11910_ (.A(_04990_),
    .B(_05010_),
    .Y(_05012_));
 sky130_fd_sc_hd__inv_2 _11911_ (.A(_05010_),
    .Y(_05013_));
 sky130_fd_sc_hd__nand3_2 _11912_ (.A(_04987_),
    .B(_04988_),
    .C(_05013_),
    .Y(_05014_));
 sky130_fd_sc_hd__nand2_1 _11913_ (.A(_05012_),
    .B(_05014_),
    .Y(_05015_));
 sky130_fd_sc_hd__nand2_1 _11914_ (.A(_04959_),
    .B(_05015_),
    .Y(_05016_));
 sky130_fd_sc_hd__nand3_2 _11915_ (.A(_04958_),
    .B(_05012_),
    .C(_05014_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _11916_ (.A(_05016_),
    .B(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__nand2_1 _11917_ (.A(_06247_),
    .B(_06221_),
    .Y(_05019_));
 sky130_fd_sc_hd__inv_2 _11918_ (.A(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__nand2_1 _11919_ (.A(_06248_),
    .B(_06218_),
    .Y(_05021_));
 sky130_fd_sc_hd__nor3_1 _11920_ (.A(_04495_),
    .B(_04854_),
    .C(_05021_),
    .Y(_05023_));
 sky130_fd_sc_hd__inv_2 _11921_ (.A(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hd__o21ai_1 _11922_ (.A1(_04495_),
    .A2(_04854_),
    .B1(_05021_),
    .Y(_05025_));
 sky130_fd_sc_hd__and2_1 _11923_ (.A(_05024_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__or2_1 _11924_ (.A(_05020_),
    .B(_05026_),
    .X(_05027_));
 sky130_fd_sc_hd__nand2_1 _11925_ (.A(_05026_),
    .B(_05020_),
    .Y(_05028_));
 sky130_fd_sc_hd__nand2_1 _11926_ (.A(_05027_),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__nand3_1 _11927_ (.A(_05029_),
    .B(_04857_),
    .C(_04861_),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_1 _11928_ (.A(_04861_),
    .B(_04857_),
    .Y(_05031_));
 sky130_fd_sc_hd__nand3_1 _11929_ (.A(_05031_),
    .B(_05027_),
    .C(_05028_),
    .Y(_05032_));
 sky130_fd_sc_hd__nand2_1 _11930_ (.A(_05030_),
    .B(_05032_),
    .Y(_05034_));
 sky130_fd_sc_hd__or3b_1 _11931_ (.A(_06250_),
    .B(_04496_),
    .C_N(_06231_),
    .X(_05035_));
 sky130_fd_sc_hd__a21o_1 _11932_ (.A1(_06299_),
    .A2(_06228_),
    .B1(_06231_),
    .X(_05036_));
 sky130_fd_sc_hd__nand2_1 _11933_ (.A(_05035_),
    .B(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _11934_ (.A(_05034_),
    .B(_05037_),
    .Y(_05038_));
 sky130_fd_sc_hd__inv_2 _11935_ (.A(_05037_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand3_1 _11936_ (.A(_05030_),
    .B(_05032_),
    .C(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_1 _11937_ (.A(_05038_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__a21oi_2 _11938_ (.A1(_04840_),
    .A2(_04823_),
    .B1(_04839_),
    .Y(_05042_));
 sky130_fd_sc_hd__inv_2 _11939_ (.A(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_1 _11940_ (.A(_05041_),
    .B(_05043_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand3_1 _11941_ (.A(_05038_),
    .B(_05042_),
    .C(_05040_),
    .Y(_05046_));
 sky130_fd_sc_hd__nand2_1 _11942_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hd__a21o_1 _11943_ (.A1(_04870_),
    .A2(_04871_),
    .B1(_04864_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_1 _11944_ (.A(_05047_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__nand3b_1 _11945_ (.A_N(_05048_),
    .B(_05045_),
    .C(_05046_),
    .Y(_05050_));
 sky130_fd_sc_hd__nand2_1 _11946_ (.A(_05049_),
    .B(_05050_),
    .Y(_05051_));
 sky130_fd_sc_hd__nand2_1 _11947_ (.A(_05018_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__inv_2 _11948_ (.A(_05051_),
    .Y(_05053_));
 sky130_fd_sc_hd__nand3_1 _11949_ (.A(_05016_),
    .B(_05017_),
    .C(_05053_),
    .Y(_05054_));
 sky130_fd_sc_hd__nand3_2 _11950_ (.A(_04957_),
    .B(_05052_),
    .C(_05054_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_1 _11951_ (.A(_05052_),
    .B(_05054_),
    .Y(_05057_));
 sky130_fd_sc_hd__a21boi_1 _11952_ (.A1(_04888_),
    .A2(_04849_),
    .B1_N(_04846_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand2_1 _11953_ (.A(_05057_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _11954_ (.A(_05056_),
    .B(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__a21oi_1 _11955_ (.A1(_04866_),
    .A2(_06225_),
    .B1(_04865_),
    .Y(_05061_));
 sky130_fd_sc_hd__nand2_1 _11956_ (.A(_04876_),
    .B(_04879_),
    .Y(_05062_));
 sky130_fd_sc_hd__nor2_1 _11957_ (.A(_04879_),
    .B(_04876_),
    .Y(_05063_));
 sky130_fd_sc_hd__a21oi_1 _11958_ (.A1(_05062_),
    .A2(_04883_),
    .B1(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__nor2_1 _11959_ (.A(_05061_),
    .B(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__inv_2 _11960_ (.A(_05065_),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_1 _11961_ (.A(_05064_),
    .B(_05061_),
    .Y(_05068_));
 sky130_fd_sc_hd__nand2_1 _11962_ (.A(_05067_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__nand2_1 _11963_ (.A(_05069_),
    .B(_04898_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand3_1 _11964_ (.A(_05067_),
    .B(_04897_),
    .C(_05068_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _11965_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(_05060_),
    .B(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__inv_2 _11967_ (.A(_05072_),
    .Y(_05074_));
 sky130_fd_sc_hd__nand3_1 _11968_ (.A(_05056_),
    .B(_05059_),
    .C(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__nand3_1 _11969_ (.A(_04955_),
    .B(_05073_),
    .C(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hd__nand2_1 _11970_ (.A(_05073_),
    .B(_05075_),
    .Y(_05078_));
 sky130_fd_sc_hd__a21boi_1 _11971_ (.A1(_04914_),
    .A2(_04893_),
    .B1_N(_04890_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2_1 _11972_ (.A(_05078_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand2_1 _11973_ (.A(_05076_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__nand2_1 _11974_ (.A(_04910_),
    .B(_04905_),
    .Y(_05082_));
 sky130_fd_sc_hd__inv_2 _11975_ (.A(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _11976_ (.A(_05081_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__nand3_1 _11977_ (.A(_05076_),
    .B(_05080_),
    .C(_05082_),
    .Y(_05085_));
 sky130_fd_sc_hd__nand3_1 _11978_ (.A(_04954_),
    .B(_05084_),
    .C(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__inv_2 _11979_ (.A(_04928_),
    .Y(_05087_));
 sky130_fd_sc_hd__nand2_1 _11980_ (.A(_05084_),
    .B(_05085_),
    .Y(_05089_));
 sky130_fd_sc_hd__a21boi_1 _11981_ (.A1(_04920_),
    .A2(_04918_),
    .B1_N(_04916_),
    .Y(_05090_));
 sky130_fd_sc_hd__nand2_1 _11982_ (.A(_05089_),
    .B(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__nand3_1 _11983_ (.A(_05086_),
    .B(_05087_),
    .C(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__nand2_1 _11984_ (.A(_05086_),
    .B(_05091_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _11985_ (.A(_05093_),
    .B(_04928_),
    .Y(_05094_));
 sky130_fd_sc_hd__nand2_1 _11986_ (.A(_05092_),
    .B(_05094_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _11987_ (.A(_04952_),
    .B(_04932_),
    .Y(_05096_));
 sky130_fd_sc_hd__xnor2_1 _11988_ (.A(_05095_),
    .B(_05096_),
    .Y(\m1.out[33] ));
 sky130_fd_sc_hd__nand2_1 _11989_ (.A(_05085_),
    .B(_05076_),
    .Y(_05097_));
 sky130_fd_sc_hd__nand2_1 _11990_ (.A(_05075_),
    .B(_05056_),
    .Y(_05099_));
 sky130_fd_sc_hd__nand2_1 _11991_ (.A(_05054_),
    .B(_05017_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _11992_ (.A(_05014_),
    .B(_04988_),
    .Y(_05101_));
 sky130_fd_sc_hd__nand2_1 _11993_ (.A(_04985_),
    .B(_04973_),
    .Y(_05102_));
 sky130_fd_sc_hd__or3_1 _11994_ (.A(_04962_),
    .B(_00700_),
    .C(_04801_),
    .X(_05103_));
 sky130_fd_sc_hd__a21o_1 _11995_ (.A1(_06280_),
    .A2(_02423_),
    .B1(_06291_),
    .X(_05104_));
 sky130_fd_sc_hd__nand2_1 _11996_ (.A(_05103_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__nand2_1 _11997_ (.A(_06279_),
    .B(_02181_),
    .Y(_05106_));
 sky130_fd_sc_hd__nand2_1 _11998_ (.A(_05105_),
    .B(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__nand3b_1 _11999_ (.A_N(_05106_),
    .B(_05103_),
    .C(_05104_),
    .Y(_05108_));
 sky130_fd_sc_hd__nand2_1 _12000_ (.A(_05107_),
    .B(_05108_),
    .Y(_05110_));
 sky130_fd_sc_hd__nand2_1 _12001_ (.A(_04970_),
    .B(_04963_),
    .Y(_05111_));
 sky130_fd_sc_hd__nand2b_1 _12002_ (.A_N(_05110_),
    .B(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__nand3_1 _12003_ (.A(_05110_),
    .B(_04963_),
    .C(_04970_),
    .Y(_05113_));
 sky130_fd_sc_hd__nand2_1 _12004_ (.A(_05112_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__and4_1 _12005_ (.A(_01831_),
    .B(_01158_),
    .C(_06175_),
    .D(_06187_),
    .X(_05115_));
 sky130_fd_sc_hd__a22o_1 _12006_ (.A1(_01831_),
    .A2(_06175_),
    .B1(_01158_),
    .B2(_06187_),
    .X(_05116_));
 sky130_fd_sc_hd__nand2b_1 _12007_ (.A_N(_05115_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _12008_ (.A(_06238_),
    .B(_06178_),
    .Y(_05118_));
 sky130_fd_sc_hd__nand2_1 _12009_ (.A(_05117_),
    .B(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hd__inv_2 _12010_ (.A(_05118_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand3b_1 _12011_ (.A_N(_05115_),
    .B(_05121_),
    .C(_05116_),
    .Y(_05122_));
 sky130_fd_sc_hd__nand2_1 _12012_ (.A(_05119_),
    .B(_05122_),
    .Y(_05123_));
 sky130_fd_sc_hd__nand2_1 _12013_ (.A(_05114_),
    .B(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__inv_2 _12014_ (.A(_05123_),
    .Y(_05125_));
 sky130_fd_sc_hd__nand3_1 _12015_ (.A(_05112_),
    .B(_05125_),
    .C(_05113_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand3_1 _12016_ (.A(_05102_),
    .B(_05124_),
    .C(_05126_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _12017_ (.A(_05124_),
    .B(_05126_),
    .Y(_05128_));
 sky130_fd_sc_hd__a21boi_1 _12018_ (.A1(_04984_),
    .A2(_04974_),
    .B1_N(_04973_),
    .Y(_05129_));
 sky130_fd_sc_hd__nand2_1 _12019_ (.A(_05128_),
    .B(_05129_),
    .Y(_05130_));
 sky130_fd_sc_hd__nand2_1 _12020_ (.A(_05127_),
    .B(_05130_),
    .Y(_05132_));
 sky130_fd_sc_hd__inv_2 _12021_ (.A(_04976_),
    .Y(_05133_));
 sky130_fd_sc_hd__a21oi_1 _12022_ (.A1(_04979_),
    .A2(_05133_),
    .B1(_04977_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_1 _12023_ (.A(_01858_),
    .B(_00918_),
    .Y(_05135_));
 sky130_fd_sc_hd__inv_2 _12024_ (.A(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__nand2_1 _12025_ (.A(_06241_),
    .B(_01278_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand2_1 _12026_ (.A(_06235_),
    .B(_06171_),
    .Y(_05138_));
 sky130_fd_sc_hd__xor2_1 _12027_ (.A(_05137_),
    .B(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__or2_1 _12028_ (.A(_05136_),
    .B(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__nand2_1 _12029_ (.A(_05139_),
    .B(_05136_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2_1 _12030_ (.A(_05140_),
    .B(_05141_),
    .Y(_05143_));
 sky130_fd_sc_hd__or2_1 _12031_ (.A(_05134_),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__nand2_1 _12032_ (.A(_05143_),
    .B(_05134_),
    .Y(_05145_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_05144_),
    .B(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hd__and4_1 _12034_ (.A(_06236_),
    .B(_06238_),
    .C(_06172_),
    .D(_06174_),
    .X(_05147_));
 sky130_fd_sc_hd__inv_2 _12035_ (.A(_04999_),
    .Y(_05148_));
 sky130_fd_sc_hd__nor2_1 _12036_ (.A(_05147_),
    .B(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__nand2_1 _12037_ (.A(_05146_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__nand3b_1 _12038_ (.A_N(_05149_),
    .B(_05144_),
    .C(_05145_),
    .Y(_05151_));
 sky130_fd_sc_hd__nand2_1 _12039_ (.A(_05150_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__nand2_1 _12040_ (.A(_05132_),
    .B(_05152_),
    .Y(_05154_));
 sky130_fd_sc_hd__inv_2 _12041_ (.A(_05152_),
    .Y(_05155_));
 sky130_fd_sc_hd__nand3_1 _12042_ (.A(_05127_),
    .B(_05130_),
    .C(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__nand3_2 _12043_ (.A(_05101_),
    .B(_05154_),
    .C(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2_1 _12044_ (.A(_05154_),
    .B(_05156_),
    .Y(_05158_));
 sky130_fd_sc_hd__a21boi_1 _12045_ (.A1(_04987_),
    .A2(_05013_),
    .B1_N(_04988_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2_1 _12046_ (.A(_05158_),
    .B(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__nand2_1 _12047_ (.A(_05157_),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__nand2_1 _12048_ (.A(_06247_),
    .B(_06218_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(_06248_),
    .B(_06223_),
    .Y(_05163_));
 sky130_fd_sc_hd__xor2_1 _12050_ (.A(_05162_),
    .B(_05163_),
    .X(_05165_));
 sky130_fd_sc_hd__nand2_1 _12051_ (.A(_03905_),
    .B(_06221_),
    .Y(_05166_));
 sky130_fd_sc_hd__inv_2 _12052_ (.A(_05166_),
    .Y(_05167_));
 sky130_fd_sc_hd__nand2_1 _12053_ (.A(_05165_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__or2_1 _12054_ (.A(_05167_),
    .B(_05165_),
    .X(_05169_));
 sky130_fd_sc_hd__nand2_1 _12055_ (.A(_05028_),
    .B(_05024_),
    .Y(_05170_));
 sky130_fd_sc_hd__a21o_1 _12056_ (.A1(_05168_),
    .A2(_05169_),
    .B1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nand3_1 _12057_ (.A(_05170_),
    .B(_05168_),
    .C(_05169_),
    .Y(_05172_));
 sky130_fd_sc_hd__nand2_1 _12058_ (.A(_05171_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__nand2_1 _12059_ (.A(_05173_),
    .B(_04496_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand3_1 _12060_ (.A(_05171_),
    .B(_06228_),
    .C(_05172_),
    .Y(_05176_));
 sky130_fd_sc_hd__nand2_1 _12061_ (.A(_05174_),
    .B(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__nand2_1 _12062_ (.A(_05009_),
    .B(_05002_),
    .Y(_05178_));
 sky130_fd_sc_hd__inv_2 _12063_ (.A(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand2_1 _12064_ (.A(_05177_),
    .B(_05179_),
    .Y(_05180_));
 sky130_fd_sc_hd__nand3_1 _12065_ (.A(_05178_),
    .B(_05174_),
    .C(_05176_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _12066_ (.A(_05180_),
    .B(_05181_),
    .Y(_05182_));
 sky130_fd_sc_hd__nand2_1 _12067_ (.A(_05040_),
    .B(_05032_),
    .Y(_05183_));
 sky130_fd_sc_hd__inv_2 _12068_ (.A(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__nand2_1 _12069_ (.A(_05182_),
    .B(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__nand3_1 _12070_ (.A(_05180_),
    .B(_05181_),
    .C(_05183_),
    .Y(_05187_));
 sky130_fd_sc_hd__nand2_1 _12071_ (.A(_05185_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand2_1 _12072_ (.A(_05161_),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__inv_2 _12073_ (.A(_05188_),
    .Y(_05190_));
 sky130_fd_sc_hd__nand3_1 _12074_ (.A(_05157_),
    .B(_05160_),
    .C(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__nand3_2 _12075_ (.A(_05100_),
    .B(_05189_),
    .C(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__nand2_1 _12076_ (.A(_05189_),
    .B(_05191_),
    .Y(_05193_));
 sky130_fd_sc_hd__a21boi_1 _12077_ (.A1(_05016_),
    .A2(_05053_),
    .B1_N(_05017_),
    .Y(_05194_));
 sky130_fd_sc_hd__nand2_1 _12078_ (.A(_05193_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__nand2_1 _12079_ (.A(_05192_),
    .B(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__o21a_1 _12080_ (.A1(_05041_),
    .A2(_05042_),
    .B1(_05049_),
    .X(_05198_));
 sky130_fd_sc_hd__nor2_1 _12081_ (.A(_05035_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__inv_2 _12082_ (.A(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__nand2_1 _12083_ (.A(_05198_),
    .B(_05035_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(_05200_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__nand2_1 _12085_ (.A(_05196_),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__inv_2 _12086_ (.A(_05202_),
    .Y(_05204_));
 sky130_fd_sc_hd__nand3_1 _12087_ (.A(_05192_),
    .B(_05195_),
    .C(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hd__nand3_1 _12088_ (.A(_05099_),
    .B(_05203_),
    .C(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_1 _12089_ (.A(_05203_),
    .B(_05205_),
    .Y(_05207_));
 sky130_fd_sc_hd__a21boi_1 _12090_ (.A1(_05074_),
    .A2(_05059_),
    .B1_N(_05056_),
    .Y(_05209_));
 sky130_fd_sc_hd__nand2_1 _12091_ (.A(_05207_),
    .B(_05209_),
    .Y(_05210_));
 sky130_fd_sc_hd__nand2_1 _12092_ (.A(_05206_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__nand2_2 _12093_ (.A(_05071_),
    .B(_05067_),
    .Y(_05212_));
 sky130_fd_sc_hd__inv_2 _12094_ (.A(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__nand2_1 _12095_ (.A(_05211_),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__nand3_1 _12096_ (.A(_05206_),
    .B(_05210_),
    .C(_05212_),
    .Y(_05215_));
 sky130_fd_sc_hd__nand3_2 _12097_ (.A(_05097_),
    .B(_05214_),
    .C(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_1 _12098_ (.A(_05214_),
    .B(_05215_),
    .Y(_05217_));
 sky130_fd_sc_hd__a21boi_1 _12099_ (.A1(_05082_),
    .A2(_05080_),
    .B1_N(_05076_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand2_1 _12100_ (.A(_05217_),
    .B(_05218_),
    .Y(_05220_));
 sky130_fd_sc_hd__nand2_1 _12101_ (.A(_05216_),
    .B(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__nand2_1 _12102_ (.A(_05221_),
    .B(_05086_),
    .Y(_05222_));
 sky130_fd_sc_hd__nor2_1 _12103_ (.A(_05090_),
    .B(_05089_),
    .Y(_05223_));
 sky130_fd_sc_hd__nand3_2 _12104_ (.A(_05216_),
    .B(_05223_),
    .C(_05220_),
    .Y(_05224_));
 sky130_fd_sc_hd__nand2_1 _12105_ (.A(_05222_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__inv_2 _12106_ (.A(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__nor2_1 _12107_ (.A(_04933_),
    .B(_05095_),
    .Y(_05227_));
 sky130_fd_sc_hd__inv_2 _12108_ (.A(_05094_),
    .Y(_05228_));
 sky130_fd_sc_hd__o21ai_1 _12109_ (.A1(_04932_),
    .A2(_05228_),
    .B1(_05092_),
    .Y(_05229_));
 sky130_fd_sc_hd__a21o_1 _12110_ (.A1(_04950_),
    .A2(_05227_),
    .B1(_05229_),
    .X(_05231_));
 sky130_fd_sc_hd__or2_1 _12111_ (.A(_05226_),
    .B(_05231_),
    .X(_05232_));
 sky130_fd_sc_hd__nand2_1 _12112_ (.A(_05231_),
    .B(_05226_),
    .Y(_05233_));
 sky130_fd_sc_hd__and2_1 _12113_ (.A(_05232_),
    .B(_05233_),
    .X(_05234_));
 sky130_fd_sc_hd__clkbuf_1 _12114_ (.A(_05234_),
    .X(\m1.out[34] ));
 sky130_fd_sc_hd__nand2_1 _12115_ (.A(_05215_),
    .B(_05206_),
    .Y(_05235_));
 sky130_fd_sc_hd__nand2_1 _12116_ (.A(_05205_),
    .B(_05192_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_1 _12117_ (.A(_05191_),
    .B(_05157_),
    .Y(_05237_));
 sky130_fd_sc_hd__inv_2 _12118_ (.A(_06278_),
    .Y(_05238_));
 sky130_fd_sc_hd__or3_1 _12119_ (.A(_05238_),
    .B(_00700_),
    .C(_04801_),
    .X(_05239_));
 sky130_fd_sc_hd__a21o_1 _12120_ (.A1(_00701_),
    .A2(_06183_),
    .B1(_00849_),
    .X(_05241_));
 sky130_fd_sc_hd__nand2_1 _12121_ (.A(_05239_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__nand2_1 _12122_ (.A(_06283_),
    .B(_02180_),
    .Y(_05243_));
 sky130_fd_sc_hd__nand2_1 _12123_ (.A(_05242_),
    .B(_05243_),
    .Y(_05244_));
 sky130_fd_sc_hd__inv_2 _12124_ (.A(_05243_),
    .Y(_05245_));
 sky130_fd_sc_hd__nand3_1 _12125_ (.A(_05239_),
    .B(_05245_),
    .C(_05241_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand2_1 _12126_ (.A(_05244_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__and2_1 _12127_ (.A(_05108_),
    .B(_05103_),
    .X(_05248_));
 sky130_fd_sc_hd__nor2_1 _12128_ (.A(_05247_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__inv_2 _12129_ (.A(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__nand2_1 _12130_ (.A(_05248_),
    .B(_05247_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_1 _12131_ (.A(_05250_),
    .B(_05252_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand2_1 _12132_ (.A(_06236_),
    .B(_06179_),
    .Y(_05254_));
 sky130_fd_sc_hd__nand2_1 _12133_ (.A(_06238_),
    .B(_06176_),
    .Y(_05255_));
 sky130_fd_sc_hd__nor3_1 _12134_ (.A(_01422_),
    .B(_06188_),
    .C(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__o21ai_1 _12135_ (.A1(_01422_),
    .A2(_06188_),
    .B1(_05255_),
    .Y(_05257_));
 sky130_fd_sc_hd__and2b_1 _12136_ (.A_N(_05256_),
    .B(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__xor2_1 _12137_ (.A(_05254_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__nand2_1 _12138_ (.A(_05253_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand3b_1 _12139_ (.A_N(_05259_),
    .B(_05250_),
    .C(_05252_),
    .Y(_05261_));
 sky130_fd_sc_hd__nand2_1 _12140_ (.A(_05260_),
    .B(_05261_),
    .Y(_05263_));
 sky130_fd_sc_hd__nand2_1 _12141_ (.A(_05126_),
    .B(_05112_),
    .Y(_05264_));
 sky130_fd_sc_hd__inv_2 _12142_ (.A(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand2_1 _12143_ (.A(_05263_),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__nand3_1 _12144_ (.A(_05264_),
    .B(_05260_),
    .C(_05261_),
    .Y(_05267_));
 sky130_fd_sc_hd__nand2_1 _12145_ (.A(_05266_),
    .B(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hd__a21oi_1 _12146_ (.A1(_05116_),
    .A2(_05121_),
    .B1(_05115_),
    .Y(_05269_));
 sky130_fd_sc_hd__nand2_1 _12147_ (.A(_02095_),
    .B(_00918_),
    .Y(_05270_));
 sky130_fd_sc_hd__inv_2 _12148_ (.A(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__nand2_1 _12149_ (.A(_01858_),
    .B(_01278_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand2_1 _12150_ (.A(_06242_),
    .B(_06171_),
    .Y(_05274_));
 sky130_fd_sc_hd__xor2_1 _12151_ (.A(_05272_),
    .B(_05274_),
    .X(_05275_));
 sky130_fd_sc_hd__or2_1 _12152_ (.A(_05271_),
    .B(_05275_),
    .X(_05276_));
 sky130_fd_sc_hd__nand2_1 _12153_ (.A(_05275_),
    .B(_05271_),
    .Y(_05277_));
 sky130_fd_sc_hd__nand2_1 _12154_ (.A(_05276_),
    .B(_05277_),
    .Y(_05278_));
 sky130_fd_sc_hd__or2_1 _12155_ (.A(_05269_),
    .B(_05278_),
    .X(_05279_));
 sky130_fd_sc_hd__nand2_1 _12156_ (.A(_05278_),
    .B(_05269_),
    .Y(_05280_));
 sky130_fd_sc_hd__and4_1 _12157_ (.A(_06236_),
    .B(_06243_),
    .C(_06172_),
    .D(_06174_),
    .X(_05281_));
 sky130_fd_sc_hd__inv_2 _12158_ (.A(_05141_),
    .Y(_05282_));
 sky130_fd_sc_hd__nor2_1 _12159_ (.A(_05281_),
    .B(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__inv_2 _12160_ (.A(_05283_),
    .Y(_05285_));
 sky130_fd_sc_hd__a21o_1 _12161_ (.A1(_05279_),
    .A2(_05280_),
    .B1(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__nand3_1 _12162_ (.A(_05279_),
    .B(_05285_),
    .C(_05280_),
    .Y(_05287_));
 sky130_fd_sc_hd__nand2_1 _12163_ (.A(_05286_),
    .B(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__nand2_1 _12164_ (.A(_05268_),
    .B(_05288_),
    .Y(_05289_));
 sky130_fd_sc_hd__inv_2 _12165_ (.A(_05288_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand3_1 _12166_ (.A(_05266_),
    .B(_05267_),
    .C(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__nand2_1 _12167_ (.A(_05289_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nand2_1 _12168_ (.A(_05156_),
    .B(_05127_),
    .Y(_05293_));
 sky130_fd_sc_hd__inv_2 _12169_ (.A(_05293_),
    .Y(_05294_));
 sky130_fd_sc_hd__nand2_1 _12170_ (.A(_05292_),
    .B(_05294_),
    .Y(_05296_));
 sky130_fd_sc_hd__nand3_1 _12171_ (.A(_05293_),
    .B(_05289_),
    .C(_05291_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand2_1 _12172_ (.A(_05296_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__o21a_1 _12173_ (.A1(_05162_),
    .A2(_05163_),
    .B1(_05168_),
    .X(_05299_));
 sky130_fd_sc_hd__and4_1 _12174_ (.A(_06246_),
    .B(_06298_),
    .C(_06218_),
    .D(_06223_),
    .X(_05300_));
 sky130_fd_sc_hd__a22o_1 _12175_ (.A1(_06246_),
    .A2(_06223_),
    .B1(_03905_),
    .B2(_06218_),
    .X(_05301_));
 sky130_fd_sc_hd__and2b_1 _12176_ (.A_N(_05300_),
    .B(_05301_),
    .X(_05302_));
 sky130_fd_sc_hd__or2_1 _12177_ (.A(_06221_),
    .B(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__nand2_1 _12178_ (.A(_05302_),
    .B(_06221_),
    .Y(_05304_));
 sky130_fd_sc_hd__nand2_1 _12179_ (.A(_05303_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__or2_1 _12180_ (.A(_05299_),
    .B(_05305_),
    .X(_05307_));
 sky130_fd_sc_hd__nand2_1 _12181_ (.A(_05305_),
    .B(_05299_),
    .Y(_05308_));
 sky130_fd_sc_hd__nand2_1 _12182_ (.A(_05307_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__nand3_1 _12183_ (.A(_05309_),
    .B(_05144_),
    .C(_05151_),
    .Y(_05310_));
 sky130_fd_sc_hd__nand2_1 _12184_ (.A(_05151_),
    .B(_05144_),
    .Y(_05311_));
 sky130_fd_sc_hd__nand3_1 _12185_ (.A(_05311_),
    .B(_05308_),
    .C(_05307_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2_1 _12186_ (.A(_05310_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__nand2_1 _12187_ (.A(_05176_),
    .B(_05172_),
    .Y(_05314_));
 sky130_fd_sc_hd__inv_2 _12188_ (.A(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_1 _12189_ (.A(_05313_),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__nand3_1 _12190_ (.A(_05310_),
    .B(_05314_),
    .C(_05312_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand2_1 _12191_ (.A(_05316_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__nand2_1 _12192_ (.A(_05298_),
    .B(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__inv_2 _12193_ (.A(_05319_),
    .Y(_05321_));
 sky130_fd_sc_hd__nand3_1 _12194_ (.A(_05296_),
    .B(_05297_),
    .C(_05321_),
    .Y(_05322_));
 sky130_fd_sc_hd__nand3_1 _12195_ (.A(_05237_),
    .B(_05320_),
    .C(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__nand2_1 _12196_ (.A(_05320_),
    .B(_05322_),
    .Y(_05324_));
 sky130_fd_sc_hd__a21boi_1 _12197_ (.A1(_05190_),
    .A2(_05160_),
    .B1_N(_05157_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_1 _12198_ (.A(_05324_),
    .B(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__nand2_1 _12199_ (.A(_05323_),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__nand2_1 _12200_ (.A(_05187_),
    .B(_05181_),
    .Y(_05329_));
 sky130_fd_sc_hd__inv_2 _12201_ (.A(_05329_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _12202_ (.A(_05327_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__nand3_1 _12203_ (.A(_05323_),
    .B(_05326_),
    .C(_05329_),
    .Y(_05332_));
 sky130_fd_sc_hd__nand3_1 _12204_ (.A(_05236_),
    .B(_05331_),
    .C(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(_05331_),
    .B(_05332_),
    .Y(_05334_));
 sky130_fd_sc_hd__a21boi_1 _12206_ (.A1(_05204_),
    .A2(_05195_),
    .B1_N(_05192_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand2_1 _12207_ (.A(_05334_),
    .B(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__nand3_1 _12208_ (.A(_05333_),
    .B(_05336_),
    .C(_05199_),
    .Y(_05337_));
 sky130_fd_sc_hd__nand2_1 _12209_ (.A(_05333_),
    .B(_05336_),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _12210_ (.A(_05338_),
    .B(_05200_),
    .Y(_05340_));
 sky130_fd_sc_hd__nand3_1 _12211_ (.A(_05235_),
    .B(_05337_),
    .C(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__nand2_1 _12212_ (.A(_05340_),
    .B(_05337_),
    .Y(_05342_));
 sky130_fd_sc_hd__a21boi_1 _12213_ (.A1(_05212_),
    .A2(_05210_),
    .B1_N(_05206_),
    .Y(_05343_));
 sky130_fd_sc_hd__nand2_1 _12214_ (.A(_05342_),
    .B(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(_05341_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_1 _12216_ (.A(_05345_),
    .B(_05216_),
    .Y(_05346_));
 sky130_fd_sc_hd__nor2_1 _12217_ (.A(_05218_),
    .B(_05217_),
    .Y(_05347_));
 sky130_fd_sc_hd__nand3_1 _12218_ (.A(_05341_),
    .B(_05347_),
    .C(_05344_),
    .Y(_05348_));
 sky130_fd_sc_hd__nand2_1 _12219_ (.A(_05346_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _12220_ (.A(_05233_),
    .B(_05224_),
    .Y(_05351_));
 sky130_fd_sc_hd__xnor2_1 _12221_ (.A(_05349_),
    .B(_05351_),
    .Y(\m1.out[35] ));
 sky130_fd_sc_hd__nand2_1 _12222_ (.A(_05337_),
    .B(_05333_),
    .Y(_05352_));
 sky130_fd_sc_hd__and2_1 _12223_ (.A(_05332_),
    .B(_05323_),
    .X(_05353_));
 sky130_fd_sc_hd__nand2_1 _12224_ (.A(_05261_),
    .B(_05250_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand2_2 _12225_ (.A(_06241_),
    .B(_06177_),
    .Y(_05355_));
 sky130_fd_sc_hd__inv_2 _12226_ (.A(_06237_),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_1 _12227_ (.A(_06234_),
    .B(_06175_),
    .Y(_05357_));
 sky130_fd_sc_hd__nor3_1 _12228_ (.A(_05356_),
    .B(_06188_),
    .C(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hd__o21ai_1 _12229_ (.A1(_05356_),
    .A2(_06188_),
    .B1(_05357_),
    .Y(_05359_));
 sky130_fd_sc_hd__and2b_1 _12230_ (.A_N(_05358_),
    .B(_05359_),
    .X(_05361_));
 sky130_fd_sc_hd__xor2_1 _12231_ (.A(_05355_),
    .B(_05361_),
    .X(_05362_));
 sky130_fd_sc_hd__inv_2 _12232_ (.A(_06283_),
    .Y(_05363_));
 sky130_fd_sc_hd__or3_1 _12233_ (.A(_05238_),
    .B(_05363_),
    .C(_04801_),
    .X(_05364_));
 sky130_fd_sc_hd__a21o_1 _12234_ (.A1(_01158_),
    .A2(_06183_),
    .B1(_06279_),
    .X(_05365_));
 sky130_fd_sc_hd__nand2_1 _12235_ (.A(_05364_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _12236_ (.A(_01831_),
    .B(_02180_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _12237_ (.A(_05366_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__inv_2 _12238_ (.A(_05367_),
    .Y(_05369_));
 sky130_fd_sc_hd__nand3_1 _12239_ (.A(_05364_),
    .B(_05369_),
    .C(_05365_),
    .Y(_05370_));
 sky130_fd_sc_hd__nand2_1 _12240_ (.A(_05368_),
    .B(_05370_),
    .Y(_05372_));
 sky130_fd_sc_hd__and2_1 _12241_ (.A(_05246_),
    .B(_05239_),
    .X(_05373_));
 sky130_fd_sc_hd__or2_1 _12242_ (.A(_05372_),
    .B(_05373_),
    .X(_05374_));
 sky130_fd_sc_hd__nand2_1 _12243_ (.A(_05373_),
    .B(_05372_),
    .Y(_05375_));
 sky130_fd_sc_hd__nand3b_2 _12244_ (.A_N(_05362_),
    .B(_05374_),
    .C(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand2_1 _12245_ (.A(_05374_),
    .B(_05375_),
    .Y(_05377_));
 sky130_fd_sc_hd__nand2_1 _12246_ (.A(_05377_),
    .B(_05362_),
    .Y(_05378_));
 sky130_fd_sc_hd__nand3_2 _12247_ (.A(_05354_),
    .B(_05376_),
    .C(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__inv_2 _12248_ (.A(_05354_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand2_1 _12249_ (.A(_05378_),
    .B(_05376_),
    .Y(_05381_));
 sky130_fd_sc_hd__nand2_1 _12250_ (.A(_05380_),
    .B(_05381_),
    .Y(_05383_));
 sky130_fd_sc_hd__nand2_1 _12251_ (.A(_05379_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__a31oi_1 _12252_ (.A1(_05257_),
    .A2(_06236_),
    .A3(_06179_),
    .B1(_05256_),
    .Y(_05385_));
 sky130_fd_sc_hd__nand2_1 _12253_ (.A(_06247_),
    .B(_06222_),
    .Y(_05386_));
 sky130_fd_sc_hd__and4_1 _12254_ (.A(_06239_),
    .B(net13),
    .C(_01280_),
    .D(_06173_),
    .X(_05387_));
 sky130_fd_sc_hd__a22o_1 _12255_ (.A1(_06239_),
    .A2(_01280_),
    .B1(net13),
    .B2(_06173_),
    .X(_05388_));
 sky130_fd_sc_hd__nand2b_1 _12256_ (.A_N(_05387_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__or2_1 _12257_ (.A(_05386_),
    .B(_05389_),
    .X(_05390_));
 sky130_fd_sc_hd__nand2_1 _12258_ (.A(_05389_),
    .B(_05386_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _12259_ (.A(_05390_),
    .B(_05391_),
    .Y(_05392_));
 sky130_fd_sc_hd__nor2_1 _12260_ (.A(_05385_),
    .B(_05392_),
    .Y(_05394_));
 sky130_fd_sc_hd__inv_2 _12261_ (.A(_05394_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand2_1 _12262_ (.A(_05392_),
    .B(_05385_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand2_1 _12263_ (.A(_05395_),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__and4_1 _12264_ (.A(_06240_),
    .B(_06243_),
    .C(_06172_),
    .D(_06174_),
    .X(_05398_));
 sky130_fd_sc_hd__inv_2 _12265_ (.A(_05277_),
    .Y(_05399_));
 sky130_fd_sc_hd__nor2_1 _12266_ (.A(_05398_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_1 _12267_ (.A(_05397_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__inv_2 _12268_ (.A(_05400_),
    .Y(_05402_));
 sky130_fd_sc_hd__nand3_1 _12269_ (.A(_05395_),
    .B(_05402_),
    .C(_05396_),
    .Y(_05403_));
 sky130_fd_sc_hd__nand2_1 _12270_ (.A(_05401_),
    .B(_05403_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_1 _12271_ (.A(_05384_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hd__inv_2 _12272_ (.A(_05405_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand3_1 _12273_ (.A(_05407_),
    .B(_05379_),
    .C(_05383_),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_1 _12274_ (.A(_05406_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand2_1 _12275_ (.A(_05291_),
    .B(_05267_),
    .Y(_05410_));
 sky130_fd_sc_hd__inv_2 _12276_ (.A(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_1 _12277_ (.A(_05409_),
    .B(_05411_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand3_1 _12278_ (.A(_05410_),
    .B(_05406_),
    .C(_05408_),
    .Y(_05413_));
 sky130_fd_sc_hd__nand2_1 _12279_ (.A(_05412_),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hd__or3b_2 _12280_ (.A(_06250_),
    .B(_04854_),
    .C_N(_06218_),
    .X(_05416_));
 sky130_fd_sc_hd__a21o_1 _12281_ (.A1(_03905_),
    .A2(_06223_),
    .B1(_06218_),
    .X(_05417_));
 sky130_fd_sc_hd__nand2_1 _12282_ (.A(_05416_),
    .B(_05417_),
    .Y(_05418_));
 sky130_fd_sc_hd__a21oi_1 _12283_ (.A1(_05301_),
    .A2(_06221_),
    .B1(_05300_),
    .Y(_05419_));
 sky130_fd_sc_hd__nor2_1 _12284_ (.A(_05418_),
    .B(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__inv_2 _12285_ (.A(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__nand2_1 _12286_ (.A(_05419_),
    .B(_05418_),
    .Y(_05422_));
 sky130_fd_sc_hd__nand2_1 _12287_ (.A(_05421_),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hd__a21o_1 _12288_ (.A1(_05287_),
    .A2(_05279_),
    .B1(_05423_),
    .X(_05424_));
 sky130_fd_sc_hd__nand3_1 _12289_ (.A(_05287_),
    .B(_05279_),
    .C(_05423_),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _12290_ (.A(_05424_),
    .B(_05425_),
    .Y(_05427_));
 sky130_fd_sc_hd__or2_1 _12291_ (.A(_05307_),
    .B(_05427_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_1 _12292_ (.A(_05427_),
    .B(_05307_),
    .Y(_05429_));
 sky130_fd_sc_hd__nand2_1 _12293_ (.A(_05428_),
    .B(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _12294_ (.A(_05414_),
    .B(_05430_),
    .Y(_05431_));
 sky130_fd_sc_hd__inv_2 _12295_ (.A(_05430_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand3_2 _12296_ (.A(_05412_),
    .B(_05413_),
    .C(_05432_),
    .Y(_05433_));
 sky130_fd_sc_hd__nand2_1 _12297_ (.A(_05431_),
    .B(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__nand2_1 _12298_ (.A(_05322_),
    .B(_05297_),
    .Y(_05435_));
 sky130_fd_sc_hd__inv_2 _12299_ (.A(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hd__nand2_1 _12300_ (.A(_05434_),
    .B(_05436_),
    .Y(_05438_));
 sky130_fd_sc_hd__nand3_2 _12301_ (.A(_05435_),
    .B(_05431_),
    .C(_05433_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_1 _12302_ (.A(_05438_),
    .B(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_1 _12303_ (.A(_05318_),
    .B(_05312_),
    .Y(_05441_));
 sky130_fd_sc_hd__inv_2 _12304_ (.A(_05441_),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_1 _12305_ (.A(_05440_),
    .B(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__nand3_1 _12306_ (.A(_05438_),
    .B(_05439_),
    .C(_05441_),
    .Y(_05444_));
 sky130_fd_sc_hd__nand2_1 _12307_ (.A(_05443_),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__nand2_1 _12308_ (.A(_05353_),
    .B(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__nor2_1 _12309_ (.A(_05445_),
    .B(_05353_),
    .Y(_05447_));
 sky130_fd_sc_hd__inv_2 _12310_ (.A(_05447_),
    .Y(_05449_));
 sky130_fd_sc_hd__nand3_1 _12311_ (.A(_05352_),
    .B(_05446_),
    .C(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__nand2_1 _12312_ (.A(_05449_),
    .B(_05446_),
    .Y(_05451_));
 sky130_fd_sc_hd__nor2_1 _12313_ (.A(_05335_),
    .B(_05334_),
    .Y(_05452_));
 sky130_fd_sc_hd__a21oi_1 _12314_ (.A1(_05336_),
    .A2(_05199_),
    .B1(_05452_),
    .Y(_05453_));
 sky130_fd_sc_hd__nand2_1 _12315_ (.A(_05451_),
    .B(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__nand2_1 _12316_ (.A(_05450_),
    .B(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand2_1 _12317_ (.A(_05455_),
    .B(_05341_),
    .Y(_05456_));
 sky130_fd_sc_hd__nor2_1 _12318_ (.A(_05343_),
    .B(_05342_),
    .Y(_05457_));
 sky130_fd_sc_hd__nand3_1 _12319_ (.A(_05457_),
    .B(_05450_),
    .C(_05454_),
    .Y(_05458_));
 sky130_fd_sc_hd__and2_1 _12320_ (.A(_05456_),
    .B(_05458_),
    .X(_05460_));
 sky130_fd_sc_hd__nor2_1 _12321_ (.A(_05225_),
    .B(_05349_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand2_1 _12322_ (.A(_05461_),
    .B(_05227_),
    .Y(_05462_));
 sky130_fd_sc_hd__inv_2 _12323_ (.A(_05462_),
    .Y(_05463_));
 sky130_fd_sc_hd__nand2_1 _12324_ (.A(_04950_),
    .B(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__nand2_1 _12325_ (.A(_05229_),
    .B(_05461_),
    .Y(_05465_));
 sky130_fd_sc_hd__inv_2 _12326_ (.A(_05224_),
    .Y(_05466_));
 sky130_fd_sc_hd__a21boi_1 _12327_ (.A1(_05466_),
    .A2(_05346_),
    .B1_N(_05348_),
    .Y(_05467_));
 sky130_fd_sc_hd__nand2_1 _12328_ (.A(_05465_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__inv_2 _12329_ (.A(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__nand2_1 _12330_ (.A(_05464_),
    .B(_05469_),
    .Y(_05471_));
 sky130_fd_sc_hd__or2_1 _12331_ (.A(_05460_),
    .B(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__nand2_1 _12332_ (.A(_05471_),
    .B(_05460_),
    .Y(_05473_));
 sky130_fd_sc_hd__and2_1 _12333_ (.A(_05472_),
    .B(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_1 _12334_ (.A(_05474_),
    .X(\m1.out[36] ));
 sky130_fd_sc_hd__nand2_1 _12335_ (.A(_05408_),
    .B(_05379_),
    .Y(_05475_));
 sky130_fd_sc_hd__or3_1 _12336_ (.A(_01422_),
    .B(_05363_),
    .C(_04801_),
    .X(_05476_));
 sky130_fd_sc_hd__a21o_1 _12337_ (.A1(_01831_),
    .A2(_06183_),
    .B1(_01158_),
    .X(_05477_));
 sky130_fd_sc_hd__nand2_1 _12338_ (.A(_05476_),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__nand2_1 _12339_ (.A(_01211_),
    .B(_02181_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_1 _12340_ (.A(_05478_),
    .B(_05479_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand3b_1 _12341_ (.A_N(_05479_),
    .B(_05476_),
    .C(_05477_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand2_1 _12342_ (.A(_05481_),
    .B(_05482_),
    .Y(_05483_));
 sky130_fd_sc_hd__and2_1 _12343_ (.A(_05370_),
    .B(_05364_),
    .X(_05484_));
 sky130_fd_sc_hd__or2_1 _12344_ (.A(_05483_),
    .B(_05484_),
    .X(_05485_));
 sky130_fd_sc_hd__nand2_1 _12345_ (.A(_05484_),
    .B(_05483_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand2_1 _12346_ (.A(_06240_),
    .B(_06179_),
    .Y(_05487_));
 sky130_fd_sc_hd__inv_2 _12347_ (.A(_06234_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand2_1 _12348_ (.A(_06242_),
    .B(_01692_),
    .Y(_05489_));
 sky130_fd_sc_hd__nor3_1 _12349_ (.A(_05488_),
    .B(_06188_),
    .C(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__o21ai_1 _12350_ (.A1(_05488_),
    .A2(_06188_),
    .B1(_05489_),
    .Y(_05492_));
 sky130_fd_sc_hd__and2b_1 _12351_ (.A_N(_05490_),
    .B(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__xor2_1 _12352_ (.A(_05487_),
    .B(_05493_),
    .X(_05494_));
 sky130_fd_sc_hd__inv_2 _12353_ (.A(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__a21o_1 _12354_ (.A1(_05485_),
    .A2(_05486_),
    .B1(_05495_),
    .X(_05496_));
 sky130_fd_sc_hd__nand3_1 _12355_ (.A(_05485_),
    .B(_05495_),
    .C(_05486_),
    .Y(_05497_));
 sky130_fd_sc_hd__nand2_1 _12356_ (.A(_05496_),
    .B(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__nand2_1 _12357_ (.A(_05376_),
    .B(_05374_),
    .Y(_05499_));
 sky130_fd_sc_hd__inv_2 _12358_ (.A(_05499_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_1 _12359_ (.A(_05498_),
    .B(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hd__nand3_1 _12360_ (.A(_05499_),
    .B(_05496_),
    .C(_05497_),
    .Y(_05503_));
 sky130_fd_sc_hd__nand2_1 _12361_ (.A(_05501_),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__nand2_1 _12362_ (.A(_03905_),
    .B(_06222_),
    .Y(_05505_));
 sky130_fd_sc_hd__and4_1 _12363_ (.A(_06245_),
    .B(net13),
    .C(net41),
    .D(net40),
    .X(_05506_));
 sky130_fd_sc_hd__a22o_1 _12364_ (.A1(net14),
    .A2(net40),
    .B1(net13),
    .B2(_01280_),
    .X(_05507_));
 sky130_fd_sc_hd__or2b_1 _12365_ (.A(_05506_),
    .B_N(_05507_),
    .X(_05508_));
 sky130_fd_sc_hd__or2_1 _12366_ (.A(_05505_),
    .B(_05508_),
    .X(_05509_));
 sky130_fd_sc_hd__nand2_1 _12367_ (.A(_05508_),
    .B(_05505_),
    .Y(_05510_));
 sky130_fd_sc_hd__nand2_1 _12368_ (.A(_05509_),
    .B(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__inv_2 _12369_ (.A(_05355_),
    .Y(_05512_));
 sky130_fd_sc_hd__a21oi_1 _12370_ (.A1(_05359_),
    .A2(_05512_),
    .B1(_05358_),
    .Y(_05514_));
 sky130_fd_sc_hd__inv_2 _12371_ (.A(_05514_),
    .Y(_05515_));
 sky130_fd_sc_hd__or2b_1 _12372_ (.A(_05511_),
    .B_N(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_1 _12373_ (.A(_05511_),
    .B(_05514_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_1 _12374_ (.A(_05516_),
    .B(_05517_),
    .Y(_05518_));
 sky130_fd_sc_hd__and2b_1 _12375_ (.A_N(_05387_),
    .B(_05390_),
    .X(_05519_));
 sky130_fd_sc_hd__nand2_1 _12376_ (.A(_05518_),
    .B(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__nand3b_1 _12377_ (.A_N(_05519_),
    .B(_05516_),
    .C(_05517_),
    .Y(_05521_));
 sky130_fd_sc_hd__nand2_1 _12378_ (.A(_05520_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nand2_1 _12379_ (.A(_05504_),
    .B(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__nand3b_1 _12380_ (.A_N(_05522_),
    .B(_05501_),
    .C(_05503_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand3_1 _12381_ (.A(_05475_),
    .B(_05523_),
    .C(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_1 _12382_ (.A(_05523_),
    .B(_05525_),
    .Y(_05527_));
 sky130_fd_sc_hd__a21boi_1 _12383_ (.A1(_05407_),
    .A2(_05383_),
    .B1_N(_05379_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _12384_ (.A(_05527_),
    .B(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__nand2_1 _12385_ (.A(_05526_),
    .B(_05529_),
    .Y(_05530_));
 sky130_fd_sc_hd__nand2_1 _12386_ (.A(_05416_),
    .B(_06223_),
    .Y(_05531_));
 sky130_fd_sc_hd__a21oi_1 _12387_ (.A1(_05396_),
    .A2(_05402_),
    .B1(_05394_),
    .Y(_05532_));
 sky130_fd_sc_hd__or2_1 _12388_ (.A(_05531_),
    .B(_05532_),
    .X(_05533_));
 sky130_fd_sc_hd__nand2_1 _12389_ (.A(_05532_),
    .B(_05531_),
    .Y(_05534_));
 sky130_fd_sc_hd__nand2_1 _12390_ (.A(_05533_),
    .B(_05534_),
    .Y(_05536_));
 sky130_fd_sc_hd__nand2_1 _12391_ (.A(_05536_),
    .B(_05421_),
    .Y(_05537_));
 sky130_fd_sc_hd__nand3_1 _12392_ (.A(_05533_),
    .B(_05420_),
    .C(_05534_),
    .Y(_05538_));
 sky130_fd_sc_hd__nand2_1 _12393_ (.A(_05537_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__nand2_1 _12394_ (.A(_05530_),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__nand3b_1 _12395_ (.A_N(_05539_),
    .B(_05526_),
    .C(_05529_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand2_1 _12396_ (.A(_05540_),
    .B(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand2_1 _12397_ (.A(_05433_),
    .B(_05413_),
    .Y(_05543_));
 sky130_fd_sc_hd__inv_2 _12398_ (.A(_05543_),
    .Y(_05544_));
 sky130_fd_sc_hd__nand2_1 _12399_ (.A(_05542_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__nand3_1 _12400_ (.A(_05543_),
    .B(_05540_),
    .C(_05541_),
    .Y(_05547_));
 sky130_fd_sc_hd__nand2_1 _12401_ (.A(_05545_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__nand2_1 _12402_ (.A(_05428_),
    .B(_05424_),
    .Y(_05549_));
 sky130_fd_sc_hd__inv_2 _12403_ (.A(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2_1 _12404_ (.A(_05548_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand3_2 _12405_ (.A(_05545_),
    .B(_05547_),
    .C(_05549_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand2_1 _12406_ (.A(_05551_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__nand3_1 _12407_ (.A(_05553_),
    .B(_05439_),
    .C(_05444_),
    .Y(_05554_));
 sky130_fd_sc_hd__nand2_1 _12408_ (.A(_05444_),
    .B(_05439_),
    .Y(_05555_));
 sky130_fd_sc_hd__nand3_2 _12409_ (.A(_05555_),
    .B(_05551_),
    .C(_05552_),
    .Y(_05556_));
 sky130_fd_sc_hd__nand2_1 _12410_ (.A(_05554_),
    .B(_05556_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_1 _12411_ (.A(_05558_),
    .B(_05449_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand3_2 _12412_ (.A(_05554_),
    .B(_05447_),
    .C(_05556_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_05559_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__nand2_1 _12414_ (.A(_05561_),
    .B(_05450_),
    .Y(_05562_));
 sky130_fd_sc_hd__nor2_1 _12415_ (.A(_05453_),
    .B(_05451_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand3_1 _12416_ (.A(_05563_),
    .B(_05559_),
    .C(_05560_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand2_1 _12417_ (.A(_05562_),
    .B(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__inv_2 _12418_ (.A(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand2_1 _12419_ (.A(_05473_),
    .B(_05458_),
    .Y(_05567_));
 sky130_fd_sc_hd__xor2_1 _12420_ (.A(_05566_),
    .B(_05567_),
    .X(\m1.out[37] ));
 sky130_fd_sc_hd__nand2_1 _12421_ (.A(_05541_),
    .B(_05526_),
    .Y(_05569_));
 sky130_fd_sc_hd__inv_2 _12422_ (.A(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__nand2_1 _12423_ (.A(_05482_),
    .B(_05476_),
    .Y(_05571_));
 sky130_fd_sc_hd__inv_2 _12424_ (.A(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2_1 _12425_ (.A(_06235_),
    .B(_02180_),
    .Y(_05573_));
 sky130_fd_sc_hd__or3_1 _12426_ (.A(_01422_),
    .B(_05356_),
    .C(_04801_),
    .X(_05574_));
 sky130_fd_sc_hd__a21o_1 _12427_ (.A1(_06237_),
    .A2(net47),
    .B1(_06281_),
    .X(_05575_));
 sky130_fd_sc_hd__nand2_1 _12428_ (.A(_05574_),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__or2_1 _12429_ (.A(_05573_),
    .B(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__nand2_1 _12430_ (.A(_05576_),
    .B(_05573_),
    .Y(_05579_));
 sky130_fd_sc_hd__nand2_1 _12431_ (.A(_05577_),
    .B(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__or2_1 _12432_ (.A(_05572_),
    .B(_05580_),
    .X(_05581_));
 sky130_fd_sc_hd__nand2_1 _12433_ (.A(_05580_),
    .B(_05572_),
    .Y(_05582_));
 sky130_fd_sc_hd__nand2_1 _12434_ (.A(_05581_),
    .B(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__nand2_1 _12435_ (.A(_06248_),
    .B(_06179_),
    .Y(_05584_));
 sky130_fd_sc_hd__and4_1 _12436_ (.A(_01858_),
    .B(_06241_),
    .C(_06175_),
    .D(_06187_),
    .X(_05585_));
 sky130_fd_sc_hd__inv_2 _12437_ (.A(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__a22o_1 _12438_ (.A1(_06240_),
    .A2(_06176_),
    .B1(_06243_),
    .B2(_01922_),
    .X(_05587_));
 sky130_fd_sc_hd__nand2_1 _12439_ (.A(_05586_),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__xnor2_1 _12440_ (.A(_05584_),
    .B(_05588_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand2_1 _12441_ (.A(_05583_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__nand3b_2 _12442_ (.A_N(_05590_),
    .B(_05581_),
    .C(_05582_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand2_1 _12443_ (.A(_05591_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__nand3_1 _12444_ (.A(_05593_),
    .B(_05485_),
    .C(_05497_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_1 _12445_ (.A(_05497_),
    .B(_05485_),
    .Y(_05595_));
 sky130_fd_sc_hd__nand3_2 _12446_ (.A(_05591_),
    .B(_05592_),
    .C(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__nand2_1 _12447_ (.A(_05594_),
    .B(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__a31oi_2 _12448_ (.A1(_05492_),
    .A2(_06240_),
    .A3(_06179_),
    .B1(_05490_),
    .Y(_05598_));
 sky130_fd_sc_hd__and4_1 _12449_ (.A(_06245_),
    .B(net15),
    .C(net41),
    .D(_06173_),
    .X(_05599_));
 sky130_fd_sc_hd__inv_2 _12450_ (.A(_05599_),
    .Y(_05601_));
 sky130_fd_sc_hd__a22o_1 _12451_ (.A1(_06245_),
    .A2(_06171_),
    .B1(_06298_),
    .B2(_01278_),
    .X(_05602_));
 sky130_fd_sc_hd__nand2_1 _12452_ (.A(_05601_),
    .B(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__inv_2 _12453_ (.A(_05603_),
    .Y(_05604_));
 sky130_fd_sc_hd__or2_1 _12454_ (.A(_06222_),
    .B(_05604_),
    .X(_05605_));
 sky130_fd_sc_hd__nand2_1 _12455_ (.A(_05604_),
    .B(_06222_),
    .Y(_05606_));
 sky130_fd_sc_hd__nand2_1 _12456_ (.A(_05605_),
    .B(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hd__or2_1 _12457_ (.A(_05598_),
    .B(_05607_),
    .X(_05608_));
 sky130_fd_sc_hd__nand2_1 _12458_ (.A(_05607_),
    .B(_05598_),
    .Y(_05609_));
 sky130_fd_sc_hd__nand2_1 _12459_ (.A(_05608_),
    .B(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__and2b_1 _12460_ (.A_N(_05506_),
    .B(_05509_),
    .X(_05612_));
 sky130_fd_sc_hd__nand2_1 _12461_ (.A(_05610_),
    .B(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand3b_1 _12462_ (.A_N(_05612_),
    .B(_05608_),
    .C(_05609_),
    .Y(_05614_));
 sky130_fd_sc_hd__nand2_1 _12463_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand2_1 _12464_ (.A(_05597_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__nand3b_2 _12465_ (.A_N(_05615_),
    .B(_05594_),
    .C(_05596_),
    .Y(_05617_));
 sky130_fd_sc_hd__nand2_1 _12466_ (.A(_05616_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__nand2_1 _12467_ (.A(_05525_),
    .B(_05503_),
    .Y(_05619_));
 sky130_fd_sc_hd__inv_2 _12468_ (.A(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__nand2_1 _12469_ (.A(_05618_),
    .B(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__nand3_1 _12470_ (.A(_05619_),
    .B(_05616_),
    .C(_05617_),
    .Y(_05623_));
 sky130_fd_sc_hd__nand2_1 _12471_ (.A(_05621_),
    .B(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__and2_1 _12472_ (.A(_05521_),
    .B(_05516_),
    .X(_05625_));
 sky130_fd_sc_hd__nor2_1 _12473_ (.A(_05416_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__inv_2 _12474_ (.A(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand2_1 _12475_ (.A(_05625_),
    .B(_05416_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_1 _12476_ (.A(_05627_),
    .B(_05628_),
    .Y(_05629_));
 sky130_fd_sc_hd__nand2_1 _12477_ (.A(_05624_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand3b_1 _12478_ (.A_N(_05629_),
    .B(_05621_),
    .C(_05623_),
    .Y(_05631_));
 sky130_fd_sc_hd__nand2_1 _12479_ (.A(_05630_),
    .B(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__nand2_1 _12480_ (.A(_05570_),
    .B(_05632_),
    .Y(_05634_));
 sky130_fd_sc_hd__nand3_1 _12481_ (.A(_05569_),
    .B(_05630_),
    .C(_05631_),
    .Y(_05635_));
 sky130_fd_sc_hd__nand2_1 _12482_ (.A(_05634_),
    .B(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__nand2_1 _12483_ (.A(_05538_),
    .B(_05533_),
    .Y(_05637_));
 sky130_fd_sc_hd__inv_2 _12484_ (.A(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__nand2_1 _12485_ (.A(_05636_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__nand3_1 _12486_ (.A(_05634_),
    .B(_05635_),
    .C(_05637_),
    .Y(_05640_));
 sky130_fd_sc_hd__nand2_1 _12487_ (.A(_05639_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(_05552_),
    .B(_05547_),
    .Y(_05642_));
 sky130_fd_sc_hd__inv_2 _12489_ (.A(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__nand2_1 _12490_ (.A(_05641_),
    .B(_05643_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand3_2 _12491_ (.A(_05642_),
    .B(_05639_),
    .C(_05640_),
    .Y(_05646_));
 sky130_fd_sc_hd__nand3b_2 _12492_ (.A_N(_05556_),
    .B(_05645_),
    .C(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_1 _12493_ (.A(_05645_),
    .B(_05646_),
    .Y(_05648_));
 sky130_fd_sc_hd__nand2_1 _12494_ (.A(_05648_),
    .B(_05556_),
    .Y(_05649_));
 sky130_fd_sc_hd__nand3b_1 _12495_ (.A_N(_05560_),
    .B(_05647_),
    .C(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__nand2_1 _12496_ (.A(_05649_),
    .B(_05647_),
    .Y(_05651_));
 sky130_fd_sc_hd__nand2_1 _12497_ (.A(_05651_),
    .B(_05560_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_1 _12498_ (.A(_05650_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__inv_2 _12499_ (.A(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_1 _12500_ (.A(_05460_),
    .B(_05566_),
    .Y(_05656_));
 sky130_fd_sc_hd__inv_2 _12501_ (.A(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand2_1 _12502_ (.A(_05471_),
    .B(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__o21ai_1 _12503_ (.A1(_05458_),
    .A2(_05565_),
    .B1(_05564_),
    .Y(_05659_));
 sky130_fd_sc_hd__inv_2 _12504_ (.A(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__nand2_1 _12505_ (.A(_05658_),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__or2_1 _12506_ (.A(_05654_),
    .B(_05661_),
    .X(_05662_));
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(_05661_),
    .B(_05654_),
    .Y(_05663_));
 sky130_fd_sc_hd__and2_1 _12508_ (.A(_05662_),
    .B(_05663_),
    .X(_05664_));
 sky130_fd_sc_hd__clkbuf_1 _12509_ (.A(_05664_),
    .X(\m1.out[38] ));
 sky130_fd_sc_hd__nand2_1 _12510_ (.A(_05663_),
    .B(_05650_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand2_1 _12511_ (.A(_06234_),
    .B(net47),
    .Y(_05667_));
 sky130_fd_sc_hd__xor2_1 _12512_ (.A(_06237_),
    .B(_05667_),
    .X(_05668_));
 sky130_fd_sc_hd__or3_1 _12513_ (.A(_04853_),
    .B(_06185_),
    .C(_05668_),
    .X(_05669_));
 sky130_fd_sc_hd__o21ai_1 _12514_ (.A1(_04853_),
    .A2(_06186_),
    .B1(_05668_),
    .Y(_05670_));
 sky130_fd_sc_hd__nand2_1 _12515_ (.A(_05669_),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__and2_1 _12516_ (.A(_05577_),
    .B(_05574_),
    .X(_05672_));
 sky130_fd_sc_hd__or2_1 _12517_ (.A(_05671_),
    .B(_05672_),
    .X(_05673_));
 sky130_fd_sc_hd__nand2_1 _12518_ (.A(_05672_),
    .B(_05671_),
    .Y(_05674_));
 sky130_fd_sc_hd__nand2_1 _12519_ (.A(_05673_),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__nand2_1 _12520_ (.A(_06246_),
    .B(_06178_),
    .Y(_05677_));
 sky130_fd_sc_hd__and4_1 _12521_ (.A(net11),
    .B(net13),
    .C(net43),
    .D(_06187_),
    .X(_05678_));
 sky130_fd_sc_hd__inv_2 _12522_ (.A(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__a22o_1 _12523_ (.A1(_01858_),
    .A2(_01921_),
    .B1(_02095_),
    .B2(_01692_),
    .X(_05680_));
 sky130_fd_sc_hd__nand2_1 _12524_ (.A(_05679_),
    .B(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__xnor2_1 _12525_ (.A(_05677_),
    .B(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__nand2_1 _12526_ (.A(_05675_),
    .B(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand3b_1 _12527_ (.A_N(_05682_),
    .B(_05673_),
    .C(_05674_),
    .Y(_05684_));
 sky130_fd_sc_hd__nand2_1 _12528_ (.A(_05683_),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand2_1 _12529_ (.A(_05592_),
    .B(_05581_),
    .Y(_05686_));
 sky130_fd_sc_hd__inv_2 _12530_ (.A(_05686_),
    .Y(_05688_));
 sky130_fd_sc_hd__nand2_1 _12531_ (.A(_05685_),
    .B(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__nand3_1 _12532_ (.A(_05686_),
    .B(_05683_),
    .C(_05684_),
    .Y(_05690_));
 sky130_fd_sc_hd__nand2_1 _12533_ (.A(_05689_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__and3_1 _12534_ (.A(_03905_),
    .B(_06172_),
    .C(_06174_),
    .X(_05692_));
 sky130_fd_sc_hd__inv_2 _12535_ (.A(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__a21o_1 _12536_ (.A1(_06299_),
    .A2(_06172_),
    .B1(_06174_),
    .X(_05694_));
 sky130_fd_sc_hd__nand2_1 _12537_ (.A(_05693_),
    .B(_05694_),
    .Y(_05695_));
 sky130_fd_sc_hd__o21a_1 _12538_ (.A1(_05584_),
    .A2(_05588_),
    .B1(_05586_),
    .X(_05696_));
 sky130_fd_sc_hd__nor2_1 _12539_ (.A(_05695_),
    .B(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hd__inv_2 _12540_ (.A(_05697_),
    .Y(_05699_));
 sky130_fd_sc_hd__nand2_1 _12541_ (.A(_05696_),
    .B(_05695_),
    .Y(_05700_));
 sky130_fd_sc_hd__nand2_1 _12542_ (.A(_05606_),
    .B(_05601_),
    .Y(_05701_));
 sky130_fd_sc_hd__a21o_1 _12543_ (.A1(_05699_),
    .A2(_05700_),
    .B1(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__nand3_1 _12544_ (.A(_05699_),
    .B(_05701_),
    .C(_05700_),
    .Y(_05703_));
 sky130_fd_sc_hd__nand2_1 _12545_ (.A(_05702_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__nand2_1 _12546_ (.A(_05691_),
    .B(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand3b_1 _12547_ (.A_N(_05704_),
    .B(_05689_),
    .C(_05690_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand2_1 _12548_ (.A(_05705_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__nand3_1 _12549_ (.A(_05707_),
    .B(_05596_),
    .C(_05617_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_1 _12550_ (.A(_05617_),
    .B(_05596_),
    .Y(_05710_));
 sky130_fd_sc_hd__nand3_1 _12551_ (.A(_05710_),
    .B(_05705_),
    .C(_05706_),
    .Y(_05711_));
 sky130_fd_sc_hd__nand2_1 _12552_ (.A(_05708_),
    .B(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__nand2_1 _12553_ (.A(_05614_),
    .B(_05608_),
    .Y(_05713_));
 sky130_fd_sc_hd__inv_2 _12554_ (.A(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__nand2_1 _12555_ (.A(_05712_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__nand3_1 _12556_ (.A(_05708_),
    .B(_05711_),
    .C(_05713_),
    .Y(_05716_));
 sky130_fd_sc_hd__nand2_1 _12557_ (.A(_05715_),
    .B(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__nand2_1 _12558_ (.A(_05631_),
    .B(_05623_),
    .Y(_05718_));
 sky130_fd_sc_hd__inv_2 _12559_ (.A(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__nand2_1 _12560_ (.A(_05717_),
    .B(_05719_),
    .Y(_05721_));
 sky130_fd_sc_hd__nand3_1 _12561_ (.A(_05718_),
    .B(_05715_),
    .C(_05716_),
    .Y(_05722_));
 sky130_fd_sc_hd__nand2_1 _12562_ (.A(_05721_),
    .B(_05722_),
    .Y(_05723_));
 sky130_fd_sc_hd__nand2_1 _12563_ (.A(_05723_),
    .B(_05627_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand3_1 _12564_ (.A(_05721_),
    .B(_05722_),
    .C(_05626_),
    .Y(_05725_));
 sky130_fd_sc_hd__nand2_1 _12565_ (.A(_05724_),
    .B(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_1 _12566_ (.A(_05640_),
    .B(_05635_),
    .Y(_05727_));
 sky130_fd_sc_hd__inv_2 _12567_ (.A(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__nand2_1 _12568_ (.A(_05726_),
    .B(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__nand3_2 _12569_ (.A(_05727_),
    .B(_05724_),
    .C(_05725_),
    .Y(_05730_));
 sky130_fd_sc_hd__nand3b_2 _12570_ (.A_N(_05646_),
    .B(_05729_),
    .C(_05730_),
    .Y(_05732_));
 sky130_fd_sc_hd__nand2_1 _12571_ (.A(_05729_),
    .B(_05730_),
    .Y(_05733_));
 sky130_fd_sc_hd__nand2_1 _12572_ (.A(_05733_),
    .B(_05646_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand3b_1 _12573_ (.A_N(_05647_),
    .B(_05732_),
    .C(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__nand2_1 _12574_ (.A(_05732_),
    .B(_05734_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand2_1 _12575_ (.A(_05736_),
    .B(_05647_),
    .Y(_05737_));
 sky130_fd_sc_hd__nand2_1 _12576_ (.A(_05735_),
    .B(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__nand2_1 _12577_ (.A(_05666_),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__inv_2 _12578_ (.A(_05738_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand3_1 _12579_ (.A(_05663_),
    .B(_05650_),
    .C(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _12580_ (.A(_05739_),
    .B(_05741_),
    .Y(\m1.out[39] ));
 sky130_fd_sc_hd__and2_1 _12581_ (.A(_05725_),
    .B(_05722_),
    .X(_05743_));
 sky130_fd_sc_hd__nand2_1 _12582_ (.A(_05706_),
    .B(_05690_),
    .Y(_05744_));
 sky130_fd_sc_hd__inv_2 _12583_ (.A(_05744_),
    .Y(_05745_));
 sky130_fd_sc_hd__and2_1 _12584_ (.A(_05684_),
    .B(_05673_),
    .X(_05746_));
 sky130_fd_sc_hd__nand2_1 _12585_ (.A(_03905_),
    .B(_06179_),
    .Y(_05747_));
 sky130_fd_sc_hd__inv_2 _12586_ (.A(net43),
    .Y(_05748_));
 sky130_fd_sc_hd__or4_1 _12587_ (.A(_02871_),
    .B(_03411_),
    .C(_05748_),
    .D(_06188_),
    .X(_05749_));
 sky130_fd_sc_hd__a22o_1 _12588_ (.A1(_06245_),
    .A2(_01692_),
    .B1(_06248_),
    .B2(_01921_),
    .X(_05750_));
 sky130_fd_sc_hd__nand2_1 _12589_ (.A(_05749_),
    .B(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__or2_1 _12590_ (.A(_05747_),
    .B(_05751_),
    .X(_05753_));
 sky130_fd_sc_hd__nand2_1 _12591_ (.A(_05751_),
    .B(_05747_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2_1 _12592_ (.A(_05753_),
    .B(_05754_),
    .Y(_05755_));
 sky130_fd_sc_hd__nand2_1 _12593_ (.A(_06241_),
    .B(net47),
    .Y(_05756_));
 sky130_fd_sc_hd__xor2_1 _12594_ (.A(_06234_),
    .B(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__or3_1 _12595_ (.A(_04495_),
    .B(_06185_),
    .C(_05757_),
    .X(_05758_));
 sky130_fd_sc_hd__o21ai_1 _12596_ (.A1(_04495_),
    .A2(_06186_),
    .B1(_05757_),
    .Y(_05759_));
 sky130_fd_sc_hd__nand2_1 _12597_ (.A(_05758_),
    .B(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__o21a_1 _12598_ (.A1(_05356_),
    .A2(_05667_),
    .B1(_05669_),
    .X(_05761_));
 sky130_fd_sc_hd__nor2_1 _12599_ (.A(_05760_),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand2_1 _12600_ (.A(_05761_),
    .B(_05760_),
    .Y(_05764_));
 sky130_fd_sc_hd__nand2b_1 _12601_ (.A_N(_05762_),
    .B(_05764_),
    .Y(_05765_));
 sky130_fd_sc_hd__nor2_1 _12602_ (.A(_05755_),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__inv_2 _12603_ (.A(_05766_),
    .Y(_05767_));
 sky130_fd_sc_hd__nand2_1 _12604_ (.A(_05765_),
    .B(_05755_),
    .Y(_05768_));
 sky130_fd_sc_hd__nand2_1 _12605_ (.A(_05767_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__nor2_1 _12606_ (.A(_05746_),
    .B(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__inv_2 _12607_ (.A(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _12608_ (.A(_05769_),
    .B(_05746_),
    .Y(_05772_));
 sky130_fd_sc_hd__inv_2 _12609_ (.A(_06172_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21a_1 _12610_ (.A1(_05677_),
    .A2(_05681_),
    .B1(_05679_),
    .X(_05775_));
 sky130_fd_sc_hd__nor2_1 _12611_ (.A(_05773_),
    .B(_05775_),
    .Y(_05776_));
 sky130_fd_sc_hd__inv_2 _12612_ (.A(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_1 _12613_ (.A(_05775_),
    .B(_05773_),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_1 _12614_ (.A(_05777_),
    .B(_05778_),
    .Y(_05779_));
 sky130_fd_sc_hd__or2_1 _12615_ (.A(_05693_),
    .B(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__nand2_1 _12616_ (.A(_05779_),
    .B(_05693_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_1 _12617_ (.A(_05780_),
    .B(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__inv_2 _12618_ (.A(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__a21o_1 _12619_ (.A1(_05771_),
    .A2(_05772_),
    .B1(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__nand3_1 _12620_ (.A(_05771_),
    .B(_05783_),
    .C(_05772_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand2_1 _12621_ (.A(_05784_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__or2_1 _12622_ (.A(_05745_),
    .B(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__nand2_1 _12623_ (.A(_05787_),
    .B(_05745_),
    .Y(_05789_));
 sky130_fd_sc_hd__nand2_1 _12624_ (.A(_05703_),
    .B(_05699_),
    .Y(_05790_));
 sky130_fd_sc_hd__a21o_1 _12625_ (.A1(_05788_),
    .A2(_05789_),
    .B1(_05790_),
    .X(_05791_));
 sky130_fd_sc_hd__nand3_1 _12626_ (.A(_05788_),
    .B(_05790_),
    .C(_05789_),
    .Y(_05792_));
 sky130_fd_sc_hd__nand2_1 _12627_ (.A(_05791_),
    .B(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__nand2_1 _12628_ (.A(_05716_),
    .B(_05711_),
    .Y(_05794_));
 sky130_fd_sc_hd__inv_2 _12629_ (.A(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand2_1 _12630_ (.A(_05793_),
    .B(_05795_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand3_1 _12631_ (.A(_05791_),
    .B(_05794_),
    .C(_05792_),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_1 _12632_ (.A(_05797_),
    .B(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__nor2_1 _12633_ (.A(_05743_),
    .B(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__inv_2 _12634_ (.A(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__nand2_1 _12635_ (.A(_05799_),
    .B(_05743_),
    .Y(_05802_));
 sky130_fd_sc_hd__nand2_1 _12636_ (.A(_05801_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand2_1 _12637_ (.A(_05803_),
    .B(_05730_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand3b_2 _12638_ (.A_N(_05730_),
    .B(_05801_),
    .C(_05802_),
    .Y(_05805_));
 sky130_fd_sc_hd__nand2_1 _12639_ (.A(_05804_),
    .B(_05805_),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_1 _12640_ (.A(_05806_),
    .B(_05732_),
    .Y(_05808_));
 sky130_fd_sc_hd__inv_2 _12641_ (.A(_05732_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand3_1 _12642_ (.A(_05804_),
    .B(_05805_),
    .C(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__nand2_1 _12643_ (.A(_05808_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__inv_2 _12644_ (.A(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__nand2_1 _12645_ (.A(_05740_),
    .B(_05654_),
    .Y(_05813_));
 sky130_fd_sc_hd__nor3_1 _12646_ (.A(_05813_),
    .B(_05656_),
    .C(_05462_),
    .Y(_05814_));
 sky130_fd_sc_hd__nand2_1 _12647_ (.A(_04950_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__nor2_1 _12648_ (.A(_05813_),
    .B(_05656_),
    .Y(_05816_));
 sky130_fd_sc_hd__nor2_1 _12649_ (.A(_05653_),
    .B(_05738_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_1 _12650_ (.A(_05659_),
    .B(_05817_),
    .Y(_05819_));
 sky130_fd_sc_hd__nor2_1 _12651_ (.A(_05560_),
    .B(_05651_),
    .Y(_05820_));
 sky130_fd_sc_hd__a21boi_1 _12652_ (.A1(_05820_),
    .A2(_05737_),
    .B1_N(_05735_),
    .Y(_05821_));
 sky130_fd_sc_hd__nand2_1 _12653_ (.A(_05819_),
    .B(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__a21oi_1 _12654_ (.A1(_05468_),
    .A2(_05816_),
    .B1(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__nand2_1 _12655_ (.A(_05815_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__or2_1 _12656_ (.A(_05812_),
    .B(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__nand2_1 _12657_ (.A(_05824_),
    .B(_05812_),
    .Y(_05826_));
 sky130_fd_sc_hd__and2_1 _12658_ (.A(_05825_),
    .B(_05826_),
    .X(_05827_));
 sky130_fd_sc_hd__clkbuf_1 _12659_ (.A(_05827_),
    .X(\m1.out[40] ));
 sky130_fd_sc_hd__nand2_1 _12660_ (.A(_05786_),
    .B(_05771_),
    .Y(_05829_));
 sky130_fd_sc_hd__inv_2 _12661_ (.A(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__nor2_1 _12662_ (.A(_05762_),
    .B(_05766_),
    .Y(_05831_));
 sky130_fd_sc_hd__inv_2 _12663_ (.A(_06179_),
    .Y(_05832_));
 sky130_fd_sc_hd__or4_1 _12664_ (.A(_02871_),
    .B(_06250_),
    .C(_05748_),
    .D(_06188_),
    .X(_05833_));
 sky130_fd_sc_hd__a22o_1 _12665_ (.A1(_06246_),
    .A2(_01922_),
    .B1(_03905_),
    .B2(_06176_),
    .X(_05834_));
 sky130_fd_sc_hd__nand2_1 _12666_ (.A(_05833_),
    .B(_05834_),
    .Y(_05835_));
 sky130_fd_sc_hd__or2_1 _12667_ (.A(_05832_),
    .B(_05835_),
    .X(_05836_));
 sky130_fd_sc_hd__nand2_1 _12668_ (.A(_05835_),
    .B(_05832_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_1 _12669_ (.A(_05836_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_1 _12670_ (.A(_06239_),
    .B(net47),
    .Y(_05840_));
 sky130_fd_sc_hd__xor2_1 _12671_ (.A(_06241_),
    .B(_05840_),
    .X(_05841_));
 sky130_fd_sc_hd__or3_1 _12672_ (.A(_03411_),
    .B(_06185_),
    .C(_05841_),
    .X(_05842_));
 sky130_fd_sc_hd__o21ai_1 _12673_ (.A1(_03411_),
    .A2(_06186_),
    .B1(_05841_),
    .Y(_05843_));
 sky130_fd_sc_hd__nand2_1 _12674_ (.A(_05842_),
    .B(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__o21a_1 _12675_ (.A1(_05488_),
    .A2(_05756_),
    .B1(_05758_),
    .X(_05845_));
 sky130_fd_sc_hd__nor2_1 _12676_ (.A(_05844_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _12677_ (.A(_05845_),
    .B(_05844_),
    .Y(_05847_));
 sky130_fd_sc_hd__nand2b_1 _12678_ (.A_N(_05846_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__nor2_1 _12679_ (.A(_05838_),
    .B(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__inv_2 _12680_ (.A(_05849_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand2_1 _12681_ (.A(_05848_),
    .B(_05838_),
    .Y(_05852_));
 sky130_fd_sc_hd__nand2_1 _12682_ (.A(_05851_),
    .B(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__nor2_1 _12683_ (.A(_05831_),
    .B(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__inv_2 _12684_ (.A(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__nand2_1 _12685_ (.A(_05853_),
    .B(_05831_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(_05753_),
    .B(_05749_),
    .Y(_05857_));
 sky130_fd_sc_hd__a21o_1 _12687_ (.A1(_05855_),
    .A2(_05856_),
    .B1(_05857_),
    .X(_05858_));
 sky130_fd_sc_hd__nand3_1 _12688_ (.A(_05855_),
    .B(_05857_),
    .C(_05856_),
    .Y(_05859_));
 sky130_fd_sc_hd__nand2_1 _12689_ (.A(_05858_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__or2_1 _12690_ (.A(_05830_),
    .B(_05860_),
    .X(_05862_));
 sky130_fd_sc_hd__nand2_1 _12691_ (.A(_05860_),
    .B(_05830_),
    .Y(_05863_));
 sky130_fd_sc_hd__nand2_1 _12692_ (.A(_05780_),
    .B(_05777_),
    .Y(_05864_));
 sky130_fd_sc_hd__a21o_1 _12693_ (.A1(_05862_),
    .A2(_05863_),
    .B1(_05864_),
    .X(_05865_));
 sky130_fd_sc_hd__nand3_1 _12694_ (.A(_05862_),
    .B(_05864_),
    .C(_05863_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand2_1 _12695_ (.A(_05865_),
    .B(_05866_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand2_1 _12696_ (.A(_05792_),
    .B(_05788_),
    .Y(_05868_));
 sky130_fd_sc_hd__inv_2 _12697_ (.A(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__nand2_1 _12698_ (.A(_05867_),
    .B(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__nand3_2 _12699_ (.A(_05865_),
    .B(_05868_),
    .C(_05866_),
    .Y(_05871_));
 sky130_fd_sc_hd__nand3b_1 _12700_ (.A_N(_05798_),
    .B(_05870_),
    .C(_05871_),
    .Y(_05873_));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(_05870_),
    .B(_05871_),
    .Y(_05874_));
 sky130_fd_sc_hd__nand2_1 _12702_ (.A(_05874_),
    .B(_05798_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand2_1 _12703_ (.A(_05873_),
    .B(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__nand2_1 _12704_ (.A(_05876_),
    .B(_05801_),
    .Y(_05877_));
 sky130_fd_sc_hd__nand3_1 _12705_ (.A(_05873_),
    .B(_05800_),
    .C(_05875_),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_1 _12706_ (.A(_05877_),
    .B(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__xor2_1 _12707_ (.A(_05805_),
    .B(_05879_),
    .X(_05880_));
 sky130_fd_sc_hd__nand2_1 _12708_ (.A(_05826_),
    .B(_05810_),
    .Y(_05881_));
 sky130_fd_sc_hd__xor2_1 _12709_ (.A(_05880_),
    .B(_05881_),
    .X(\m1.out[41] ));
 sky130_fd_sc_hd__and2_1 _12710_ (.A(_05859_),
    .B(_05855_),
    .X(_05883_));
 sky130_fd_sc_hd__nand2_1 _12711_ (.A(_05836_),
    .B(_05833_),
    .Y(_05884_));
 sky130_fd_sc_hd__nor2_1 _12712_ (.A(_05846_),
    .B(_05849_),
    .Y(_05885_));
 sky130_fd_sc_hd__and3_1 _12713_ (.A(_06299_),
    .B(_06176_),
    .C(_01922_),
    .X(_05886_));
 sky130_fd_sc_hd__inv_2 _12714_ (.A(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__a21o_1 _12715_ (.A1(_06299_),
    .A2(_01922_),
    .B1(_06176_),
    .X(_05888_));
 sky130_fd_sc_hd__nand2_1 _12716_ (.A(_05887_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__nand2_1 _12717_ (.A(_02095_),
    .B(_06183_),
    .Y(_05890_));
 sky130_fd_sc_hd__xor2_1 _12718_ (.A(_01858_),
    .B(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__or3_1 _12719_ (.A(_02871_),
    .B(_06186_),
    .C(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__o21ai_1 _12720_ (.A1(_02871_),
    .A2(_06186_),
    .B1(_05891_),
    .Y(_05894_));
 sky130_fd_sc_hd__nand2_1 _12721_ (.A(_05892_),
    .B(_05894_),
    .Y(_05895_));
 sky130_fd_sc_hd__o21a_1 _12722_ (.A1(_04853_),
    .A2(_05840_),
    .B1(_05842_),
    .X(_05896_));
 sky130_fd_sc_hd__nor2_1 _12723_ (.A(_05895_),
    .B(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_1 _12724_ (.A(_05896_),
    .B(_05895_),
    .Y(_05898_));
 sky130_fd_sc_hd__nand2b_1 _12725_ (.A_N(_05897_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__or2_1 _12726_ (.A(_05889_),
    .B(_05899_),
    .X(_05900_));
 sky130_fd_sc_hd__nand2_1 _12727_ (.A(_05899_),
    .B(_05889_),
    .Y(_05901_));
 sky130_fd_sc_hd__nand2_1 _12728_ (.A(_05900_),
    .B(_05901_),
    .Y(_05902_));
 sky130_fd_sc_hd__nor2_1 _12729_ (.A(_05885_),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__nand2_1 _12730_ (.A(_05902_),
    .B(_05885_),
    .Y(_05905_));
 sky130_fd_sc_hd__nand2b_1 _12731_ (.A_N(_05903_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__xor2_1 _12732_ (.A(_05884_),
    .B(_05906_),
    .X(_05907_));
 sky130_fd_sc_hd__nor2_1 _12733_ (.A(_05883_),
    .B(_05907_),
    .Y(_05908_));
 sky130_fd_sc_hd__nand2_1 _12734_ (.A(_05907_),
    .B(_05883_),
    .Y(_05909_));
 sky130_fd_sc_hd__or2b_1 _12735_ (.A(_05908_),
    .B_N(_05909_),
    .X(_05910_));
 sky130_fd_sc_hd__a21boi_1 _12736_ (.A1(_05864_),
    .A2(_05863_),
    .B1_N(_05862_),
    .Y(_05911_));
 sky130_fd_sc_hd__or2_1 _12737_ (.A(_05910_),
    .B(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__nand2_1 _12738_ (.A(_05911_),
    .B(_05910_),
    .Y(_05913_));
 sky130_fd_sc_hd__nand2_1 _12739_ (.A(_05912_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__nand2_1 _12740_ (.A(_05914_),
    .B(_05871_),
    .Y(_05916_));
 sky130_fd_sc_hd__inv_2 _12741_ (.A(_05871_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand3_2 _12742_ (.A(_05917_),
    .B(_05912_),
    .C(_05913_),
    .Y(_05918_));
 sky130_fd_sc_hd__nand2_1 _12743_ (.A(_05916_),
    .B(_05918_),
    .Y(_05919_));
 sky130_fd_sc_hd__nand2_1 _12744_ (.A(_05919_),
    .B(_05873_),
    .Y(_05920_));
 sky130_fd_sc_hd__nor2_1 _12745_ (.A(_05798_),
    .B(_05874_),
    .Y(_05921_));
 sky130_fd_sc_hd__nand3_1 _12746_ (.A(_05921_),
    .B(_05916_),
    .C(_05918_),
    .Y(_05922_));
 sky130_fd_sc_hd__nand2_1 _12747_ (.A(_05920_),
    .B(_05922_),
    .Y(_05923_));
 sky130_fd_sc_hd__or2_1 _12748_ (.A(_05878_),
    .B(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__nand2_1 _12749_ (.A(_05923_),
    .B(_05878_),
    .Y(_05925_));
 sky130_fd_sc_hd__nand2_1 _12750_ (.A(_05924_),
    .B(_05925_),
    .Y(_05927_));
 sky130_fd_sc_hd__inv_2 _12751_ (.A(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _12752_ (.A(_05812_),
    .B(_05880_),
    .Y(_05929_));
 sky130_fd_sc_hd__inv_2 _12753_ (.A(_05929_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand2_1 _12754_ (.A(_05824_),
    .B(_05930_),
    .Y(_05931_));
 sky130_fd_sc_hd__inv_2 _12755_ (.A(_05810_),
    .Y(_05932_));
 sky130_fd_sc_hd__nand2_1 _12756_ (.A(_05879_),
    .B(_05805_),
    .Y(_05933_));
 sky130_fd_sc_hd__nor2_1 _12757_ (.A(_05805_),
    .B(_05879_),
    .Y(_05934_));
 sky130_fd_sc_hd__a21o_1 _12758_ (.A1(_05932_),
    .A2(_05933_),
    .B1(_05934_),
    .X(_05935_));
 sky130_fd_sc_hd__inv_2 _12759_ (.A(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__nand2_1 _12760_ (.A(_05931_),
    .B(_05936_),
    .Y(_05938_));
 sky130_fd_sc_hd__or2_1 _12761_ (.A(_05928_),
    .B(_05938_),
    .X(_05939_));
 sky130_fd_sc_hd__nand2_1 _12762_ (.A(_05938_),
    .B(_05928_),
    .Y(_05940_));
 sky130_fd_sc_hd__and2_1 _12763_ (.A(_05939_),
    .B(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__clkbuf_1 _12764_ (.A(_05941_),
    .X(\m1.out[42] ));
 sky130_fd_sc_hd__nand2_1 _12765_ (.A(_05940_),
    .B(_05924_),
    .Y(_05942_));
 sky130_fd_sc_hd__inv_2 _12766_ (.A(_05918_),
    .Y(_05943_));
 sky130_fd_sc_hd__nand2_1 _12767_ (.A(_06246_),
    .B(_02423_),
    .Y(_05944_));
 sky130_fd_sc_hd__xor2_1 _12768_ (.A(_06248_),
    .B(_05944_),
    .X(_05945_));
 sky130_fd_sc_hd__or3_1 _12769_ (.A(_06250_),
    .B(_06186_),
    .C(_05945_),
    .X(_05946_));
 sky130_fd_sc_hd__o21ai_1 _12770_ (.A1(_06250_),
    .A2(_06186_),
    .B1(_05945_),
    .Y(_05948_));
 sky130_fd_sc_hd__nand2_1 _12771_ (.A(_05946_),
    .B(_05948_),
    .Y(_05949_));
 sky130_fd_sc_hd__o21a_1 _12772_ (.A1(_04495_),
    .A2(_05890_),
    .B1(_05892_),
    .X(_05950_));
 sky130_fd_sc_hd__nor2_1 _12773_ (.A(_05949_),
    .B(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand2_1 _12774_ (.A(_05950_),
    .B(_05949_),
    .Y(_05952_));
 sky130_fd_sc_hd__or2b_1 _12775_ (.A(_05951_),
    .B_N(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__xor2_1 _12776_ (.A(_01922_),
    .B(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__and2b_1 _12777_ (.A_N(_05897_),
    .B(_05900_),
    .X(_05955_));
 sky130_fd_sc_hd__nor2_1 _12778_ (.A(_05954_),
    .B(_05955_),
    .Y(_05956_));
 sky130_fd_sc_hd__inv_2 _12779_ (.A(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__nand2_1 _12780_ (.A(_05955_),
    .B(_05954_),
    .Y(_05959_));
 sky130_fd_sc_hd__nand2_1 _12781_ (.A(_05957_),
    .B(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__or2_1 _12782_ (.A(_05887_),
    .B(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__nand2_1 _12783_ (.A(_05960_),
    .B(_05887_),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_1 _12784_ (.A(_05961_),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__a21oi_1 _12785_ (.A1(_05905_),
    .A2(_05884_),
    .B1(_05903_),
    .Y(_05964_));
 sky130_fd_sc_hd__nand2_1 _12786_ (.A(_05963_),
    .B(_05964_),
    .Y(_05965_));
 sky130_fd_sc_hd__nand3b_2 _12787_ (.A_N(_05964_),
    .B(_05961_),
    .C(_05962_),
    .Y(_05966_));
 sky130_fd_sc_hd__a21o_1 _12788_ (.A1(_05965_),
    .A2(_05966_),
    .B1(_05908_),
    .X(_05967_));
 sky130_fd_sc_hd__nand3_1 _12789_ (.A(_05965_),
    .B(_05966_),
    .C(_05908_),
    .Y(_05968_));
 sky130_fd_sc_hd__nand2_1 _12790_ (.A(_05967_),
    .B(_05968_),
    .Y(_05970_));
 sky130_fd_sc_hd__nor2_1 _12791_ (.A(_05910_),
    .B(_05911_),
    .Y(_05971_));
 sky130_fd_sc_hd__nand2b_1 _12792_ (.A_N(_05970_),
    .B(_05971_),
    .Y(_05972_));
 sky130_fd_sc_hd__nand2_1 _12793_ (.A(_05912_),
    .B(_05970_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand3_1 _12794_ (.A(_05943_),
    .B(_05972_),
    .C(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__nand2_1 _12795_ (.A(_05972_),
    .B(_05973_),
    .Y(_05975_));
 sky130_fd_sc_hd__nand2_1 _12796_ (.A(_05975_),
    .B(_05918_),
    .Y(_05976_));
 sky130_fd_sc_hd__nand2_1 _12797_ (.A(_05974_),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__nor2_1 _12798_ (.A(_05922_),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__inv_2 _12799_ (.A(_05978_),
    .Y(_05979_));
 sky130_fd_sc_hd__nand2_1 _12800_ (.A(_05977_),
    .B(_05922_),
    .Y(_05981_));
 sky130_fd_sc_hd__nand2_1 _12801_ (.A(_05979_),
    .B(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__nand2_1 _12802_ (.A(_05942_),
    .B(_05982_),
    .Y(_05983_));
 sky130_fd_sc_hd__nand3b_1 _12803_ (.A_N(_05982_),
    .B(_05940_),
    .C(_05924_),
    .Y(_05984_));
 sky130_fd_sc_hd__nand2_1 _12804_ (.A(_05983_),
    .B(_05984_),
    .Y(\m1.out[43] ));
 sky130_fd_sc_hd__nand2_2 _12805_ (.A(_06299_),
    .B(_06184_),
    .Y(_05985_));
 sky130_fd_sc_hd__inv_2 _12806_ (.A(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__nand2_1 _12807_ (.A(_05986_),
    .B(_06247_),
    .Y(_05987_));
 sky130_fd_sc_hd__nand2_1 _12808_ (.A(_05985_),
    .B(_02871_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand2_1 _12809_ (.A(_05987_),
    .B(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__or2_1 _12810_ (.A(_06186_),
    .B(_05989_),
    .X(_05991_));
 sky130_fd_sc_hd__nand2_1 _12811_ (.A(_05989_),
    .B(_06186_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand2_1 _12812_ (.A(_05991_),
    .B(_05992_),
    .Y(_05993_));
 sky130_fd_sc_hd__o21a_1 _12813_ (.A1(_03411_),
    .A2(_05944_),
    .B1(_05946_),
    .X(_05994_));
 sky130_fd_sc_hd__nor2_1 _12814_ (.A(_05993_),
    .B(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand2_1 _12815_ (.A(_05994_),
    .B(_05993_),
    .Y(_05996_));
 sky130_fd_sc_hd__or2b_1 _12816_ (.A(_05995_),
    .B_N(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__a21oi_1 _12817_ (.A1(_05952_),
    .A2(_01922_),
    .B1(_05951_),
    .Y(_05998_));
 sky130_fd_sc_hd__nor2_1 _12818_ (.A(_05997_),
    .B(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__nand2_1 _12819_ (.A(_05998_),
    .B(_05997_),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2b_1 _12820_ (.A_N(_05999_),
    .B(_06000_),
    .Y(_06002_));
 sky130_fd_sc_hd__and2_1 _12821_ (.A(_05961_),
    .B(_05957_),
    .X(_06003_));
 sky130_fd_sc_hd__xnor2_1 _12822_ (.A(_06002_),
    .B(_06003_),
    .Y(_06004_));
 sky130_fd_sc_hd__or2_1 _12823_ (.A(_05966_),
    .B(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__nand2_1 _12824_ (.A(_06004_),
    .B(_05966_),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2_1 _12825_ (.A(_06005_),
    .B(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__or2_1 _12826_ (.A(_05968_),
    .B(_06007_),
    .X(_06008_));
 sky130_fd_sc_hd__nand2_1 _12827_ (.A(_06007_),
    .B(_05968_),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2_1 _12828_ (.A(_06008_),
    .B(_06009_),
    .Y(_06010_));
 sky130_fd_sc_hd__nor2_1 _12829_ (.A(_05972_),
    .B(_06010_),
    .Y(_06011_));
 sky130_fd_sc_hd__inv_2 _12830_ (.A(_06011_),
    .Y(_06013_));
 sky130_fd_sc_hd__nand2_1 _12831_ (.A(_06010_),
    .B(_05972_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_1 _12832_ (.A(_06013_),
    .B(_06014_),
    .Y(_06015_));
 sky130_fd_sc_hd__or2_1 _12833_ (.A(_05974_),
    .B(_06015_),
    .X(_06016_));
 sky130_fd_sc_hd__nand2_1 _12834_ (.A(_06015_),
    .B(_05974_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand2_1 _12835_ (.A(_06016_),
    .B(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__inv_2 _12836_ (.A(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__nor2_1 _12837_ (.A(_05982_),
    .B(_05927_),
    .Y(_06020_));
 sky130_fd_sc_hd__nor2b_1 _12838_ (.A(_05929_),
    .B_N(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__nand2_1 _12839_ (.A(_05824_),
    .B(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__o21ai_1 _12840_ (.A1(_05924_),
    .A2(_05982_),
    .B1(_05979_),
    .Y(_06024_));
 sky130_fd_sc_hd__a21oi_1 _12841_ (.A1(_05935_),
    .A2(_06020_),
    .B1(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2_1 _12842_ (.A(_06022_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__or2_1 _12843_ (.A(_06019_),
    .B(_06026_),
    .X(_06027_));
 sky130_fd_sc_hd__nand2_1 _12844_ (.A(_06026_),
    .B(_06019_),
    .Y(_06028_));
 sky130_fd_sc_hd__and2_1 _12845_ (.A(_06027_),
    .B(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__clkbuf_1 _12846_ (.A(_06029_),
    .X(\m1.out[44] ));
 sky130_fd_sc_hd__nand2_1 _12847_ (.A(_06028_),
    .B(_06016_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand2_1 _12848_ (.A(_06250_),
    .B(_04801_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand2_1 _12849_ (.A(_06031_),
    .B(_05985_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand2_1 _12850_ (.A(_05991_),
    .B(_05987_),
    .Y(_06034_));
 sky130_fd_sc_hd__xor2_1 _12851_ (.A(_06032_),
    .B(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__nor2_1 _12852_ (.A(_06035_),
    .B(_05995_),
    .Y(_06036_));
 sky130_fd_sc_hd__or2_1 _12853_ (.A(_06036_),
    .B(_05999_),
    .X(_06037_));
 sky130_fd_sc_hd__nand2_1 _12854_ (.A(_05999_),
    .B(_06036_),
    .Y(_06038_));
 sky130_fd_sc_hd__nand2_1 _12855_ (.A(_06037_),
    .B(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__or3_1 _12856_ (.A(_06002_),
    .B(_06039_),
    .C(_06003_),
    .X(_06040_));
 sky130_fd_sc_hd__o21ai_1 _12857_ (.A1(_06002_),
    .A2(_06003_),
    .B1(_06039_),
    .Y(_06041_));
 sky130_fd_sc_hd__and2_1 _12858_ (.A(_06040_),
    .B(_06041_),
    .X(_06042_));
 sky130_fd_sc_hd__xor2_1 _12859_ (.A(_06005_),
    .B(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__or2_1 _12860_ (.A(_06008_),
    .B(_06043_),
    .X(_06045_));
 sky130_fd_sc_hd__nand2_1 _12861_ (.A(_06043_),
    .B(_06008_),
    .Y(_06046_));
 sky130_fd_sc_hd__nand2_1 _12862_ (.A(_06045_),
    .B(_06046_),
    .Y(_06047_));
 sky130_fd_sc_hd__nor2_1 _12863_ (.A(_06013_),
    .B(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__nand2_1 _12864_ (.A(_06047_),
    .B(_06013_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand2b_1 _12865_ (.A_N(_06048_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_1 _12866_ (.A(_06030_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand3b_1 _12867_ (.A_N(_06050_),
    .B(_06028_),
    .C(_06016_),
    .Y(_06052_));
 sky130_fd_sc_hd__nand2_1 _12868_ (.A(_06051_),
    .B(_06052_),
    .Y(\m1.out[45] ));
 sky130_fd_sc_hd__nor2_1 _12869_ (.A(_06018_),
    .B(_06050_),
    .Y(_06053_));
 sky130_fd_sc_hd__nand2_1 _12870_ (.A(_06026_),
    .B(_06053_),
    .Y(_06055_));
 sky130_fd_sc_hd__o21ba_1 _12871_ (.A1(_06016_),
    .A2(_06050_),
    .B1_N(_06048_),
    .X(_06056_));
 sky130_fd_sc_hd__nand2_1 _12872_ (.A(_06055_),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__and2b_1 _12873_ (.A_N(_06005_),
    .B(_06042_),
    .X(_06058_));
 sky130_fd_sc_hd__a31o_1 _12874_ (.A1(_06031_),
    .A2(_06247_),
    .A3(_02181_),
    .B1(_05986_),
    .X(_06059_));
 sky130_fd_sc_hd__xor2_1 _12875_ (.A(_06059_),
    .B(_05995_),
    .X(_06060_));
 sky130_fd_sc_hd__xnor2_1 _12876_ (.A(_06060_),
    .B(_06038_),
    .Y(_06061_));
 sky130_fd_sc_hd__or2_1 _12877_ (.A(_06061_),
    .B(_06040_),
    .X(_06062_));
 sky130_fd_sc_hd__nand2_1 _12878_ (.A(_06040_),
    .B(_06061_),
    .Y(_06063_));
 sky130_fd_sc_hd__nand2_1 _12879_ (.A(_06062_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__or2b_1 _12880_ (.A(_06058_),
    .B_N(_06064_),
    .X(_06066_));
 sky130_fd_sc_hd__or2b_1 _12881_ (.A(_06064_),
    .B_N(_06058_),
    .X(_06067_));
 sky130_fd_sc_hd__nand2_1 _12882_ (.A(_06066_),
    .B(_06067_),
    .Y(_06068_));
 sky130_fd_sc_hd__or2_1 _12883_ (.A(_06068_),
    .B(_06045_),
    .X(_06069_));
 sky130_fd_sc_hd__nand2_1 _12884_ (.A(_06045_),
    .B(_06068_),
    .Y(_06070_));
 sky130_fd_sc_hd__nand2_1 _12885_ (.A(_06069_),
    .B(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__nand2_1 _12886_ (.A(_06057_),
    .B(_06071_),
    .Y(_06072_));
 sky130_fd_sc_hd__inv_2 _12887_ (.A(_06071_),
    .Y(_06073_));
 sky130_fd_sc_hd__nand3_1 _12888_ (.A(_06055_),
    .B(_06056_),
    .C(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__nand2_1 _12889_ (.A(_06072_),
    .B(_06074_),
    .Y(\m1.out[46] ));
 sky130_fd_sc_hd__nand2_1 _12890_ (.A(_06057_),
    .B(_06073_),
    .Y(_06076_));
 sky130_fd_sc_hd__or3b_1 _12891_ (.A(_05995_),
    .B(_06059_),
    .C_N(_06038_),
    .X(_06077_));
 sky130_fd_sc_hd__and3b_1 _12892_ (.A_N(_06077_),
    .B(_06067_),
    .C(_06062_),
    .X(_06078_));
 sky130_fd_sc_hd__nand3_1 _12893_ (.A(_06076_),
    .B(_06069_),
    .C(_06078_),
    .Y(\m1.out[47] ));
 sky130_fd_sc_hd__and2_1 _12894_ (.A(_00256_),
    .B(_00095_),
    .X(_06079_));
 sky130_fd_sc_hd__nor2_1 _12895_ (.A(_00257_),
    .B(_06079_),
    .Y(\m1.out[8] ));
 sky130_fd_sc_hd__nand2_1 _12896_ (.A(_04378_),
    .B(net123),
    .Y(_06080_));
 sky130_fd_sc_hd__o21ai_1 _12897_ (.A1(_04378_),
    .A2(_01446_),
    .B1(net124),
    .Y(_00026_));
 sky130_fd_sc_hd__nand2_1 _12898_ (.A(net129),
    .B(net126),
    .Y(_06081_));
 sky130_fd_sc_hd__inv_2 _12899_ (.A(net127),
    .Y(_06082_));
 sky130_fd_sc_hd__a21o_1 _12900_ (.A1(net162),
    .A2(_03072_),
    .B1(_06082_),
    .X(_00017_));
 sky130_fd_sc_hd__o21ai_1 _12901_ (.A1(_04378_),
    .A2(_06124_),
    .B1(net127),
    .Y(_00018_));
 sky130_fd_sc_hd__a21o_1 _12902_ (.A1(net166),
    .A2(_03072_),
    .B1(_06082_),
    .X(_00019_));
 sky130_fd_sc_hd__a21o_1 _12903_ (.A1(net175),
    .A2(_03072_),
    .B1(_06082_),
    .X(_00020_));
 sky130_fd_sc_hd__o21ai_1 _12904_ (.A1(_04378_),
    .A2(net136),
    .B1(net127),
    .Y(_00021_));
 sky130_fd_sc_hd__o21ai_1 _12905_ (.A1(_02135_),
    .A2(_05904_),
    .B1(net127),
    .Y(_00022_));
 sky130_fd_sc_hd__o21ai_1 _12906_ (.A1(_02135_),
    .A2(net147),
    .B1(net127),
    .Y(_00023_));
 sky130_fd_sc_hd__a21o_1 _12907_ (.A1(_06158_),
    .A2(_03072_),
    .B1(_06082_),
    .X(_00025_));
 sky130_fd_sc_hd__nand2_1 _12908_ (.A(net157),
    .B(_02157_),
    .Y(_06084_));
 sky130_fd_sc_hd__inv_2 _12909_ (.A(_01555_),
    .Y(_06085_));
 sky130_fd_sc_hd__nor2_1 _12910_ (.A(_01336_),
    .B(_06085_),
    .Y(_06087_));
 sky130_fd_sc_hd__a21o_1 _12911_ (.A1(_04151_),
    .A2(_06084_),
    .B1(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__nand2_1 _12912_ (.A(_02157_),
    .B(_04151_),
    .Y(_06089_));
 sky130_fd_sc_hd__nand2_1 _12913_ (.A(_01555_),
    .B(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__and2_1 _12914_ (.A(_06090_),
    .B(net142),
    .X(_06091_));
 sky130_fd_sc_hd__a211o_1 _12915_ (.A1(_06088_),
    .A2(net141),
    .B1(net130),
    .C1(_06091_),
    .X(_06092_));
 sky130_fd_sc_hd__inv_2 _12916_ (.A(net181),
    .Y(_00002_));
 sky130_fd_sc_hd__nand2_1 _12917_ (.A(net204),
    .B(net141),
    .Y(_06093_));
 sky130_fd_sc_hd__nand2_1 _12918_ (.A(_01665_),
    .B(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__and3_1 _12919_ (.A(_04314_),
    .B(net204),
    .C(_04151_),
    .X(_06095_));
 sky130_fd_sc_hd__a221o_1 _12920_ (.A1(_06090_),
    .A2(_06094_),
    .B1(_06087_),
    .B2(net204),
    .C1(_06095_),
    .X(_06097_));
 sky130_fd_sc_hd__nor2_1 _12921_ (.A(_04378_),
    .B(_06097_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_1 _12922_ (.A(_02058_),
    .B(_05655_),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_1 _12923_ (.A(_01665_),
    .B(_01643_),
    .Y(_06099_));
 sky130_fd_sc_hd__nand2_1 _12924_ (.A(_01676_),
    .B(_06099_),
    .Y(_06100_));
 sky130_fd_sc_hd__a32o_1 _12925_ (.A1(_01533_),
    .A2(_06089_),
    .A3(_01643_),
    .B1(_06090_),
    .B2(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__a221o_1 _12926_ (.A1(net206),
    .A2(_06098_),
    .B1(_06101_),
    .B2(_05655_),
    .C1(net130),
    .X(_06102_));
 sky130_fd_sc_hd__inv_2 _12927_ (.A(_06102_),
    .Y(_00024_));
 sky130_fd_sc_hd__nand2_1 _12928_ (.A(_01676_),
    .B(net192),
    .Y(_06103_));
 sky130_fd_sc_hd__or2b_1 _12929_ (.A(_01686_),
    .B_N(_06103_),
    .X(_06104_));
 sky130_fd_sc_hd__a32o_1 _12930_ (.A1(_01533_),
    .A2(_06089_),
    .A3(net192),
    .B1(_06090_),
    .B2(_06104_),
    .X(_06106_));
 sky130_fd_sc_hd__a221o_1 _12931_ (.A1(_06098_),
    .A2(net192),
    .B1(_06106_),
    .B2(_05655_),
    .C1(net130),
    .X(_06107_));
 sky130_fd_sc_hd__inv_2 _12932_ (.A(net193),
    .Y(_00027_));
 sky130_fd_sc_hd__or2_1 _12933_ (.A(net273),
    .B(_01686_),
    .X(_06108_));
 sky130_fd_sc_hd__nand2_1 _12934_ (.A(_01686_),
    .B(net273),
    .Y(_06109_));
 sky130_fd_sc_hd__nand2_1 _12935_ (.A(_06108_),
    .B(net274),
    .Y(_06110_));
 sky130_fd_sc_hd__a2bb2o_1 _12936_ (.A1_N(net273),
    .A2_N(_01478_),
    .B1(_02036_),
    .B2(net275),
    .X(_06111_));
 sky130_fd_sc_hd__a221o_1 _12937_ (.A1(_01992_),
    .A2(net275),
    .B1(_01533_),
    .B2(_01741_),
    .C1(_06111_),
    .X(_06112_));
 sky130_fd_sc_hd__mux2_1 _12938_ (.A0(net275),
    .A1(_01741_),
    .S(_04314_),
    .X(_06113_));
 sky130_fd_sc_hd__and2_1 _12939_ (.A(_06113_),
    .B(_04151_),
    .X(_06114_));
 sky130_fd_sc_hd__a211o_1 _12940_ (.A1(net276),
    .A2(_02146_),
    .B1(net130),
    .C1(_06114_),
    .X(_06116_));
 sky130_fd_sc_hd__inv_2 _12941_ (.A(net277),
    .Y(_00028_));
 sky130_fd_sc_hd__nand2_1 _12942_ (.A(net274),
    .B(_01719_),
    .Y(_06117_));
 sky130_fd_sc_hd__nand2_1 _12943_ (.A(_06117_),
    .B(_02298_),
    .Y(_06118_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(_06118_),
    .A1(_01719_),
    .S(_04314_),
    .X(_06119_));
 sky130_fd_sc_hd__inv_2 _12945_ (.A(_06087_),
    .Y(_06120_));
 sky130_fd_sc_hd__nor2_1 _12946_ (.A(net284),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__a221o_1 _12947_ (.A1(_04151_),
    .A2(_06119_),
    .B1(_06085_),
    .B2(_06118_),
    .C1(net285),
    .X(_06122_));
 sky130_fd_sc_hd__nor2_1 _12948_ (.A(_04378_),
    .B(_06122_),
    .Y(_00029_));
 sky130_fd_sc_hd__nand2_1 _12949_ (.A(_02298_),
    .B(_01796_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _12950_ (.A(_02309_),
    .B(_06123_),
    .Y(_06125_));
 sky130_fd_sc_hd__mux2_1 _12951_ (.A0(_06125_),
    .A1(_01796_),
    .S(_04314_),
    .X(_06126_));
 sky130_fd_sc_hd__nor2_1 _12952_ (.A(net264),
    .B(_06120_),
    .Y(_06127_));
 sky130_fd_sc_hd__a221o_1 _12953_ (.A1(_04151_),
    .A2(_06126_),
    .B1(_06085_),
    .B2(_06125_),
    .C1(net265),
    .X(_06128_));
 sky130_fd_sc_hd__nor2_1 _12954_ (.A(_04378_),
    .B(net266),
    .Y(_00030_));
 sky130_fd_sc_hd__nand2_1 _12955_ (.A(_02309_),
    .B(net239),
    .Y(_06129_));
 sky130_fd_sc_hd__and2_1 _12956_ (.A(_02320_),
    .B(_06129_),
    .X(_06130_));
 sky130_fd_sc_hd__mux2_1 _12957_ (.A0(_06130_),
    .A1(net238),
    .S(_04314_),
    .X(_06131_));
 sky130_fd_sc_hd__or2_1 _12958_ (.A(_06130_),
    .B(_01555_),
    .X(_06132_));
 sky130_fd_sc_hd__nand2_1 _12959_ (.A(_06087_),
    .B(net239),
    .Y(_06133_));
 sky130_fd_sc_hd__o2111a_1 _12960_ (.A1(_02124_),
    .A2(_06131_),
    .B1(_03072_),
    .C1(_06132_),
    .D1(net240),
    .X(_00031_));
 sky130_fd_sc_hd__or2_1 _12961_ (.A(_01851_),
    .B(_01818_),
    .X(_06135_));
 sky130_fd_sc_hd__nand2_1 _12962_ (.A(_06135_),
    .B(_01862_),
    .Y(_06136_));
 sky130_fd_sc_hd__mux2_1 _12963_ (.A0(_06136_),
    .A1(_01840_),
    .S(_04314_),
    .X(_06137_));
 sky130_fd_sc_hd__nand2_1 _12964_ (.A(_06137_),
    .B(_04151_),
    .Y(_06138_));
 sky130_fd_sc_hd__nand2_1 _12965_ (.A(_06085_),
    .B(_06136_),
    .Y(_06139_));
 sky130_fd_sc_hd__o2111a_1 _12966_ (.A1(_01851_),
    .A2(_06120_),
    .B1(_03072_),
    .C1(_06138_),
    .D1(_06139_),
    .X(_00032_));
 sky130_fd_sc_hd__dfrtp_1 _12967_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00002_),
    .RESET_B(net109),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _12968_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00013_),
    .RESET_B(net109),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _12969_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00024_),
    .RESET_B(net109),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _12970_ (.CLK(clknet_3_5__leaf_clk),
    .D(net194),
    .RESET_B(net109),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _12971_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00028_),
    .RESET_B(net110),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _12972_ (.CLK(clknet_3_3__leaf_clk),
    .D(_00029_),
    .RESET_B(net110),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _12973_ (.CLK(clknet_3_3__leaf_clk),
    .D(net267),
    .RESET_B(net110),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _12974_ (.CLK(clknet_3_3__leaf_clk),
    .D(net241),
    .RESET_B(net110),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _12975_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00032_),
    .RESET_B(net110),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _12976_ (.CLK(clknet_3_5__leaf_clk),
    .D(net186),
    .RESET_B(net109),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _12977_ (.CLK(clknet_3_5__leaf_clk),
    .D(net236),
    .RESET_B(net109),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _12978_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00004_),
    .RESET_B(net109),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _12979_ (.CLK(clknet_3_5__leaf_clk),
    .D(_00005_),
    .RESET_B(net109),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _12980_ (.CLK(clknet_3_5__leaf_clk),
    .D(net213),
    .RESET_B(net109),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _12981_ (.CLK(clknet_3_5__leaf_clk),
    .D(net254),
    .RESET_B(net109),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _12982_ (.CLK(clknet_3_4__leaf_clk),
    .D(_00008_),
    .RESET_B(net110),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _12983_ (.CLK(clknet_3_4__leaf_clk),
    .D(_00009_),
    .RESET_B(net115),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _12984_ (.CLK(clknet_3_4__leaf_clk),
    .D(net224),
    .RESET_B(net115),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _12985_ (.CLK(clknet_3_4__leaf_clk),
    .D(_00011_),
    .RESET_B(net115),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _12986_ (.CLK(clknet_3_4__leaf_clk),
    .D(net247),
    .RESET_B(net115),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _12987_ (.CLK(clknet_3_7__leaf_clk),
    .D(_00014_),
    .RESET_B(net115),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _12988_ (.CLK(clknet_3_7__leaf_clk),
    .D(_00015_),
    .RESET_B(net115),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _12989_ (.CLK(clknet_3_7__leaf_clk),
    .D(net154),
    .RESET_B(net115),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _12990_ (.CLK(clknet_3_7__leaf_clk),
    .D(net163),
    .RESET_B(net115),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _12991_ (.CLK(clknet_3_7__leaf_clk),
    .D(net131),
    .RESET_B(net115),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _12992_ (.CLK(clknet_3_7__leaf_clk),
    .D(net167),
    .RESET_B(net115),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _12993_ (.CLK(clknet_3_7__leaf_clk),
    .D(net176),
    .RESET_B(net114),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _12994_ (.CLK(clknet_3_7__leaf_clk),
    .D(net137),
    .RESET_B(net114),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _12995_ (.CLK(clknet_3_7__leaf_clk),
    .D(net128),
    .RESET_B(net114),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _12996_ (.CLK(clknet_3_7__leaf_clk),
    .D(net148),
    .RESET_B(net114),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _12997_ (.CLK(clknet_3_6__leaf_clk),
    .D(_00025_),
    .RESET_B(net114),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _12998_ (.CLK(clknet_3_7__leaf_clk),
    .D(net125),
    .RESET_B(net114),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _12999_ (.CLK(clknet_3_7__leaf_clk),
    .D(_00034_),
    .RESET_B(net114),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _13000_ (.CLK(clknet_3_6__leaf_clk),
    .D(_00035_),
    .RESET_B(net114),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _13001_ (.CLK(clknet_3_7__leaf_clk),
    .D(net287),
    .RESET_B(net114),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _13002_ (.CLK(clknet_3_7__leaf_clk),
    .D(net122),
    .RESET_B(net114),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _13003_ (.CLK(clknet_3_7__leaf_clk),
    .D(_00000_),
    .RESET_B(net116),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _13004_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[0] ),
    .RESET_B(net106),
    .Q(\M000[0] ));
 sky130_fd_sc_hd__dfrtp_1 _13005_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[1] ),
    .RESET_B(net106),
    .Q(\M000[1] ));
 sky130_fd_sc_hd__dfrtp_1 _13006_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[2] ),
    .RESET_B(net106),
    .Q(\M000[2] ));
 sky130_fd_sc_hd__dfrtp_1 _13007_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[3] ),
    .RESET_B(net106),
    .Q(\M000[3] ));
 sky130_fd_sc_hd__dfrtp_1 _13008_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[4] ),
    .RESET_B(net107),
    .Q(\M000[4] ));
 sky130_fd_sc_hd__dfrtp_1 _13009_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[5] ),
    .RESET_B(net107),
    .Q(\M000[5] ));
 sky130_fd_sc_hd__dfrtp_1 _13010_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[6] ),
    .RESET_B(net107),
    .Q(\M000[6] ));
 sky130_fd_sc_hd__dfrtp_1 _13011_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[7] ),
    .RESET_B(net107),
    .Q(\M000[7] ));
 sky130_fd_sc_hd__dfrtp_1 _13012_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[8] ),
    .RESET_B(net107),
    .Q(\M000[8] ));
 sky130_fd_sc_hd__dfrtp_1 _13013_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[9] ),
    .RESET_B(net107),
    .Q(\M000[9] ));
 sky130_fd_sc_hd__dfrtp_1 _13014_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[10] ),
    .RESET_B(net106),
    .Q(\M000[10] ));
 sky130_fd_sc_hd__dfrtp_1 _13015_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[11] ),
    .RESET_B(net106),
    .Q(\M000[11] ));
 sky130_fd_sc_hd__dfrtp_1 _13016_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[12] ),
    .RESET_B(net106),
    .Q(\M000[12] ));
 sky130_fd_sc_hd__dfrtp_1 _13017_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[13] ),
    .RESET_B(net106),
    .Q(\M000[13] ));
 sky130_fd_sc_hd__dfrtp_1 _13018_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[14] ),
    .RESET_B(net106),
    .Q(\M000[14] ));
 sky130_fd_sc_hd__dfrtp_1 _13019_ (.CLK(clknet_3_0__leaf_clk),
    .D(\m1.out[15] ),
    .RESET_B(net106),
    .Q(\M000[15] ));
 sky130_fd_sc_hd__dfrtp_1 _13020_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[16] ),
    .RESET_B(net108),
    .Q(\M000[16] ));
 sky130_fd_sc_hd__dfrtp_1 _13021_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[17] ),
    .RESET_B(net108),
    .Q(\M000[17] ));
 sky130_fd_sc_hd__dfrtp_1 _13022_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[18] ),
    .RESET_B(net108),
    .Q(\M000[18] ));
 sky130_fd_sc_hd__dfrtp_1 _13023_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[19] ),
    .RESET_B(net108),
    .Q(\M000[19] ));
 sky130_fd_sc_hd__dfrtp_1 _13024_ (.CLK(clknet_3_3__leaf_clk),
    .D(\m1.out[20] ),
    .RESET_B(net108),
    .Q(\M000[20] ));
 sky130_fd_sc_hd__dfrtp_1 _13025_ (.CLK(clknet_3_1__leaf_clk),
    .D(\m1.out[21] ),
    .RESET_B(net108),
    .Q(\M000[21] ));
 sky130_fd_sc_hd__dfrtp_1 _13026_ (.CLK(clknet_3_3__leaf_clk),
    .D(\m1.out[22] ),
    .RESET_B(net111),
    .Q(\M000[22] ));
 sky130_fd_sc_hd__dfrtp_1 _13027_ (.CLK(clknet_3_3__leaf_clk),
    .D(\m1.out[23] ),
    .RESET_B(net111),
    .Q(\M000[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13028_ (.CLK(clknet_3_2__leaf_clk),
    .D(\m1.out[24] ),
    .RESET_B(net111),
    .Q(\M000[24] ));
 sky130_fd_sc_hd__dfrtp_1 _13029_ (.CLK(clknet_3_2__leaf_clk),
    .D(\m1.out[25] ),
    .RESET_B(net117),
    .Q(\M000[25] ));
 sky130_fd_sc_hd__dfrtp_1 _13030_ (.CLK(clknet_3_2__leaf_clk),
    .D(\m1.out[26] ),
    .RESET_B(net111),
    .Q(\M000[26] ));
 sky130_fd_sc_hd__dfrtp_1 _13031_ (.CLK(clknet_3_2__leaf_clk),
    .D(\m1.out[27] ),
    .RESET_B(net111),
    .Q(\M000[27] ));
 sky130_fd_sc_hd__dfrtp_1 _13032_ (.CLK(clknet_3_3__leaf_clk),
    .D(\m1.out[28] ),
    .RESET_B(net111),
    .Q(\M000[28] ));
 sky130_fd_sc_hd__dfrtp_1 _13033_ (.CLK(clknet_3_5__leaf_clk),
    .D(\m1.out[29] ),
    .RESET_B(net111),
    .Q(\M000[29] ));
 sky130_fd_sc_hd__dfrtp_1 _13034_ (.CLK(clknet_3_2__leaf_clk),
    .D(\m1.out[30] ),
    .RESET_B(net117),
    .Q(\M000[30] ));
 sky130_fd_sc_hd__dfrtp_1 _13035_ (.CLK(clknet_3_6__leaf_clk),
    .D(\m1.out[31] ),
    .RESET_B(net112),
    .Q(\M000[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13036_ (.CLK(clknet_3_7__leaf_clk),
    .D(\m1.out[32] ),
    .RESET_B(net113),
    .Q(\M000[32] ));
 sky130_fd_sc_hd__dfrtp_1 _13037_ (.CLK(clknet_3_6__leaf_clk),
    .D(\m1.out[33] ),
    .RESET_B(net112),
    .Q(\M000[33] ));
 sky130_fd_sc_hd__dfrtp_1 _13038_ (.CLK(clknet_3_6__leaf_clk),
    .D(\m1.out[34] ),
    .RESET_B(net112),
    .Q(\M000[34] ));
 sky130_fd_sc_hd__dfrtp_1 _13039_ (.CLK(clknet_3_6__leaf_clk),
    .D(\m1.out[35] ),
    .RESET_B(net112),
    .Q(\M000[35] ));
 sky130_fd_sc_hd__dfrtp_1 _13040_ (.CLK(clknet_3_6__leaf_clk),
    .D(\m1.out[36] ),
    .RESET_B(net112),
    .Q(\M000[36] ));
 sky130_fd_sc_hd__dfrtp_1 _13041_ (.CLK(clknet_3_7__leaf_clk),
    .D(\m1.out[37] ),
    .RESET_B(net113),
    .Q(\M000[37] ));
 sky130_fd_sc_hd__dfrtp_1 _13042_ (.CLK(clknet_3_6__leaf_clk),
    .D(\m1.out[38] ),
    .RESET_B(net112),
    .Q(\M000[38] ));
 sky130_fd_sc_hd__dfrtp_1 _13043_ (.CLK(clknet_3_6__leaf_clk),
    .D(\m1.out[39] ),
    .RESET_B(net112),
    .Q(\M000[39] ));
 sky130_fd_sc_hd__dfrtp_1 _13044_ (.CLK(clknet_3_7__leaf_clk),
    .D(\m1.out[40] ),
    .RESET_B(net113),
    .Q(\M000[40] ));
 sky130_fd_sc_hd__dfrtp_1 _13045_ (.CLK(clknet_3_4__leaf_clk),
    .D(\m1.out[41] ),
    .RESET_B(net113),
    .Q(\M000[41] ));
 sky130_fd_sc_hd__dfrtp_1 _13046_ (.CLK(clknet_3_4__leaf_clk),
    .D(\m1.out[42] ),
    .RESET_B(net113),
    .Q(\M000[42] ));
 sky130_fd_sc_hd__dfrtp_1 _13047_ (.CLK(clknet_3_4__leaf_clk),
    .D(\m1.out[43] ),
    .RESET_B(net113),
    .Q(\M000[43] ));
 sky130_fd_sc_hd__dfrtp_1 _13048_ (.CLK(clknet_3_4__leaf_clk),
    .D(\m1.out[44] ),
    .RESET_B(net113),
    .Q(\M000[44] ));
 sky130_fd_sc_hd__dfrtp_1 _13049_ (.CLK(clknet_3_5__leaf_clk),
    .D(\m1.out[45] ),
    .RESET_B(net113),
    .Q(\M000[45] ));
 sky130_fd_sc_hd__dfrtp_1 _13050_ (.CLK(clknet_3_5__leaf_clk),
    .D(\m1.out[46] ),
    .RESET_B(net111),
    .Q(\M000[46] ));
 sky130_fd_sc_hd__dfrtp_1 _13051_ (.CLK(clknet_3_2__leaf_clk),
    .D(\m1.out[47] ),
    .RESET_B(net111),
    .Q(\M000[47] ));
 sky130_fd_sc_hd__dfrtp_1 _13052_ (.CLK(clknet_3_6__leaf_clk),
    .D(net118),
    .RESET_B(net116),
    .Q(done0_reg));
 sky130_fd_sc_hd__conb_1 _13052__118 (.HI(net118));
 sky130_fd_sc_hd__dfrtp_1 _13053_ (.CLK(clknet_3_7__leaf_clk),
    .D(inv_f_c),
    .RESET_B(net112),
    .Q(inv_f));
 sky130_fd_sc_hd__dfrtp_1 _13054_ (.CLK(clknet_3_6__leaf_clk),
    .D(\out_f_c[23] ),
    .RESET_B(net112),
    .Q(\out_f[23] ));
 sky130_fd_sc_hd__dfrtp_1 _13055_ (.CLK(clknet_3_6__leaf_clk),
    .D(\out_f_c[31] ),
    .RESET_B(net113),
    .Q(\out_f[31] ));
 sky130_fd_sc_hd__dfrtp_1 _13056_ (.CLK(clknet_3_6__leaf_clk),
    .D(forward_c),
    .RESET_B(net112),
    .Q(forward));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(net108),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net117),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net117),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net116),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(net116),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net68),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net286),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00022_),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_04173_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\M000[40] ),
    .X(net219));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold102 (.A(_03333_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_03454_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_03465_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_03476_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_00010_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\M000[34] ),
    .X(net225));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold108 (.A(_02254_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_02408_),
    .X(net227));
 sky130_fd_sc_hd__buf_1 hold11 (.A(net187),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_02418_),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_02429_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_02440_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\M000[33] ),
    .X(net231));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold114 (.A(_01915_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_02200_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_02211_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_02222_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_00003_),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\M000[30] ),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 hold12 (.A(_01588_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_01763_),
    .X(net238));
 sky130_fd_sc_hd__buf_1 hold121 (.A(_01774_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_06133_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_00031_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\M000[42] ),
    .X(net242));
 sky130_fd_sc_hd__buf_1 hold125 (.A(_03682_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_03813_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_03824_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_03835_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_00012_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_00018_),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\M000[37] ),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 hold131 (.A(_02810_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_02920_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_02931_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_02942_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_02953_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_00007_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\M000[39] ),
    .X(net255));
 sky130_fd_sc_hd__buf_1 hold138 (.A(_03148_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_03529_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\M000[22] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\M000[35] ),
    .X(net258));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold141 (.A(_02461_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_02593_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_02604_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_02615_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\M000[29] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_01785_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_06127_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_06128_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_00030_),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 hold15 (.A(_01369_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\M000[38] ),
    .X(net268));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold151 (.A(_02984_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_03170_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_03181_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\M000[27] ),
    .X(net272));
 sky130_fd_sc_hd__buf_1 hold155 (.A(_01730_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_06109_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_06110_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_06112_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_06116_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_05731_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\M000[31] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_01829_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_02331_),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_03039_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_03061_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\M000[28] ),
    .X(net283));
 sky130_fd_sc_hd__buf_1 hold166 (.A(_01708_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_06121_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net288),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net119),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_05742_),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(done0_reg),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_05818_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_00021_),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(inv_f),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\M000[24] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_01172_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_01183_),
    .X(net140));
 sky130_fd_sc_hd__buf_1 hold23 (.A(net180),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_01205_),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_01380_),
    .X(net143));
 sky130_fd_sc_hd__buf_1 hold26 (.A(_01391_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_2 hold27 (.A(_01566_),
    .X(net145));
 sky130_fd_sc_hd__buf_1 hold28 (.A(_01577_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_05687_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_04347_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00023_),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\M000[46] ),
    .X(net149));
 sky130_fd_sc_hd__buf_1 hold32 (.A(_04205_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_04270_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_04281_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_04303_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_00016_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\M000[21] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_01227_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_2 hold39 (.A(_01292_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00001_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 hold40 (.A(_01402_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_06044_),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_06054_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_06065_),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_06165_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_00017_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 hold46 (.A(net205),
    .X(net164));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold47 (.A(_01117_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_05958_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_00019_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\out_f[31] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\M000[43] ),
    .X(net168));
 sky130_fd_sc_hd__buf_1 hold51 (.A(_03856_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_03867_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_04913_),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_04956_),
    .X(net172));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold55 (.A(_04967_),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_05044_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_05098_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_00020_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\out_f[23] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_06080_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_06081_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\M000[23] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_01194_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_06092_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\M000[32] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_01139_),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_01150_),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 hold67 (.A(_01161_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_00033_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(forward),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_00026_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net129),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\M000[26] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_01599_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_01610_),
    .X(net191));
 sky130_fd_sc_hd__buf_1 hold74 (.A(_01621_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_06107_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_00027_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\M000[41] ),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 hold78 (.A(_03496_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_03878_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net177),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_03889_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_03987_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_03998_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_04009_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\M000[25] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_01632_),
    .X(net203));
 sky130_fd_sc_hd__buf_1 hold86 (.A(_01654_),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\M000[47] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_01643_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\M000[36] ),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 hold9 (.A(net178),
    .X(net127));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold90 (.A(_02647_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_02756_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_02767_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_02778_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_02789_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_00006_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\M000[44] ),
    .X(net214));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold97 (.A(_04052_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_04074_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_04085_),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(in1[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(in1[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(in1[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(in1[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_8 input13 (.A(in1[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(in1[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input15 (.A(in1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in1[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(in1[24]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(in1[25]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(in1[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_4 input2 (.A(in1[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in1[27]),
    .X(net20));
 sky130_fd_sc_hd__dlymetal6s2s_1 input21 (.A(in1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in1[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(in1[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in1[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(in1[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(in1[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(in1[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(in1[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 input29 (.A(in1[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(in1[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(in1[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(in1[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(in1[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(in2[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(in2[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(in2[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(in2[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(in2[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_4 input38 (.A(in2[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_4 input39 (.A(in2[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_8 input4 (.A(in1[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(in2[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 input41 (.A(in2[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(in2[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(in2[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input44 (.A(in2[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(in2[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 input46 (.A(in2[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_4 input47 (.A(in2[22]),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(in2[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(in2[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(in1[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(in2[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(in2[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(in2[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(in2[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(in2[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(in2[2]),
    .X(net55));
 sky130_fd_sc_hd__dlymetal6s2s_1 input56 (.A(in2[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(in2[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(in2[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(in2[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(in1[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input60 (.A(in2[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 input61 (.A(in2[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(in2[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_4 input63 (.A(in2[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_4 input64 (.A(in2[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_4 input65 (.A(round_m[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 input66 (.A(round_m[1]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(round_m[2]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(rst),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input7 (.A(in1[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(in1[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(in1[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(out[6]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(out[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(out[8]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(out[9]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(ov));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(un));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(done));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(inexact));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(inv));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(out[0]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(out[10]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(out[11]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(out[12]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(out[13]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(out[14]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(out[15]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(out[16]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(out[17]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(out[18]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(out[19]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(out[20]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(out[21]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(out[22]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(out[23]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(out[24]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(out[25]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(out[26]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(out[27]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(out[28]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(out[29]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(out[2]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(out[30]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(out[31]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(out[3]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(out[4]));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net99),
    .X(out[5]));
endmodule

