// This is the unpowered netlist.
module fp_comp (act,
    clk,
    done,
    eq,
    great,
    inv,
    less,
    rst,
    in1,
    in2);
 input act;
 input clk;
 output done;
 output eq;
 output great;
 output inv;
 output less;
 input rst;
 input [31:0] in1;
 input [31:0] in2;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire eq_f;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA__362__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__363__B (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__367__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__368__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__375__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__378__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__379__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__384__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__389__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__390__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__392__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__394__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__406__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__410__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__413__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__441__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__441__C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__442__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__442__C (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__443__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__443__D (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__444__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__444__C (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__447__C_N (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__448__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__448__B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__449__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__449__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__449__C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__449__D (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__461__RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__462__RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__463__RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__464__RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__465__RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__466__RESET_B (.DIODE(net65));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_96 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _231_ (.A(net12),
    .Y(_201_));
 sky130_fd_sc_hd__nand2_1 _232_ (.A(_201_),
    .B(net44),
    .Y(_202_));
 sky130_fd_sc_hd__inv_2 _233_ (.A(net44),
    .Y(_203_));
 sky130_fd_sc_hd__nand2_1 _234_ (.A(_203_),
    .B(net12),
    .Y(_204_));
 sky130_fd_sc_hd__inv_2 _235_ (.A(net33),
    .Y(_205_));
 sky130_fd_sc_hd__nand2_1 _236_ (.A(_205_),
    .B(net1),
    .Y(_206_));
 sky130_fd_sc_hd__nand3_1 _237_ (.A(_202_),
    .B(_204_),
    .C(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__nand2_1 _238_ (.A(_207_),
    .B(_202_),
    .Y(_208_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(net26),
    .Y(_209_));
 sky130_fd_sc_hd__nand2_1 _240_ (.A(_209_),
    .B(net58),
    .Y(_210_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(net58),
    .Y(_211_));
 sky130_fd_sc_hd__nand2_1 _242_ (.A(_211_),
    .B(net26),
    .Y(_212_));
 sky130_fd_sc_hd__nand2_1 _243_ (.A(_210_),
    .B(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__nand2b_1 _244_ (.A_N(net55),
    .B(net23),
    .Y(_214_));
 sky130_fd_sc_hd__nand2b_1 _245_ (.A_N(net23),
    .B(net55),
    .Y(_215_));
 sky130_fd_sc_hd__nand2_1 _246_ (.A(_214_),
    .B(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__nor2_1 _247_ (.A(_213_),
    .B(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__nand2_1 _248_ (.A(_208_),
    .B(_217_),
    .Y(_218_));
 sky130_fd_sc_hd__nor2_1 _249_ (.A(net26),
    .B(_211_),
    .Y(_219_));
 sky130_fd_sc_hd__nor2_1 _250_ (.A(_215_),
    .B(_213_),
    .Y(_220_));
 sky130_fd_sc_hd__nor2_1 _251_ (.A(_219_),
    .B(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__nand2_1 _252_ (.A(_218_),
    .B(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(net30),
    .Y(_223_));
 sky130_fd_sc_hd__inv_2 _254_ (.A(net62),
    .Y(_224_));
 sky130_fd_sc_hd__nand2_1 _255_ (.A(_223_),
    .B(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__nand2_1 _256_ (.A(net30),
    .B(net62),
    .Y(_226_));
 sky130_fd_sc_hd__nand2_1 _257_ (.A(_225_),
    .B(_226_),
    .Y(_227_));
 sky130_fd_sc_hd__nand2b_1 _258_ (.A_N(net61),
    .B(net29),
    .Y(_228_));
 sky130_fd_sc_hd__nand2b_1 _259_ (.A_N(net29),
    .B(net61),
    .Y(_229_));
 sky130_fd_sc_hd__nand3_1 _260_ (.A(_227_),
    .B(_228_),
    .C(_229_),
    .Y(_004_));
 sky130_fd_sc_hd__xnor2_1 _261_ (.A(net28),
    .B(net60),
    .Y(_005_));
 sky130_fd_sc_hd__nand2b_1 _262_ (.A_N(net27),
    .B(net59),
    .Y(_006_));
 sky130_fd_sc_hd__nand2b_1 _263_ (.A_N(net59),
    .B(net27),
    .Y(_007_));
 sky130_fd_sc_hd__nand3_1 _264_ (.A(_005_),
    .B(_006_),
    .C(_007_),
    .Y(_008_));
 sky130_fd_sc_hd__nor2_1 _265_ (.A(_004_),
    .B(_008_),
    .Y(_009_));
 sky130_fd_sc_hd__nand2_1 _266_ (.A(_222_),
    .B(_009_),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _267_ (.A(net28),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_1 _268_ (.A(net60),
    .B(_011_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _269_ (.A(_011_),
    .B(net60),
    .Y(_013_));
 sky130_fd_sc_hd__o21ai_1 _270_ (.A1(_012_),
    .A2(_006_),
    .B1(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__nand2_1 _271_ (.A(_223_),
    .B(net62),
    .Y(_015_));
 sky130_fd_sc_hd__nand2_1 _272_ (.A(_224_),
    .B(net30),
    .Y(_016_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(_015_),
    .B(_016_),
    .Y(_017_));
 sky130_fd_sc_hd__nand2_1 _274_ (.A(_228_),
    .B(_229_),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _275_ (.A(_017_),
    .B(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__o21ai_1 _276_ (.A1(_229_),
    .A2(_017_),
    .B1(_015_),
    .Y(_020_));
 sky130_fd_sc_hd__a21oi_1 _277_ (.A1(_014_),
    .A2(_019_),
    .B1(_020_),
    .Y(_021_));
 sky130_fd_sc_hd__nand2_1 _278_ (.A(_010_),
    .B(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__nand2b_1 _279_ (.A_N(net3),
    .B(net35),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _280_ (.A(net35),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _281_ (.A(_024_),
    .B(net3),
    .Y(_025_));
 sky130_fd_sc_hd__nand2_1 _282_ (.A(_023_),
    .B(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__nand2b_1 _283_ (.A_N(net34),
    .B(net2),
    .Y(_027_));
 sky130_fd_sc_hd__nand2b_1 _284_ (.A_N(net2),
    .B(net34),
    .Y(_028_));
 sky130_fd_sc_hd__nand2_1 _285_ (.A(_027_),
    .B(_028_),
    .Y(_029_));
 sky130_fd_sc_hd__nor2_1 _286_ (.A(_026_),
    .B(_029_),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _287_ (.A(net32),
    .Y(_031_));
 sky130_fd_sc_hd__nor2_1 _288_ (.A(net64),
    .B(_031_),
    .Y(_032_));
 sky130_fd_sc_hd__nand2_1 _289_ (.A(_031_),
    .B(net64),
    .Y(_033_));
 sky130_fd_sc_hd__and2b_1 _290_ (.A_N(_032_),
    .B(_033_),
    .X(_034_));
 sky130_fd_sc_hd__xnor2_1 _291_ (.A(net63),
    .B(net31),
    .Y(_035_));
 sky130_fd_sc_hd__nand3_1 _292_ (.A(_030_),
    .B(_034_),
    .C(_035_),
    .Y(_036_));
 sky130_fd_sc_hd__nand2b_1 _293_ (.A_N(net6),
    .B(net38),
    .Y(_037_));
 sky130_fd_sc_hd__nand2b_1 _294_ (.A_N(net38),
    .B(net6),
    .Y(_038_));
 sky130_fd_sc_hd__nand2_1 _295_ (.A(_037_),
    .B(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__xnor2_1 _296_ (.A(net7),
    .B(net39),
    .Y(_040_));
 sky130_fd_sc_hd__nor2b_1 _297_ (.A(_039_),
    .B_N(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__xnor2_1 _298_ (.A(net36),
    .B(net4),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _299_ (.A(net5),
    .Y(_043_));
 sky130_fd_sc_hd__nor2_1 _300_ (.A(net37),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__and2_1 _301_ (.A(_043_),
    .B(net37),
    .X(_045_));
 sky130_fd_sc_hd__nor2_1 _302_ (.A(_044_),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__nand3_1 _303_ (.A(_041_),
    .B(_042_),
    .C(_046_),
    .Y(_047_));
 sky130_fd_sc_hd__nor2_1 _304_ (.A(_036_),
    .B(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_1 _305_ (.A(_022_),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__nand2b_1 _306_ (.A_N(net31),
    .B(net63),
    .Y(_050_));
 sky130_fd_sc_hd__o21ai_1 _307_ (.A1(_032_),
    .A2(_050_),
    .B1(_033_),
    .Y(_051_));
 sky130_fd_sc_hd__nand2_1 _308_ (.A(_051_),
    .B(_030_),
    .Y(_052_));
 sky130_fd_sc_hd__nor2_1 _309_ (.A(net3),
    .B(_024_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _310_ (.A(_028_),
    .B(_026_),
    .Y(_054_));
 sky130_fd_sc_hd__nor2_1 _311_ (.A(_053_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__nand2_1 _312_ (.A(_052_),
    .B(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__nand2_1 _313_ (.A(_046_),
    .B(_042_),
    .Y(_057_));
 sky130_fd_sc_hd__nand2b_1 _314_ (.A_N(_039_),
    .B(_040_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _315_ (.A(_057_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__nand2b_1 _316_ (.A_N(net4),
    .B(net36),
    .Y(_060_));
 sky130_fd_sc_hd__o21bai_1 _317_ (.A1(_044_),
    .A2(_060_),
    .B1_N(_045_),
    .Y(_061_));
 sky130_fd_sc_hd__nand2_1 _318_ (.A(_041_),
    .B(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _319_ (.A(net7),
    .Y(_063_));
 sky130_fd_sc_hd__nor2_1 _320_ (.A(net39),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__nand2_1 _321_ (.A(_063_),
    .B(net39),
    .Y(_065_));
 sky130_fd_sc_hd__o21a_1 _322_ (.A1(_064_),
    .A2(_037_),
    .B1(_065_),
    .X(_066_));
 sky130_fd_sc_hd__nand2_1 _323_ (.A(_062_),
    .B(_066_),
    .Y(_067_));
 sky130_fd_sc_hd__a21oi_1 _324_ (.A1(_056_),
    .A2(_059_),
    .B1(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__nand2_1 _325_ (.A(_049_),
    .B(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _326_ (.A(net41),
    .Y(_070_));
 sky130_fd_sc_hd__nor2_1 _327_ (.A(net9),
    .B(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__nand2_1 _328_ (.A(_070_),
    .B(net9),
    .Y(_072_));
 sky130_fd_sc_hd__and2b_1 _329_ (.A_N(_071_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__inv_2 _330_ (.A(net8),
    .Y(_074_));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(_074_),
    .B(net40),
    .Y(_075_));
 sky130_fd_sc_hd__or2_1 _332_ (.A(net40),
    .B(_074_),
    .X(_076_));
 sky130_fd_sc_hd__and3_1 _333_ (.A(_073_),
    .B(_075_),
    .C(_076_),
    .X(_077_));
 sky130_fd_sc_hd__or2_1 _334_ (.A(net11),
    .B(net43),
    .X(_078_));
 sky130_fd_sc_hd__nand2_1 _335_ (.A(net11),
    .B(net43),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_1 _336_ (.A(_078_),
    .B(_079_),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _337_ (.A(net10),
    .Y(_081_));
 sky130_fd_sc_hd__or2_1 _338_ (.A(net42),
    .B(_081_),
    .X(_082_));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(_081_),
    .B(net42),
    .Y(_083_));
 sky130_fd_sc_hd__and3_1 _340_ (.A(_080_),
    .B(_082_),
    .C(_083_),
    .X(_084_));
 sky130_fd_sc_hd__and2_1 _341_ (.A(_077_),
    .B(_084_),
    .X(_085_));
 sky130_fd_sc_hd__nand2_1 _342_ (.A(_069_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__a31o_1 _343_ (.A1(_072_),
    .A2(net40),
    .A3(_074_),
    .B1(_071_),
    .X(_087_));
 sky130_fd_sc_hd__inv_2 _344_ (.A(net43),
    .Y(_088_));
 sky130_fd_sc_hd__nor2_1 _345_ (.A(net11),
    .B(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__a31o_1 _346_ (.A1(_080_),
    .A2(_081_),
    .A3(net42),
    .B1(_089_),
    .X(_090_));
 sky130_fd_sc_hd__a21oi_1 _347_ (.A1(_087_),
    .A2(_084_),
    .B1(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(_086_),
    .B(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _349_ (.A(net13),
    .Y(_093_));
 sky130_fd_sc_hd__nor2_1 _350_ (.A(net45),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _351_ (.A(net45),
    .Y(_095_));
 sky130_fd_sc_hd__nor2_1 _352_ (.A(net13),
    .B(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_2 _353_ (.A(net46),
    .Y(_097_));
 sky130_fd_sc_hd__nor2_1 _354_ (.A(net14),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__nand2_1 _355_ (.A(_097_),
    .B(net14),
    .Y(_099_));
 sky130_fd_sc_hd__nand2b_1 _356_ (.A_N(_098_),
    .B(_099_),
    .Y(_100_));
 sky130_fd_sc_hd__nor3_1 _357_ (.A(_094_),
    .B(_096_),
    .C(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__nand2_1 _358_ (.A(_092_),
    .B(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__a21oi_1 _359_ (.A1(_096_),
    .A2(_099_),
    .B1(_098_),
    .Y(_103_));
 sky130_fd_sc_hd__nand2_1 _360_ (.A(_102_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__inv_2 _361_ (.A(net47),
    .Y(_105_));
 sky130_fd_sc_hd__or2_1 _362_ (.A(net15),
    .B(_105_),
    .X(_106_));
 sky130_fd_sc_hd__nand2_1 _363_ (.A(_105_),
    .B(net15),
    .Y(_107_));
 sky130_fd_sc_hd__and2_1 _364_ (.A(_106_),
    .B(_107_),
    .X(_108_));
 sky130_fd_sc_hd__nand2_1 _365_ (.A(_104_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__inv_2 _366_ (.A(net54),
    .Y(_110_));
 sky130_fd_sc_hd__nor2_1 _367_ (.A(net22),
    .B(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__and2_1 _368_ (.A(_110_),
    .B(net22),
    .X(_112_));
 sky130_fd_sc_hd__inv_2 _369_ (.A(net24),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(_113_),
    .B(net56),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _371_ (.A(net56),
    .Y(_115_));
 sky130_fd_sc_hd__nand2_1 _372_ (.A(_115_),
    .B(net24),
    .Y(_116_));
 sky130_fd_sc_hd__nand2_1 _373_ (.A(_114_),
    .B(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__or3_1 _374_ (.A(_111_),
    .B(_112_),
    .C(_117_),
    .X(_118_));
 sky130_fd_sc_hd__inv_2 _375_ (.A(net20),
    .Y(_119_));
 sky130_fd_sc_hd__nor2_1 _376_ (.A(net52),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__inv_2 _377_ (.A(net53),
    .Y(_121_));
 sky130_fd_sc_hd__or2_1 _378_ (.A(net21),
    .B(_121_),
    .X(_122_));
 sky130_fd_sc_hd__nand2_1 _379_ (.A(_121_),
    .B(net21),
    .Y(_123_));
 sky130_fd_sc_hd__nand2_1 _380_ (.A(_122_),
    .B(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2_1 _381_ (.A(_119_),
    .B(net52),
    .Y(_125_));
 sky130_fd_sc_hd__or3b_1 _382_ (.A(_120_),
    .B(_124_),
    .C_N(_125_),
    .X(_126_));
 sky130_fd_sc_hd__nor2_1 _383_ (.A(_118_),
    .B(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__inv_2 _384_ (.A(net19),
    .Y(_128_));
 sky130_fd_sc_hd__nor2_1 _385_ (.A(net51),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__nand2_1 _386_ (.A(_128_),
    .B(net51),
    .Y(_130_));
 sky130_fd_sc_hd__nor2b_1 _387_ (.A(_129_),
    .B_N(_130_),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(net50),
    .Y(_132_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(_132_),
    .B(net18),
    .Y(_133_));
 sky130_fd_sc_hd__or2_1 _390_ (.A(net18),
    .B(_132_),
    .X(_134_));
 sky130_fd_sc_hd__and3_1 _391_ (.A(_131_),
    .B(_133_),
    .C(_134_),
    .X(_135_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(net17),
    .Y(_136_));
 sky130_fd_sc_hd__nor2_1 _393_ (.A(net49),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(net16),
    .Y(_138_));
 sky130_fd_sc_hd__nor2_1 _395_ (.A(net48),
    .B(_138_),
    .Y(_139_));
 sky130_fd_sc_hd__nand2_1 _396_ (.A(_138_),
    .B(net48),
    .Y(_140_));
 sky130_fd_sc_hd__nor2b_1 _397_ (.A(_139_),
    .B_N(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__nand2_1 _398_ (.A(_136_),
    .B(net49),
    .Y(_142_));
 sky130_fd_sc_hd__and3b_1 _399_ (.A_N(_137_),
    .B(_141_),
    .C(_142_),
    .X(_143_));
 sky130_fd_sc_hd__and3_1 _400_ (.A(_127_),
    .B(_135_),
    .C(_143_),
    .X(_144_));
 sky130_fd_sc_hd__nand3_1 _401_ (.A(_109_),
    .B(_106_),
    .C(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__o21ai_1 _402_ (.A1(_137_),
    .A2(_139_),
    .B1(_142_),
    .Y(_146_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(_135_),
    .B(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__o211ai_1 _404_ (.A1(_129_),
    .A2(_134_),
    .B1(_130_),
    .C1(_147_),
    .Y(_148_));
 sky130_fd_sc_hd__o21a_1 _405_ (.A1(_125_),
    .A2(_124_),
    .B1(_122_),
    .X(_149_));
 sky130_fd_sc_hd__or3_1 _406_ (.A(net22),
    .B(_110_),
    .C(_117_),
    .X(_150_));
 sky130_fd_sc_hd__o211a_1 _407_ (.A1(_149_),
    .A2(_118_),
    .B1(_114_),
    .C1(_150_),
    .X(_151_));
 sky130_fd_sc_hd__a21bo_1 _408_ (.A1(_127_),
    .A2(_148_),
    .B1_N(_151_),
    .X(_152_));
 sky130_fd_sc_hd__nand2_1 _409_ (.A(_145_),
    .B(_152_),
    .Y(_153_));
 sky130_fd_sc_hd__xor2_2 _410_ (.A(net25),
    .B(net57),
    .X(_154_));
 sky130_fd_sc_hd__inv_2 _411_ (.A(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__nand2_1 _412_ (.A(_153_),
    .B(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__or2b_1 _413_ (.A(net25),
    .B_N(net57),
    .X(_157_));
 sky130_fd_sc_hd__a21oi_1 _414_ (.A1(_156_),
    .A2(_157_),
    .B1(net76),
    .Y(_002_));
 sky130_fd_sc_hd__o211a_1 _415_ (.A1(net1),
    .A2(_205_),
    .B1(_108_),
    .C1(_101_),
    .X(_158_));
 sky130_fd_sc_hd__and3b_1 _416_ (.A_N(_207_),
    .B(_158_),
    .C(_217_),
    .X(_159_));
 sky130_fd_sc_hd__and3_1 _417_ (.A(_077_),
    .B(_084_),
    .C(_009_),
    .X(_160_));
 sky130_fd_sc_hd__nand3_1 _418_ (.A(_159_),
    .B(_048_),
    .C(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__or3b_1 _419_ (.A(net72),
    .B(_154_),
    .C_N(_144_),
    .X(_162_));
 sky130_fd_sc_hd__o2bb2ai_1 _420_ (.A1_N(net72),
    .A2_N(net73),
    .B1(_161_),
    .B2(_162_),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_1 _421_ (.A(_109_),
    .B(_106_),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(_163_),
    .B(_161_),
    .Y(_164_));
 sky130_fd_sc_hd__nand2_1 _423_ (.A(_164_),
    .B(_144_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _424_ (.A(_165_),
    .B(_152_),
    .Y(_166_));
 sky130_fd_sc_hd__or2b_1 _425_ (.A(net76),
    .B_N(_157_),
    .X(_167_));
 sky130_fd_sc_hd__a21oi_1 _426_ (.A1(_166_),
    .A2(_155_),
    .B1(_167_),
    .Y(_003_));
 sky130_fd_sc_hd__or3_1 _427_ (.A(net29),
    .B(net61),
    .C(_225_),
    .X(_168_));
 sky130_fd_sc_hd__or4_1 _428_ (.A(net32),
    .B(net64),
    .C(net63),
    .D(net31),
    .X(_169_));
 sky130_fd_sc_hd__or4_1 _429_ (.A(net3),
    .B(net35),
    .C(net2),
    .D(net34),
    .X(_170_));
 sky130_fd_sc_hd__or4_1 _430_ (.A(net28),
    .B(net60),
    .C(net59),
    .D(net27),
    .X(_171_));
 sky130_fd_sc_hd__or4_1 _431_ (.A(_168_),
    .B(_169_),
    .C(_170_),
    .D(_171_),
    .X(_172_));
 sky130_fd_sc_hd__or3_1 _432_ (.A(net10),
    .B(net42),
    .C(_078_),
    .X(_173_));
 sky130_fd_sc_hd__or4_1 _433_ (.A(net9),
    .B(net41),
    .C(net40),
    .D(net8),
    .X(_174_));
 sky130_fd_sc_hd__or4_1 _434_ (.A(net5),
    .B(net37),
    .C(net36),
    .D(net4),
    .X(_175_));
 sky130_fd_sc_hd__or4_1 _435_ (.A(net7),
    .B(net39),
    .C(net6),
    .D(net38),
    .X(_176_));
 sky130_fd_sc_hd__or4_1 _436_ (.A(_173_),
    .B(_174_),
    .C(_175_),
    .D(_176_),
    .X(_177_));
 sky130_fd_sc_hd__nor2_1 _437_ (.A(_172_),
    .B(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__nand2_1 _438_ (.A(_097_),
    .B(_095_),
    .Y(_179_));
 sky130_fd_sc_hd__or2_1 _439_ (.A(net14),
    .B(net13),
    .X(_180_));
 sky130_fd_sc_hd__or4_1 _440_ (.A(net56),
    .B(net24),
    .C(_179_),
    .D(_180_),
    .X(_181_));
 sky130_fd_sc_hd__or4_1 _441_ (.A(net52),
    .B(net20),
    .C(net19),
    .D(net51),
    .X(_182_));
 sky130_fd_sc_hd__or4_1 _442_ (.A(net22),
    .B(net54),
    .C(net21),
    .D(net53),
    .X(_183_));
 sky130_fd_sc_hd__or4_1 _443_ (.A(net48),
    .B(net16),
    .C(net47),
    .D(net15),
    .X(_184_));
 sky130_fd_sc_hd__or4_1 _444_ (.A(net18),
    .B(net50),
    .C(net17),
    .D(net49),
    .X(_185_));
 sky130_fd_sc_hd__or4_1 _445_ (.A(_182_),
    .B(_183_),
    .C(_184_),
    .D(_185_),
    .X(_186_));
 sky130_fd_sc_hd__nor2_1 _446_ (.A(_181_),
    .B(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__or3b_1 _447_ (.A(_113_),
    .B(_180_),
    .C_N(net22),
    .X(_188_));
 sky130_fd_sc_hd__or4_1 _448_ (.A(net15),
    .B(net25),
    .C(_136_),
    .D(_138_),
    .X(_189_));
 sky130_fd_sc_hd__and4_1 _449_ (.A(net21),
    .B(net20),
    .C(net19),
    .D(net18),
    .X(_190_));
 sky130_fd_sc_hd__or3b_1 _450_ (.A(_188_),
    .B(_189_),
    .C_N(_190_),
    .X(_191_));
 sky130_fd_sc_hd__and4b_1 _451_ (.A_N(net57),
    .B(net49),
    .C(_105_),
    .D(net48),
    .X(_192_));
 sky130_fd_sc_hd__and4_1 _452_ (.A(net53),
    .B(net52),
    .C(net51),
    .D(net50),
    .X(_193_));
 sky130_fd_sc_hd__nor3_1 _453_ (.A(_115_),
    .B(_110_),
    .C(_179_),
    .Y(_194_));
 sky130_fd_sc_hd__nand3_1 _454_ (.A(_192_),
    .B(_193_),
    .C(_194_),
    .Y(_195_));
 sky130_fd_sc_hd__or4_1 _455_ (.A(net12),
    .B(net44),
    .C(net1),
    .D(net33),
    .X(_196_));
 sky130_fd_sc_hd__or4_1 _456_ (.A(net26),
    .B(net58),
    .C(net23),
    .D(net55),
    .X(_197_));
 sky130_fd_sc_hd__nor2_1 _457_ (.A(_196_),
    .B(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__and4_1 _458_ (.A(_191_),
    .B(_154_),
    .C(_195_),
    .D(_198_),
    .X(_199_));
 sky130_fd_sc_hd__and3_1 _459_ (.A(_178_),
    .B(_187_),
    .C(_199_),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_1 _460_ (.A(_200_),
    .X(_001_));
 sky130_fd_sc_hd__dfrtp_1 _461_ (.CLK(clknet_1_0__leaf_clk),
    .D(net74),
    .RESET_B(net65),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _462_ (.CLK(clknet_1_0__leaf_clk),
    .D(_002_),
    .RESET_B(net65),
    .Q(net68));
 sky130_fd_sc_hd__dfrtp_1 _463_ (.CLK(clknet_1_1__leaf_clk),
    .D(_003_),
    .RESET_B(net65),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _464_ (.CLK(clknet_1_1__leaf_clk),
    .D(net71),
    .RESET_B(net65),
    .Q(net66));
 sky130_fd_sc_hd__conb_1 _464__71 (.HI(net71));
 sky130_fd_sc_hd__dfrtp_1 _465_ (.CLK(clknet_1_1__leaf_clk),
    .D(net76),
    .RESET_B(net65),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _466_ (.CLK(clknet_1_0__leaf_clk),
    .D(_001_),
    .RESET_B(net65),
    .Q(eq_f));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__buf_1 hold1 (.A(net75),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net77),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_000_),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net66),
    .X(net75));
 sky130_fd_sc_hd__buf_1 hold5 (.A(net72),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(eq_f),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input1 (.A(in1[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(in1[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(in1[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(in1[1]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(in1[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(in1[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(in1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in1[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(in1[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in1[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in1[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(in1[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in1[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in1[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(in1[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in1[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(in1[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(in1[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(in1[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(in1[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(in1[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(in1[11]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(in1[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(in1[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(in1[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(in2[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(in2[10]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(in2[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(in2[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(in2[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(in2[14]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(in2[15]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(in1[12]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(in2[16]),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(in2[17]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(in2[18]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(in2[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(in2[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(in2[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(in2[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(in2[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(in2[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(in2[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(in1[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(in2[25]),
    .X(net50));
 sky130_fd_sc_hd__dlymetal6s2s_1 input51 (.A(in2[26]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(in2[27]),
    .X(net52));
 sky130_fd_sc_hd__dlymetal6s2s_1 input53 (.A(in2[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(in2[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(in2[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(in2[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(in2[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(in2[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(in2[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input6 (.A(in1[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input60 (.A(in2[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(in2[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(in2[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(in2[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(in2[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(rst),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in1[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(in1[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(in1[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(done));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(eq));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(great));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(inv));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(less));
endmodule

