// This is the unpowered netlist.
module fp_div (act,
    clk,
    div_zero,
    done,
    inexact,
    inv,
    ov,
    rst,
    un,
    in1,
    in2,
    out,
    round_m);
 input act;
 input clk;
 output div_zero;
 output done;
 output inexact;
 output inv;
 output ov;
 input rst;
 output un;
 input [31:0] in1;
 input [31:0] in2;
 output [31:0] out;
 input [2:0] round_m;

 wire \M00r[0] ;
 wire \M00r[10] ;
 wire \M00r[11] ;
 wire \M00r[12] ;
 wire \M00r[13] ;
 wire \M00r[14] ;
 wire \M00r[15] ;
 wire \M00r[16] ;
 wire \M00r[17] ;
 wire \M00r[18] ;
 wire \M00r[19] ;
 wire \M00r[1] ;
 wire \M00r[20] ;
 wire \M00r[21] ;
 wire \M00r[22] ;
 wire \M00r[23] ;
 wire \M00r[24] ;
 wire \M00r[2] ;
 wire \M00r[3] ;
 wire \M00r[4] ;
 wire \M00r[5] ;
 wire \M00r[6] ;
 wire \M00r[7] ;
 wire \M00r[8] ;
 wire \M00r[9] ;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire \div1i.quot[0] ;
 wire \div1i.quot[10] ;
 wire \div1i.quot[11] ;
 wire \div1i.quot[12] ;
 wire \div1i.quot[13] ;
 wire \div1i.quot[14] ;
 wire \div1i.quot[15] ;
 wire \div1i.quot[16] ;
 wire \div1i.quot[17] ;
 wire \div1i.quot[18] ;
 wire \div1i.quot[19] ;
 wire \div1i.quot[1] ;
 wire \div1i.quot[20] ;
 wire \div1i.quot[21] ;
 wire \div1i.quot[22] ;
 wire \div1i.quot[23] ;
 wire \div1i.quot[2] ;
 wire \div1i.quot[3] ;
 wire \div1i.quot[4] ;
 wire \div1i.quot[5] ;
 wire \div1i.quot[6] ;
 wire \div1i.quot[7] ;
 wire \div1i.quot[8] ;
 wire \div1i.quot[9] ;
 wire div_zero_f;
 wire div_zero_f_c;
 wire done0_reg;
 wire forward;
 wire forward_c;
 wire inv_f;
 wire inv_f_c;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \out_f[22] ;
 wire \out_f[23] ;
 wire \out_f[31] ;
 wire \out_f_c[22] ;
 wire \out_f_c[23] ;
 wire \out_f_c[31] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA__14293__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__14294__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__14295__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14295__B (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14295__C (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14296__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__A (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14297__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__14299__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__14300__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__14301__B (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14303__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__14304__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__14305__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__14306__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__A (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__B (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__C (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14307__D (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__14308__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__14310__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__14311__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__14312__B (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14313__A (.DIODE(_05386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14314__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__14315__B (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14316__A (.DIODE(_05386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14316__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__14321__A (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__A (.DIODE(_05496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14323__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__14327__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__14328__A (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14330__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14332__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__14336__B (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14340__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__14341__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__14342__A (.DIODE(_05705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14344__A (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14345__B (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14347__A (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14351__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__14352__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14354__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__14355__A (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14357__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__14367__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__14368__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__14369__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__14370__A (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14370__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__14372__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__14373__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__14373__B (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14374__A_N (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__14374__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__14377__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__14378__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__14379__A (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14379__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__14381__A_N (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14381__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__14382__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__A (.DIODE(_06155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14383__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14388__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__14390__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__14391__A (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14393__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__14396__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__14397__A (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14399__A (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14401__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__14418__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__14419__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__14419__B (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14420__A (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14420__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__14422__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__14423__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__14423__B (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14424__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__14425__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__14428__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14428__B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__14430__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__14431__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__14432__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__14433__A (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14433__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__14435__A (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__A (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14436__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__14437__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__14438__B (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14440__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__14441__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__14442__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__14443__A (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14443__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__14444__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__14445__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__14446__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14446__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__14456__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__14457__A2 (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14461__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__A (.DIODE(_07011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14465__B (.DIODE(_07055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14467__A (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14469__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__14474__A (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14475__A (.DIODE(_07011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14476__A (.DIODE(_07055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14478__A (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14482__C (.DIODE(_07242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14483__A (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14484__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__14488__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14488__B (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14488__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__14492__A (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14494__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__14495__A (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14500__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14501__A (.DIODE(_07011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14501__C (.DIODE(_07055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14504__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14507__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14507__B (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14509__B (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14510__A (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14511__C (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__14519__C (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__14521__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__14522__B (.DIODE(_05705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14524__B (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14525__A (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14526__C (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__14530__C (.DIODE(_07055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14532__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14541__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14543__A (.DIODE(_07011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14543__C (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__14545__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__14546__C (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__A (.DIODE(_07011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14551__C (.DIODE(_07055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14553__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__14556__A (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14557__B (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14558__C (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14569__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14570__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__14570__C (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__14573__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__14574__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__14576__B (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14577__A (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14578__C (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14580__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__14581__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__14583__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__14586__B (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14588__C (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14591__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14591__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__14592__C (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__14594__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__14597__B (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14598__A (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14599__C (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14601__A (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14604__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14604__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__14605__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__14612__A (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14614__B (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14616__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14617__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__14619__B1 (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14620__C (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14622__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14623__A (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14625__A (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14627__B1 (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14628__C (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14631__A (.DIODE(_07297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__B (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14634__C (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14635__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__14637__B (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14638__A (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14639__B (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14641__A (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14644__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__14647__B (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14649__C (.DIODE(_09076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14654__A (.DIODE(_08197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14672__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__B (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14673__C (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14675__B (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14676__A (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14677__B (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14680__A (.DIODE(_08197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14692__A (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14694__B (.DIODE(_09559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14696__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__14696__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__14696__S (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14697__B (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14698__S (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14699__B (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14704__A (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14705__B (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14709__B (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14712__S (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14713__B (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__14714__S (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__A1 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14726__B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__B (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__C (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__14727__D (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__A (.DIODE(_09943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14728__B (.DIODE(_05386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14732__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14734__B (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14742__A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__14742__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__14742__S (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14743__B (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14744__S (.DIODE(_07077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14751__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14752__B (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14755__A (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14756__B (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14763__A0 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__14763__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__14763__S (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14764__A (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14765__B (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14771__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__A (.DIODE(_10426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14772__B (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14774__A (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14777__B (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14781__B (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14784__A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__14784__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__14784__S (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14792__A (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14793__B (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14796__A (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14797__B (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14798__B (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14805__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__14805__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__14805__S (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14806__A (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14807__B (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14814__B (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14816__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14821__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14826__B1 (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14832__B (.DIODE(_08197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14833__A (.DIODE(_08197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14835__B (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14836__A (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14837__B (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14851__B (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14858__B (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14859__B (.DIODE(_09076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14861__A (.DIODE(_08197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14868__B (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14869__C (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14877__B (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14886__B (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14887__B (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14895__B (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14897__B (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14899__A1 (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14899__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__14899__B1 (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14902__B (.DIODE(_07242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14906__A (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14908__B (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14918__B (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14920__B (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14928__B (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14929__B (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14938__A (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14951__B (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14956__B (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14957__B (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14960__B (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14973__B (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14974__B (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14989__B (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14990__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14994__B (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14999__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__14999__A2 (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__14999__B1 (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15002__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15004__A (.DIODE(_12974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15007__A (.DIODE(_12974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15013__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15013__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15014__C (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15015__A (.DIODE(_12974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15017__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__15018__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15019__A (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15020__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15020__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15021__C (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15024__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__15024__B (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15026__B (.DIODE(_07242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15029__A (.DIODE(_13104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15030__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15032__B (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15033__C (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15037__B (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15038__A (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15043__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__15044__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15044__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15045__C (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15047__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__15048__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15048__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15049__C (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15055__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__15056__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15056__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15058__B (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15060__C (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15065__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__15066__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15066__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15068__B (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15069__C (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15074__A (.DIODE(_13104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15075__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15077__B (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15078__C (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15083__A (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15084__B (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15086__A (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15087__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15087__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15088__C (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15089__C (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15092__A (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15101__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__15102__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15102__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15104__B (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15105__C (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15112__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15114__B (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15115__C (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15127__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15128__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15135__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__15136__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15136__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15138__B (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15139__C (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15145__A (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15146__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15146__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15149__C (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15154__A (.DIODE(_12974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15155__A (.DIODE(_13072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15155__C (.DIODE(_12952_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15157__B (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15158__B (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15163__A (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15164__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15164__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15166__B (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15167__C (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15171__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__15172__A (.DIODE(_13137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15172__C (.DIODE(_13148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15174__B (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15175__C (.DIODE(_09076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15204__B (.DIODE(_13104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15205__A2 (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15206__A (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15208__B (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15210__A (.DIODE(_12974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15217__A (.DIODE(_13104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15219__A (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15220__B (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15231__B (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15233__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15234__C (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15238__B (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15241__B (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15255__B (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15258__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15259__B (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15266__B (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15269__B (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15270__B (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15276__B (.DIODE(_13104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15281__B (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15287__B (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15290__B (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15291__B (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15311__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15312__A (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15313__A (.DIODE(_02112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15314__A (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15316__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15321__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__15323__B (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15324__C (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15338__B (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15340__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15341__B (.DIODE(_09559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15345__A (.DIODE(_02112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15346__B (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15347__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15349__B (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15359__B (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15360__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15362__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15363__B (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15375__B (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15376__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15378__B (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15386__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__15387__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15389__B (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15393__B (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15400__B (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15401__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15403__B (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15404__B (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15414__B (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15415__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15417__B (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15418__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15423__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15424__B (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15428__B1 (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15435__B (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__15436__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15446__B (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15447__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15449__B (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15450__B (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15460__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15463__A (.DIODE(_02112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15465__B (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15466__B (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15479__B (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15480__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15482__B (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15483__B (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15488__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15496__B (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15497__B (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15499__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15505__A (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15506__B (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15509__B (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15511__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15514__B (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15516__B (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15517__C (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15520__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15523__B (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15525__B (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15526__C (.DIODE(_09076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15533__B1 (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15534__A (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15546__A (.DIODE(_02112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15547__B (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15549__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15554__A (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15555__C (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15558__B (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15561__C (.DIODE(_02090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15565__B (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15566__B (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15567__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15568__A (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15569__B (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15572__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15575__A (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15577__B (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15578__B (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15584__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15587__A (.DIODE(_02112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15588__B (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15589__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15591__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__15592__B (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15596__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15599__A (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15601__B (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15602__B (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__A (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15604__B (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15606__B (.DIODE(_07242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15610__B (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15611__B (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15615__A (.DIODE(_02142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15616__A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__15617__B (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15620__B (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15621__A (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15622__A2 (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15623__B (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15626__B (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15627__B (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15643__B (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15654__S (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15655__C (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15657__A (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15669__B (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15671__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15672__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15674__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15675__B (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15684__B (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15685__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15687__B (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15688__B (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15695__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15696__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15698__A (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15701__B (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__15702__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15704__B (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15708__B (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15723__B (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15724__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15725__B (.DIODE(_09559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15729__B1 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15730__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15732__B (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15733__B (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15739__B1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15740__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15742__B (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15743__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__15746__B1 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15747__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15749__A (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15750__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15754__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15763__B (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15767__A (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15768__B (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15770__A (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15777__B1 (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15778__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15780__B (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15781__B (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15784__B (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15792__B (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15793__B1 (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15794__C (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15795__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15798__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15799__B1 (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15802__B (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15810__B (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15811__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15813__A (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15814__B (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15818__B (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15819__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15820__B1 (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15821__B (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15826__B (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15827__A (.DIODE(_05023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15829__B (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15830__B (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15834__B (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15835__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15838__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__15855__A (.DIODE(_05212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15855__C (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15860__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__15861__C (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15862__A (.DIODE(_05212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15865__A (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15869__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15870__C (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15873__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15874__C (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15880__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__15881__C (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15884__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__15885__C (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15890__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15892__B (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15893__C (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15902__A (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15903__C (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15906__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15907__C (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15910__A (.DIODE(_05120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15910__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15910__C (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15917__A (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15918__C (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15920__A (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__15921__C (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15925__C (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15926__C (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15931__A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__15932__C (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15936__B (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15937__C (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15941__B (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15942__C (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15950__B1 (.DIODE(_09559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15957__A (.DIODE(_05115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15960__S (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15961__B (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15962__A_N (.DIODE(_05328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15962__B (.DIODE(_05115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15965__A (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15975__S (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15976__A (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15987__B (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__15989__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__15991__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__16001__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16004__A (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16005__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__16008__B (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16014__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__16025__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16026__B (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16031__B (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16034__B (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16035__A (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16035__B (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16038__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16039__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16042__A1 (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16049__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__16050__B (.DIODE(_05705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16054__B (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16056__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16066__B (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16067__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__16073__B (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16074__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__16083__B (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16084__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__16087__B (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16088__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__16105__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__16106__B (.DIODE(_06155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16110__A (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16113__B (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16114__A (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16118__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__16121__A (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16123__A (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16128__B (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16131__B (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16133__B (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16141__B (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16151__B (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16157__B (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16160__C (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16161__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16161__C (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16165__A (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16168__A (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16171__B (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16172__C (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16176__A (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16180__B (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16181__C (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16186__A (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16190__B (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16191__C (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16194__A (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16198__B (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16199__C (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16220__B (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16221__B (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16222__A (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16223__A2 (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16224__A (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16225__B (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16230__B (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16231__B_N (.DIODE(_05333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16233__B (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16234__C (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16237__A (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16258__B (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__16259__B (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16267__B (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16268__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__16278__B (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16279__B (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16281__B (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16282__B (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16283__S (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16284__A (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16285__B (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16298__B (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16299__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__16313__B (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16314__B (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16319__B (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16320__A (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16322__B (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16323__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16324__S (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16326__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__16327__B (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16340__S (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16341__A (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16342__B (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16350__S (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16351__A (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16352__B (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16356__B (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16358__C (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__16370__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__16371__B (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16372__B (.DIODE(_10426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16373__B (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16388__B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__16389__B (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16394__B (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16395__B (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16397__B (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16398__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16399__S (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16400__A (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16401__B (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16415__B (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16420__A (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16420__B (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16428__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__16429__B (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16435__B (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16439__B (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16440__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__16441__A1 (.DIODE(_05496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16441__A2 (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16441__B1 (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16446__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__16451__B (.DIODE(_05705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16452__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__16459__B (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16462__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16471__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__16472__B (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16478__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__16480__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16484__B (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__B (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16489__C (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16492__B (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16493__B (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16500__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16503__A (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16504__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16513__B (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16514__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__16521__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__16523__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16534__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16535__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16536__B1 (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16538__B (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16544__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16547__A (.DIODE(_09076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16555__B (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16555__C (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16557__A (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16558__B (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16559__A (.DIODE(_05496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16559__B (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16560__A (.DIODE(_07242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16564__A (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16564__B (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16566__B (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16569__B (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16570__C (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16573__A (.DIODE(_11777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16580__A (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16580__B (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16582__B (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16583__B (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__A (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16589__B (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16591__B (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16592__B (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__A (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16601__B (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16603__A (.DIODE(_12029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16604__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16605__B (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16611__A (.DIODE(_05831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16611__B (.DIODE(_05832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16613__B (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16614__A (.DIODE(_07703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16615__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16631__A (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16632__A (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16641__B (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16642__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__16650__B (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16651__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__16664__B (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__16665__B (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16671__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16674__B (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16675__B (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16686__B (.DIODE(_06155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16687__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__16696__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16697__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16700__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__16704__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16707__A (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16708__A (.DIODE(_08384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16709__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16715__A (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16717__A (.DIODE(_08274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16718__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16719__B (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16731__B (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16732__B (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16741__B (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16743__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__16757__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__16761__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__16762__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16763__B (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16766__B (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16775__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16777__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16778__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16781__B (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16782__B (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16788__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16789__A (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16791__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__16792__B (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16796__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16797__A (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16799__A (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16800__B (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16805__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16806__A (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16808__A (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16809__B (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16821__B (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16823__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__16837__B (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16838__B (.DIODE(_10426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16846__B (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16847__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__16859__B (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__16860__B (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16865__C (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16866__B (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16868__B (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16869__B (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16877__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16878__A (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16880__B (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16881__B (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16886__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16887__A (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16890__B (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16891__B (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16901__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16902__B (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16904__B (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16905__A (.DIODE(_10690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16906__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16919__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__A (.DIODE(_06383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16924__B (.DIODE(_06385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16926__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16935__B (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16937__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__16939__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__16949__B (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16953__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__16956__B (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__16960__B (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16970__B (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16971__A1 (.DIODE(_05496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16971__A2 (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__16971__B1 (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16972__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__16978__B (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16981__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__16988__B (.DIODE(_05705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16989__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__16996__A (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16997__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__16999__A (.DIODE(_05738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17010__B (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17013__B (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17014__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__17017__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17026__B (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17040__B (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17041__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__17047__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__17048__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17049__B (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17066__B (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__17067__B (.DIODE(_06155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17074__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17075__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17077__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__17078__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17080__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17087__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17088__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17090__A (.DIODE(_08527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17091__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17092__A (.DIODE(_08505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17093__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17104__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17105__A (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17106__B (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17108__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17109__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17110__B (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17112__A (.DIODE(_08406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17113__B1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17119__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17124__B (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17125__A (.DIODE(_07242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17126__A (.DIODE(_05496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17126__B (.DIODE(_06223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17127__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17130__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17133__A (.DIODE(_07539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17134__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17137__A (.DIODE(_07560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17138__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17139__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17139__B (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17139__C (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17142__A (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17150__A (.DIODE(_06383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17152__A (.DIODE(_13588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17153__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17154__A (.DIODE(_11579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17155__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17158__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17163__A (.DIODE(_08066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17164__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17165__A (.DIODE(_08055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17166__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17177__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17178__B (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17186__B (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17187__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17205__A (.DIODE(_11140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17206__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17207__A (.DIODE(_08746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17208__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17214__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17215__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17217__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17218__B (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17226__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17227__A (.DIODE(_06388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17229__A (.DIODE(_09054_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17230__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17231__A (.DIODE(_09076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17232__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17234__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17236__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17238__A (.DIODE(_08966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17239__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17240__A (.DIODE(_08944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17241__C (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17253__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17259__A (.DIODE(_09361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17265__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17266__B (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17274__B (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17275__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__17276__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17286__A (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17288__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17289__A (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17291__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17295__B (.DIODE(_06548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17296__A (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17298__A (.DIODE(_09548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17299__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17300__A (.DIODE(_09559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17301__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17305__A (.DIODE(_09383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17306__B (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17309__A (.DIODE(_09987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17317__B (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17318__A (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17319__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17325__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__17326__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17327__B (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17337__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17338__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17340__A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17341__A (.DIODE(_09735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17344__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17345__A (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17347__A (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17348__B (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17353__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17359__A (.DIODE(_10426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17360__B (.DIODE(_10426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17366__B (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17368__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__17369__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17379__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17380__A (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17382__B (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17383__B (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17389__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17390__A (.DIODE(_10240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17391__B (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17392__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17394__A (.DIODE(_10251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17395__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17402__A (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17403__B (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17409__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17410__B (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17412__B (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17413__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17424__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__17425__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17426__B (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17431__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17432__B (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17434__A (.DIODE(_10887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17435__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17436__A (.DIODE(_10909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17437__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17451__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17456__A (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17456__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17458__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17464__A (.DIODE(_05496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17465__A (.DIODE(_05474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17466__A1 (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17466__A2 (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17467__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17468__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17469__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__17470__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17473__C (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17475__B (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17476__A (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17476__B (.DIODE(_06784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17477__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17481__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17483__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17486__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17487__A (.DIODE(_07308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17488__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17491__A (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17503__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__17504__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17505__A (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17506__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17512__A (.DIODE(_05705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17513__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17514__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__17515__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17523__A (.DIODE(_05178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17524__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17527__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__17528__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17534__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17537__B (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17543__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17545__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17546__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17552__A (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17552__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17554__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17555__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17564__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17566__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17567__A (.DIODE(_12051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17568__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17574__B (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17576__A (.DIODE(_07725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17577__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17578__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17600__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__17601__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17602__A (.DIODE(_05299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17603__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17609__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17616__A (.DIODE(_05310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17617__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17619__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__17621__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17624__A (.DIODE(_05321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17625__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17626__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__17627__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17633__B (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17641__B (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17642__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17644__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17645__B (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17653__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17655__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17656__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17660__A (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17661__A1 (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17661__A2 (.DIODE(_06970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17663__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17664__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17669__A (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17672__A (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17673__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17689__A (.DIODE(_05288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17690__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17691__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__17692__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17708__A (.DIODE(_06045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17709__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17710__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__17711__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17717__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17718__B (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17734__A (.DIODE(_06155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17735__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17736__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__17737__C (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17742__B (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17743__B (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17745__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17746__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17753__B (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17754__A (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17756__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17757__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17761__B (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17762__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17764__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17765__B (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17769__B (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17770__A (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17772__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17773__A (.DIODE(_08296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17774__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17789__B (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17790__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17806__B (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17807__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17812__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17813__B (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17827__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17828__B (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17832__A (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17834__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17835__A (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17837__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17838__B (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17843__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17844__A (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17846__B (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17847__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__17848__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17852__B (.DIODE(_07171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17853__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__17855__A (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17856__B (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17860__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17861__A (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17863__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17864__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17877__B (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17878__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17893__A (.DIODE(_10426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17894__B (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17895__B (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17903__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__17904__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17905__B (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17911__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17912__B (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17914__A (.DIODE(_10701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17915__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17916__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17930__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17931__B (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17936__C (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17937__B (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17939__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17940__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17945__C (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17946__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17948__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17949__B (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17954__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17955__A (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__17956__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17958__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17970__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17975__A (.DIODE(_07540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17975__B (.DIODE(_07538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17977__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17988__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17990__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__17992__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18002__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18006__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18009__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18013__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18023__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18024__A1 (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18024__A2 (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18025__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18031__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18034__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18041__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18042__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18049__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18051__A (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18062__B (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18065__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18066__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18069__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18078__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18092__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18093__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18099__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18100__A (.DIODE(_06012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18101__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18118__B (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18119__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18126__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18128__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18129__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18137__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18139__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18140__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18152__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18153__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18156__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18157__B (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18159__B1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18165__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18168__B (.DIODE(_07538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18168__C (.DIODE(_07540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18170__B (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__A (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18171__B (.DIODE(_07383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18172__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18176__A (.DIODE(_07538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18176__B (.DIODE(_07540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18178__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18181__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18182__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18182__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18185__A (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18193__A (.DIODE(_07538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18193__B (.DIODE(_07540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18195__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18196__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18199__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__A (.DIODE(_07538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18202__B (.DIODE(_07540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18204__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18205__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18214__A (.DIODE(_07538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18214__B (.DIODE(_07540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18216__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18217__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18223__B (.DIODE(_07540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18225__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18226__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18244__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18245__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18252__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18254__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18255__B (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18264__A (.DIODE(_07542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18266__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18267__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18273__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18274__C (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18286__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18298__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18299__B (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18307__A (.DIODE(_05375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18308__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18309__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18321__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18322__A (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18324__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18328__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18329__A (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18331__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18332__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18336__B (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18345__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18346__A (.DIODE(_06737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18347__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18353__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18354__A (.DIODE(_06814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18355__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18365__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18366__A (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18368__A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18371__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18372__A (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18374__A (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18375__B (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18379__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18385__A (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18386__B (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18394__A (.DIODE(_06704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18395__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18396__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18409__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18410__A (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18412__A (.DIODE(_10481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18413__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18414__B (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18420__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18421__B (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18423__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18424__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18430__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18431__A (.DIODE(_06550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18432__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18438__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18439__B (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18441__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18442__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18456__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18457__B (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18462__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18463__B (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18465__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18466__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18479__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__A (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18484__B (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18486__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__A1 (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18492__A2 (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18493__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18494__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18497__B (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18497__C (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18499__B (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__A (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18500__B (.DIODE(_07918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18501__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18505__A (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18505__B (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18507__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18510__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18511__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18514__A (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18526__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18527__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18533__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18534__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18542__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18545__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18551__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18554__A (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18555__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18561__A (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18561__B (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18563__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18564__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18570__A (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18570__B (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18572__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18573__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18582__A (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18582__B (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18584__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18585__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18591__A (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18591__B (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18593__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18594__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18616__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18617__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18623__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18630__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18633__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18636__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18637__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18643__B (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18651__B (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18652__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__18654__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18655__B (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18663__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__18665__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18666__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18670__A (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18671__A1 (.DIODE(_08096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18671__A2 (.DIODE(_08098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18673__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18674__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18679__A (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18682__A (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18683__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18699__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18700__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18716__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18717__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18723__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18724__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18740__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18741__C (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18746__B (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18747__B (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18749__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18750__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18757__B (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18758__A (.DIODE(\div1i.quot[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18760__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18761__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18765__B (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18766__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__18768__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18769__B (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18773__A (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18774__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18775__A (.DIODE(\div1i.quot[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18777__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18778__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18793__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18794__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18810__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18811__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18816__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18817__A (.DIODE(_05408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18818__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18832__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18833__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18838__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18839__A (.DIODE(\div1i.quot[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18841__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18842__B (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18847__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18848__A (.DIODE(\div1i.quot[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18850__B (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18851__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18855__B (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18856__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__18858__A (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18859__B (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18863__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18864__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__18866__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18867__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18881__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18882__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18897__B (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18898__A (.DIODE(_06649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18899__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18904__C (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18905__B (.DIODE(_08280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18907__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18908__B (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18914__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18915__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__18917__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18918__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18924__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18925__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18931__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18932__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__18934__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18935__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18949__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18950__A (.DIODE(_06594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18951__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18956__C (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18957__B (.DIODE(\div1i.quot[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__18959__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18960__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18974__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18979__A (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18979__B (.DIODE(_08640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18992__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18994__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__18996__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19006__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19010__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19013__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19017__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19027__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19028__A1 (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19028__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__19029__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19035__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19038__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19045__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19046__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19053__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19055__A (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19066__A (.DIODE(_05255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19067__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19070__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19071__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19074__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19083__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19097__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19098__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19104__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19105__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19122__B (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19123__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19132__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19133__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19143__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19144__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19157__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19161__B (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19163__B1 (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19172__B (.DIODE(_08640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19172__C (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19174__A (.DIODE(_05983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19176__A (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19176__B (.DIODE(_08416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19177__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19181__A (.DIODE(_08640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19181__B (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19183__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19186__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19187__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__A (.DIODE(_08640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19198__B (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19200__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19201__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19207__A (.DIODE(_08640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19207__B (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19209__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19210__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19219__A (.DIODE(_08640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19219__B (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19221__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19222__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__A (.DIODE(_08640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19228__B (.DIODE(_08642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19230__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19231__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19249__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19250__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19259__B (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19260__A (.DIODE(_08834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19261__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19272__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19273__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19279__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19280__C (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19292__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19304__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19305__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19313__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19314__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19326__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19327__A (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19329__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19333__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19334__A (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19336__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19337__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19341__B (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19350__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19351__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19357__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19358__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19368__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19369__A (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19371__A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19374__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19375__A (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19377__A (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19378__B (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19382__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19389__A (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19390__B (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19398__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19399__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19412__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19413__A (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19415__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19416__B (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19422__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19423__B (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19425__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19426__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19433__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19434__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19440__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19441__B (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19443__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19444__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19457__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19458__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19463__C (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19464__B (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19466__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19467__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19480__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19485__A (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19485__B (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19487__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__A1 (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19493__A2 (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19494__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19495__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19498__B (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19498__C (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19501__A (.DIODE(_06979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19502__B (.DIODE(_09022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19503__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__A (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19507__B (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19509__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19512__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__B (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19514__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19529__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19530__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19536__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19537__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19545__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19548__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19554__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19557__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19563__A (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19563__B (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19565__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19566__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19572__A (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19572__B (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19574__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19575__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19584__A (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19584__B (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19586__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19587__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19593__A (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19593__B (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19595__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19596__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19618__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19619__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19625__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19632__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19635__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19638__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19639__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19645__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19653__B (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19656__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19657__B (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19664__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__19665__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__19667__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19668__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19672__A (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19673__A1 (.DIODE(_09195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19673__A2 (.DIODE(_09198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19675__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19676__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19678__A (.DIODE(_05915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19682__A (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19685__A (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19686__B (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19702__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19703__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19719__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19720__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19726__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19727__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19743__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19744__C (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19749__B (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19750__B (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19752__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19753__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19760__B (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19761__A (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19763__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19764__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19768__B (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19769__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__19771__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19772__B (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19776__A (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19777__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19778__A (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19780__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19781__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19796__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19797__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19813__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19814__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19819__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19820__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19834__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19835__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19840__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19841__A (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19843__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19844__B (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19849__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19850__A (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19852__B (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19853__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19857__B (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19858__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__19860__A (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19861__B (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19865__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19866__A (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19868__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19869__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19883__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19884__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19899__B (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19900__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19905__C (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19906__B (.DIODE(_09380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19908__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19909__A (.DIODE(_06348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19910__B (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19916__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19917__A (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19919__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19920__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19926__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19927__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19933__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19934__B (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19936__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19937__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19951__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19952__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19957__C (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19958__B (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__19960__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19961__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19975__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19980__A (.DIODE(_09740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19980__B (.DIODE(_09741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19993__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19995__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__19997__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20007__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20011__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20014__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20018__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20028__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20029__A2 (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20029__B1 (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20030__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20036__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20039__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20046__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20047__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20054__A (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20055__B (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20057__A (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20068__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20071__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20072__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20075__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20084__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20098__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20099__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20105__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20106__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20123__B (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20124__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20133__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20134__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20144__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20145__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20158__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20162__B (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20164__A (.DIODE(_06592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20165__B1 (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20174__B (.DIODE(_09740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20174__C (.DIODE(_09741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20177__B (.DIODE(_09518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20178__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20182__A (.DIODE(_09740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20182__B (.DIODE(_09741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20184__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20187__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20188__B (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20188__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20199__A (.DIODE(_09740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20199__B (.DIODE(_09741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20201__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20202__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20208__A (.DIODE(_09740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20208__B (.DIODE(_09741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20210__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20211__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20220__A (.DIODE(_09740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20220__B (.DIODE(_09741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20222__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20223__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20229__A (.DIODE(_09740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20229__B (.DIODE(_09741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20231__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20232__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20250__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20251__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20260__B (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20261__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20272__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20273__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20279__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20280__C (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20292__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20304__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20305__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20313__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20314__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20326__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20327__A (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20329__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20333__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20334__A (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20336__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20337__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20341__A (.DIODE(_06805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20342__B (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20351__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20352__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20358__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20359__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20369__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20370__A (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20372__A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20373__A (.DIODE(_06844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20376__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20377__A (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20379__A (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20380__B (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20384__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20391__A (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20392__B (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20400__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20401__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20414__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20415__A (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20417__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20418__B (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20424__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20425__B (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20427__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20428__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20435__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20436__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20442__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20443__B (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20445__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20446__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20459__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20460__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20465__C (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20466__B (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20468__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20469__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20482__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20487__A (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20487__B (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20489__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__20495__A2 (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20495__B1 (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20496__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20497__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20500__B (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20500__C (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20503__B (.DIODE(_10120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20504__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20508__A (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20508__B (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20510__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20513__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20514__B (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20514__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20529__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20530__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20536__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20537__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20545__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20548__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20554__B (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20557__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20563__A (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20563__B (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20565__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20566__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20572__A (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20572__B (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20574__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20575__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20584__A (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20584__B (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20586__B (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20587__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20593__A (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20593__B (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20595__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20596__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20618__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20619__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20625__B (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20632__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20635__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20638__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20639__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20645__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20653__B (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20654__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__20656__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20657__B (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20665__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__20667__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20668__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20672__A (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__A1 (.DIODE(_10296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20673__A2 (.DIODE(_10298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20675__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20676__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20681__A (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20684__A (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20685__B (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20701__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20702__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20718__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20719__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20725__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20726__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20742__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20743__C (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20748__B (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20749__B (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20751__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20752__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20759__B (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20760__A (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20762__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20763__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20767__B (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20768__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__20770__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20771__B (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20775__B (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20776__A (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20778__B (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20779__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20794__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20795__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20811__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20812__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20817__B (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20818__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20832__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20833__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20837__A (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20839__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20840__A (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20842__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20843__B (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20848__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20849__A (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20851__B (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20852__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20856__B (.DIODE(_10478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20857__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__20859__A (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20860__B (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20864__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20865__A (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20867__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20868__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20881__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20882__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20897__A (.DIODE(_07450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20898__B (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20899__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20907__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20908__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20914__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20915__B (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20917__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20918__B (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20932__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20933__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20938__C (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20939__B (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20941__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20942__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20947__C (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20948__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20950__A (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20951__B (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20956__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20957__A (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__20958__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20960__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20972__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20977__A (.DIODE(_10836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20977__B (.DIODE(_10835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20979__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20990__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20992__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__20994__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21004__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21008__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21011__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21015__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21025__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21026__A2 (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21026__B1 (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21027__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21033__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21036__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21043__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21044__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21051__B (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21053__A (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21064__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21067__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21068__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21071__A (.DIODE(_05896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21072__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21081__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21095__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21096__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21102__B (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21103__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21120__B (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21121__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21129__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21131__B (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21132__B (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21140__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21142__B (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21143__B (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21155__A (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21156__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21159__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21160__B (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21162__B1 (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21171__B (.DIODE(_10835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21171__C (.DIODE(_10836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21174__B (.DIODE(_10683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21175__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21179__A (.DIODE(_10835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21179__B (.DIODE(_10836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21181__B (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21184__B (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21185__B (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21185__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21190__A (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21194__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21199__A (.DIODE(_10835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21199__B (.DIODE(_10836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21201__B (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21202__B (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21205__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21208__A (.DIODE(_10835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21208__B (.DIODE(_10836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21210__B (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21211__B (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21216__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21220__A (.DIODE(_10835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21220__B (.DIODE(_10836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21222__A (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21223__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21224__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21230__A (.DIODE(_10835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21230__B (.DIODE(_10836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21232__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21233__A (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21234__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21250__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21252__B (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21253__B (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21260__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21262__B (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21263__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21272__A (.DIODE(_10838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21274__B (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21275__B (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21281__B (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21282__C (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21294__A (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21295__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21307__A (.DIODE(_06207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21308__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21309__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21317__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21318__B (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21330__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21331__A (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21333__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21338__A (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21340__B (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21341__B (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21345__B (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21353__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21354__B (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21360__B (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21361__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21371__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21372__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21374__A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21377__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21378__A (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21380__A (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21381__B (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21385__B (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21391__A (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21392__B (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21400__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21401__B (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21414__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21415__A (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21417__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21418__B (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21424__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21425__B (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21427__B (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21428__B (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21433__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21434__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21448__B (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21449__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21454__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21455__B (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21457__B (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21458__B (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21464__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21465__B (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21467__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21468__A (.DIODE(_06366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21469__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21481__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21486__A (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21486__B (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21488__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__21494__A2 (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21494__B1 (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21495__B (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21496__B (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21499__B (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21499__C (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21501__B (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21502__A (.DIODE(_06607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21503__B (.DIODE(_11222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21504__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21508__A (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21508__B (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21510__A (.DIODE(_06615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21511__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21514__A (.DIODE(_06620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21515__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21516__B (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21516__C (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21519__A (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21529__B (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21530__B (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21536__B (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21537__B (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21545__B (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21548__B (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21554__B (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21557__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21563__A (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21563__B (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21565__A (.DIODE(_06636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21566__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21567__A (.DIODE(_06639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21568__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21574__A (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21574__B (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21576__A (.DIODE(_06651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21577__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21578__A (.DIODE(_06648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21579__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21588__A (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21588__B (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21590__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21591__B (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21597__A (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21597__B (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21599__B (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21600__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21622__B (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21623__B (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21630__A (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21637__B (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21640__B (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21643__B (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21644__B (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21649__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21657__B (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21658__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__21660__A (.DIODE(_06731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21661__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21662__A (.DIODE(_06733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21663__B (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21671__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__21673__A (.DIODE(_06721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21674__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21675__A (.DIODE(_06723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21676__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21679__A1 (.DIODE(_11392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21679__A2 (.DIODE(_11395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21683__A (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21685__A (.DIODE(_06695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21686__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21687__A (.DIODE(_06697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21688__C (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21693__A (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21696__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21697__B (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21713__B (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21714__B (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21730__B (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21731__B (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21737__A (.DIODE(_06521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21738__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21739__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21755__B (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21756__C (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21761__B (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21762__B (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21764__A (.DIODE(_06554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21765__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21766__A (.DIODE(_06556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21767__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21774__B (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21775__A (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21777__A (.DIODE(_06568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21778__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21779__A (.DIODE(_06570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21780__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21784__B (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21785__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__21787__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21788__B (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21792__A (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21793__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21794__A (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21796__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21797__B (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21812__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21813__A (.DIODE(_06772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21814__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21830__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21831__A (.DIODE(_06827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21832__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21837__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21838__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21852__A (.DIODE(_06819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21853__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21854__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21859__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21860__A (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21862__A (.DIODE(_06856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21863__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21864__A (.DIODE(_06809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21865__B (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21870__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21871__A (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21873__B (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21874__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21878__B (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21879__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__21881__A (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21882__B (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21886__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21887__A (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21889__A (.DIODE(_06797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21890__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21891__A (.DIODE(_06799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21892__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21906__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21907__A (.DIODE(_06874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21908__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21923__B (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21924__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21929__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21930__B (.DIODE(_11581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21932__A (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21933__B (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21939__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21940__A (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21942__A (.DIODE(_06903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21943__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21944__A (.DIODE(_06898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21945__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21951__B (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21952__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21958__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21959__B (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21961__B (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21962__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21977__A (.DIODE(_06936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21978__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21979__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21984__C (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21985__B (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__21987__A (.DIODE(_06947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21988__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21989__A (.DIODE(_06949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__21990__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22004__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22009__A (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22009__B (.DIODE(_11969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22022__A (.DIODE(_07226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22023__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22024__A (.DIODE(_07128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22026__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22028__A (.DIODE(_07228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22029__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22039__A (.DIODE(_07146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22040__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22044__A (.DIODE(_07157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22045__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22048__A (.DIODE(_07149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22049__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22053__A (.DIODE(_07130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22054__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22064__A (.DIODE(_06982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22065__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22067__A (.DIODE(_09228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22068__A1 (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22068__A2 (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22068__B1 (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22069__A (.DIODE(_06984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22070__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22076__A (.DIODE(_07043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22077__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22080__A (.DIODE(_07048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22081__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22088__A (.DIODE(_07031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22089__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22090__A (.DIODE(_07034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22091__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22098__B (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22100__A (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22111__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22114__A (.DIODE(_07024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22115__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22116__A (.DIODE(_07021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22117__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22120__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22129__A (.DIODE(_07155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22130__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22144__A (.DIODE(_07247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22145__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22146__A (.DIODE(_07249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22147__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22153__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22154__B (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22171__A (.DIODE(_07278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22172__B (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22173__A (.DIODE(_07276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22174__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22183__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22184__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22194__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22195__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22207__A (.DIODE(_07318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22209__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22213__B (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22215__B1 (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22224__B (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22224__C (.DIODE(_11969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22226__B (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22227__A (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22227__B (.DIODE(_11731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22228__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22232__A (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22232__B (.DIODE(_11969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22234__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22237__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22238__A (.DIODE(_07004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22239__B (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22239__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22242__A (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22250__A (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22250__B (.DIODE(_11969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22252__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22253__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22259__A (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22259__B (.DIODE(_11969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22261__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22262__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22271__A (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22271__B (.DIODE(_11969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22273__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22274__A (.DIODE(_07092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22275__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22281__A (.DIODE(_11968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22281__B (.DIODE(_11969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22283__A (.DIODE(_07102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22284__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22285__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22303__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22304__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22313__B (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22314__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22325__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22326__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22332__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22333__C (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22345__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22357__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22358__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22366__B (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22367__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22379__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22380__A (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22382__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22386__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22387__A (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22389__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22390__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22394__B (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22403__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22404__B (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22410__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22411__B (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22421__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22422__A (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22424__A (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22427__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22428__A (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22430__A (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22431__B (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22435__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22442__A (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22443__B (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22451__B (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22452__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22465__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22466__A (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22468__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22469__B (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22475__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22476__B (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22478__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22479__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22486__B (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22487__A (.DIODE(_07461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22488__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22494__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22495__B (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22497__A (.DIODE(_07474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22498__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22499__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22513__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22514__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22519__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22520__B (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22522__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22523__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22536__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22541__A (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22541__B (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22543__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__22549__A1 (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22549__A2 (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22549__B1 (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22550__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22551__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22554__B (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22554__C (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22556__B (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22557__A (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22557__B (.DIODE(_12374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22558__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22562__A (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22562__B (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22564__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22567__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22568__B (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22568__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22571__A (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22583__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22584__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22590__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22591__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22599__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22602__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22608__B (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22611__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22617__A (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22617__B (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22619__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22620__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22626__A (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22626__B (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22628__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22629__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22638__A (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22638__B (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22640__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22641__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22647__A (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22647__B (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22649__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22650__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22672__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22673__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22679__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22686__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22689__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22692__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22693__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22699__B (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22707__B (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22708__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__22710__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22711__B (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22719__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__22721__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22722__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22726__A (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22727__A1 (.DIODE(_12551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22727__A2 (.DIODE(_12553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22729__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22730__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22735__A (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22738__A (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22739__A (.DIODE(_09410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22740__B (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22756__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22757__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22773__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22774__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22780__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22781__A (.DIODE(_07677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22782__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22798__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22799__C (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22804__B (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22805__B (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22807__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22808__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22815__B (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22816__A (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22818__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22819__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22823__B (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22824__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__22826__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22827__B (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22831__A (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22832__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22833__A (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22835__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22836__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22851__A (.DIODE(_07905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22852__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22853__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22869__A (.DIODE(_07957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22870__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22871__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22876__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22877__B (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22891__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22892__A (.DIODE(_07948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22893__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22898__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22899__A (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22901__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22902__B (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22907__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22908__A (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22910__B (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22911__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22915__B (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22916__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__22918__A (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22919__B (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22923__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22924__A (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22926__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22927__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22941__A (.DIODE(_08001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22942__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22943__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22958__B (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22959__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22964__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22965__B (.DIODE(_12734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22967__A (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22968__A (.DIODE(_09664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22969__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22975__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22976__A (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22978__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22979__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22985__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22986__A (.DIODE(_08041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22987__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22993__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22994__B (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__22996__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__22997__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23011__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23012__B (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23017__C (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23018__B (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23020__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23021__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23035__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23040__A (.DIODE(_13100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23040__B (.DIODE(_13098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23053__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23055__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23057__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23067__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23071__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23074__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23078__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23088__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23089__A1 (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23089__A2 (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23089__B1 (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23090__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23096__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23099__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23106__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23107__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23114__A (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23115__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23117__A (.DIODE(_09823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23128__A (.DIODE(_08738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23129__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23132__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23133__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23136__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23145__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23159__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23160__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23166__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23167__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23184__B (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23185__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23194__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23195__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23205__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23206__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23219__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23223__B (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23225__A (.DIODE(_09944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23226__B1 (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23235__B (.DIODE(_13098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23235__C (.DIODE(_13100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23237__B (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23238__A (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23238__B (.DIODE(_12872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23239__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23243__A (.DIODE(_13098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23243__B (.DIODE(_13100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23245__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23248__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23249__B (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23249__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23253__A (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23262__A (.DIODE(_13098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23262__B (.DIODE(_13100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23264__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23265__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23271__A (.DIODE(_13098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23271__B (.DIODE(_13100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23273__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23274__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23283__A (.DIODE(_13098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23283__B (.DIODE(_13100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23285__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23286__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23292__A (.DIODE(_13098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23292__B (.DIODE(_13100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23294__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23295__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23313__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23314__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23323__B (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23324__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23335__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23336__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23342__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23343__C (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23355__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23367__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23368__A (.DIODE(_08465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23369__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23377__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23378__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23390__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23391__A (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23393__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23397__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23398__A (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23400__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23401__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23405__A (.DIODE(_10138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23406__B (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23415__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23416__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23422__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23423__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23433__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23434__A (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23436__A (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23437__A (.DIODE(_10173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23440__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23441__A (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23443__A (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23444__B (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23448__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23455__A (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23456__B (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23464__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23465__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23478__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23479__A (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23481__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23482__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23488__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23489__B (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23491__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23492__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23499__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23500__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23506__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23507__B (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23509__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23510__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23523__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23524__A (.DIODE(_08611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23525__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23530__C (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23531__B (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23533__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23534__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23547__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23552__A (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23552__B (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23554__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__23560__A1 (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23560__A2 (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23560__B1 (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23561__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23562__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23565__B (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23565__C (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23567__A (.DIODE(_11069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23568__B (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23569__A (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23569__B (.DIODE(_13483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23570__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23574__A (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23574__B (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23576__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23579__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23580__B (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23580__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23583__A (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23593__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23594__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23600__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23601__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23609__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23612__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23618__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23621__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23627__A (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23627__B (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23629__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23630__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23636__A (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23636__B (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23638__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23639__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23648__A (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23648__B (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23650__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23651__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23657__A (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23657__B (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23659__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23660__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23682__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23683__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23689__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23696__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23699__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23702__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23703__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23709__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23717__B (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23718__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__23720__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23721__B (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23729__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__23731__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23732__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23736__A (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23737__A1 (.DIODE(_13660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23737__A2 (.DIODE(_13662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23739__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23740__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23745__A (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23748__A (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23749__B (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23765__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23766__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23782__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23783__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23789__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23790__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23806__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23807__C (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23812__B (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23813__B (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23815__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23816__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23823__B (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23824__A (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23826__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23827__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23831__B (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23832__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__23834__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23835__B (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23839__B (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23840__A (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23842__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23843__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23858__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23859__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23875__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23876__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23881__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23882__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23896__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23897__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23901__A (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23903__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23904__A (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23906__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23907__B (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23912__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23913__A (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23915__B (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23916__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23920__B (.DIODE(_13842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23921__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__23923__A (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23924__B (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23928__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23929__A (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23931__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23932__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23946__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23947__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23962__A (.DIODE(_10749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23963__B (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23964__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23972__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23973__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23979__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23980__B (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__23982__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23983__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23997__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__23998__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24003__C (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24004__B (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24006__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24007__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24012__C (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24013__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24015__A (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24016__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24021__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24022__A (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24023__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24025__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24037__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24042__A (.DIODE(_14198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24042__B (.DIODE(_14200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24055__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24057__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24059__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24069__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24073__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24076__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24080__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24090__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24091__A1 (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24091__A2 (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24091__B1 (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24092__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24098__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24101__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24108__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24109__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24116__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24118__A (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24129__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24132__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24133__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24136__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24145__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24159__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24160__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24166__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24167__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24184__B (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24185__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24194__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24195__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24205__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24206__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24219__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24223__B (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24225__B1 (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24234__B (.DIODE(_14198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24234__C (.DIODE(_14200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24236__B (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24237__A (.DIODE(_12032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24238__B (.DIODE(_14046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24239__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24243__A (.DIODE(_14198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24243__B (.DIODE(_14200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24245__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24248__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24249__A (.DIODE(_12033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24250__B (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24250__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24253__A (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24261__A (.DIODE(_14198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24261__B (.DIODE(_14200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24263__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24264__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24270__A (.DIODE(_14198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24270__B (.DIODE(_14200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24272__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24273__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24282__A (.DIODE(_14198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24282__B (.DIODE(_14200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24284__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24285__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24291__A (.DIODE(_14198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24291__B (.DIODE(_14200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24293__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24294__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24312__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24313__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24322__B (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24323__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24334__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24335__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24341__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24342__C (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24354__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24366__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24367__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24375__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24376__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24388__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24389__A (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24391__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24395__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24396__A (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24398__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24399__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24403__B (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24412__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24413__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24419__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24420__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24430__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24431__A (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24433__A (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24436__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24437__A (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24439__A (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24440__B (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24444__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24450__A (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24451__B (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24459__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24460__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24473__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24474__A (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24476__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24477__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24483__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24484__B (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24486__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24487__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24493__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24494__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24500__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24501__B (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24503__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24504__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24518__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24519__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24524__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24525__B (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24527__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24528__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24541__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24546__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24546__B (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24548__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__24553__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__24554__A2 (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24554__B1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24555__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24556__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24559__B (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24559__C (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24561__B (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24562__B (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24563__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24567__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24567__B (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24569__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24572__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24573__B (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24573__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24576__A (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24588__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24589__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24595__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24596__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24604__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24607__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24613__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24616__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24622__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24622__B (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24624__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24625__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24631__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24631__B (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24633__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24634__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24643__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24643__B (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24645__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24646__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24652__A (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24652__B (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24654__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24655__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24677__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24678__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24684__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24691__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24694__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24697__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24698__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24704__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24712__B (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24713__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__24715__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24716__B (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24726__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24727__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24731__A (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24732__A1 (.DIODE(_00497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24732__A2 (.DIODE(_00500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24734__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24735__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24740__A (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24743__A (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24744__B (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24760__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24761__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24777__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24778__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24784__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24785__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24801__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24802__C (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24807__B (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24808__B (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24810__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24811__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24818__B (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24819__A (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24821__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24822__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24826__B (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24827__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__24829__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24830__B (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24834__B (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24835__A (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24837__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24838__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24853__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24854__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24870__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24871__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24876__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24877__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24891__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24892__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24896__A (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24898__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24899__A (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24901__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24902__B (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24907__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24908__A (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24910__B (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24911__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24915__B (.DIODE(_00680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24916__A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__24918__A (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24919__B (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24923__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24924__A (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24926__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24927__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24941__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24942__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24957__B (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24958__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24963__C (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24964__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24966__A (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24967__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24973__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24974__A (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24976__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24977__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24983__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24984__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24990__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24991__B (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__24993__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__24994__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25008__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25009__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25014__C (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25015__B (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25017__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25018__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25032__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25037__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25037__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25039__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25050__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25052__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25054__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25064__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25068__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25071__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25075__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25085__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25086__A2 (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25086__B1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25087__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25093__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25096__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25103__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25104__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25111__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25113__A (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25124__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25127__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25128__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25131__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25140__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25154__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25155__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25161__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25162__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25179__B (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25180__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25187__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25189__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25190__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25198__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25200__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25201__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25213__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25214__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25217__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25218__B (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25220__B1 (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25226__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25229__B (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25229__C (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25231__B (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25232__B (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25233__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25237__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25237__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25239__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25242__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25243__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25243__B (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25243__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25246__A (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25254__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25254__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25256__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25257__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25263__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25263__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25265__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25266__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25275__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25275__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25277__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25278__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25284__A (.DIODE(_01037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25284__B (.DIODE(_01039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25286__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25287__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25306__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25308__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25309__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25315__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25316__C (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25321__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25323__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25324__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25330__A (.DIODE(_01041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25331__B1 (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25332__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25344__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25356__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25357__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25365__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25366__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25378__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25379__A (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25381__A (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25385__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25386__A (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25388__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25389__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25393__B (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25402__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25403__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25409__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25410__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25420__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25421__A (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25423__A (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25426__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25427__A (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25429__A (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25430__B (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25434__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25441__A (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25442__B (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25450__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25451__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25464__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25465__A (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25467__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25468__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25474__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25475__B (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25477__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25478__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25485__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25486__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25492__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25493__B (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25495__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25496__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25509__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25510__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25515__C (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25516__B (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25518__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25519__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25532__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25537__A (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25537__B (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25539__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__25540__B (.DIODE(_01412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25541__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25545__A (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25545__B (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25547__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25548__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25549__B (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25549__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25558__A2 (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25558__B1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25559__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25560__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25563__B (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25563__C (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25565__B (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25566__C (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25581__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25582__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25589__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25590__B (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25598__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25601__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25607__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25610__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25616__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__25616__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__25618__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25619__B (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25625__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__25625__B (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25627__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25628__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25637__A (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25637__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__25639__B (.DIODE(_11105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25640__B (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25646__A (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25646__B (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25648__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25649__B (.DIODE(_11117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25667__A1 (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25670__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25675__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25676__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25681__A (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25682__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__25682__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__25684__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25685__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25687__A (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25691__A (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25694__A (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25695__B (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25700__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25704__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25719__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25720__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25725__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25726__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__25726__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__25728__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25729__B (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25734__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25735__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__25737__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25738__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25753__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25754__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25769__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25770__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25776__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25777__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25793__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25794__C (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25799__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25800__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25802__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25803__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25810__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25811__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__25813__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25814__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25818__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25819__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__25820__B1 (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25822__B (.DIODE(_06149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25827__A (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25828__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25829__A (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25831__B (.DIODE(_11185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25832__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25847__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25848__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25864__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25865__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25871__B (.DIODE(_11199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25872__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25886__B (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25887__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25892__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25893__A (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25895__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25896__B (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25902__B1 (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25903__A (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25905__B (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25906__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25910__B (.DIODE(_01725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25911__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__25913__A (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25914__B (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25919__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25920__A (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25922__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25923__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25936__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25937__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25952__B (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25953__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25958__C (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25959__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25961__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25962__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25968__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25969__A (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25971__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25972__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25979__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25980__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25986__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25987__B (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__25989__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__25990__B (.DIODE(_11376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26004__B (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26005__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26010__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26011__B (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__26013__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26014__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26027__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26032__A (.DIODE(_02128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26032__B (.DIODE(_02130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26035__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__26036__B (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__26038__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__26039__B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__26041__A0 (.DIODE(\M00r[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__26041__A1 (.DIODE(\M00r[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__26048__A (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26049__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__26049__A2 (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26054__B (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26056__B (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26058__A0 (.DIODE(\M00r[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__26059__A1 (.DIODE(\M00r[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__26061__A1 (.DIODE(\M00r[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__26063__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26072__B (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26073__A1 (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26074__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26079__B (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26084__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26100__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26102__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26104__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26137__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26139__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26142__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26192__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26193__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26194__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26196__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26198__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26249__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26250__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26251__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26252__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26253__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26255__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26314__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26315__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26316__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26317__S (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26318__S (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26320__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26385__B (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26386__A1 (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26387__S (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26388__S (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26390__B (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26391__A1 (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26392__B (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26393__A1 (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26432__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__26434__A (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26434__B (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__26439__A (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26441__A (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26441__B (.DIODE(_02146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26447__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26448__B (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26452__B (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26507__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__26508__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26509__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__26517__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__26527__A (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26527__B (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26529__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26529__B (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26530__B (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26531__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26539__B (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26608__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__26608__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__26610__A1 (.DIODE(_08790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26610__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__26610__A3 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__26610__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__26621__A (.DIODE(_02774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26621__B (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26623__A (.DIODE(_02774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26709__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__26710__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__26723__B (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26802__A (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26803__B (.DIODE(_02576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26804__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__26819__A (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26910__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__26925__A (.DIODE(_03106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26926__B (.DIODE(_03106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__26928__B_N (.DIODE(_03106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27004__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__27005__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__27017__A (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27092__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__27098__A_N (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27099__B (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27100__B (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27127__B (.DIODE(_01907_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27128__A (.DIODE(_11412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27132__A (.DIODE(_02128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27132__B (.DIODE(_02130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27134__B (.DIODE(_11421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27135__B (.DIODE(_11426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27136__B (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27136__C (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27145__A2 (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27145__B1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27146__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27147__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27150__B (.DIODE(_02128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27150__C (.DIODE(_02130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27152__B (.DIODE(_13679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27153__C (.DIODE(_11799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27168__B1 (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27172__B (.DIODE(_12047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27174__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27175__C (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27181__B (.DIODE(_02128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27181__C (.DIODE(_02130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27182__B1 (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27183__C (.DIODE(_12261_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27189__A (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27190__B (.DIODE(_12270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27203__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27204__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27208__A (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27211__B (.DIODE(_11496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27212__B (.DIODE(_11494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27225__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27226__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27232__B (.DIODE(_02130_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27232__C (.DIODE(_02128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27236__B (.DIODE(_11482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27237__C (.DIODE(_11484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27243__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27244__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27247__B (.DIODE(_12085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27248__B (.DIODE(_12087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27255__A (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27259__B (.DIODE(_12030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27260__A2 (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27260__B1 (.DIODE(_00174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27261__B (.DIODE(_12035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27264__B (.DIODE(_12043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27271__B (.DIODE(_12056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27272__C (.DIODE(_12058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27282__B (.DIODE(_13182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27284__B (.DIODE(_08176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27301__B (.DIODE(_13197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27302__B (.DIODE(_10939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27309__A (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27311__B (.DIODE(_08951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27312__C (.DIODE(_12771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27321__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27322__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27328__B (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27331__B (.DIODE(_11614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27332__B (.DIODE(_11616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27337__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27339__B (.DIODE(_12101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27341__B (.DIODE(_12008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27344__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27353__B (.DIODE(_12002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27357__B (.DIODE(_12012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27374__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27375__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27380__B (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27381__B (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27383__B (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27384__B (.DIODE(_11588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27397__B (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27400__B (.DIODE(_11600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27401__B (.DIODE(_11603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27407__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27411__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27413__B (.DIODE(_12017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27415__B (.DIODE(_11986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27430__B (.DIODE(_11983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27431__B (.DIODE(_11990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27437__B (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27438__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__27439__B1 (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27440__B (.DIODE(_12187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27453__A (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27455__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27464__B (.DIODE(_11671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27465__B (.DIODE(_12817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27479__B (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27480__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__27481__B1 (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27482__B (.DIODE(_13304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27488__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27489__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27502__B (.DIODE(_12120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27503__B (.DIODE(_12118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27509__A (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27510__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27511__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__27513__B (.DIODE(_11715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27514__B (.DIODE(_11717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27527__B (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27528__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27533__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27534__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__27536__B (.DIODE(_11701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27537__B (.DIODE(_11703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27543__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27546__B (.DIODE(_12149_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27547__B (.DIODE(_12147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27550__B (.DIODE(_11754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27564__A (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27565__B (.DIODE(_12894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27572__A (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27573__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27579__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27580__A (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27582__B (.DIODE(_06754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27583__B (.DIODE(_13502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27593__B (.DIODE(_03404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27594__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__27597__B (.DIODE(_11840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27598__B (.DIODE(_11838_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27606__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27607__B (.DIODE(_11774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27612__A (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27614__B (.DIODE(_13461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27620__A (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27621__B (.DIODE(_12914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27626__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27627__A (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27629__B (.DIODE(_13537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27630__B (.DIODE(_07400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27640__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27641__C (.DIODE(_11797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27657__A (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27658__B (.DIODE(_12939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27664__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27665__A (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27667__B (.DIODE(_11811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27668__B (.DIODE(_11808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27674__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27675__B (.DIODE(_11858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27747__A (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27748__B (.DIODE(_12992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27752__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27753__B (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27755__B (.DIODE(_11896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27756__B (.DIODE(_11899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27765__A (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27766__B (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27772__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27773__A (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27775__B (.DIODE(_08020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27776__B (.DIODE(_13022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27786__A (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27787__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27791__C (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27792__B (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27794__A (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27795__B (.DIODE(_12506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27806__A (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27807__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27812__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27813__B (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27815__B (.DIODE(_11948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27816__B (.DIODE(_11946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27823__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27835__C (.DIODE(_05167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27854__A (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__27854__B (.DIODE(_12221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27855__B (.DIODE(_04126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27857__A (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27865__B (.DIODE(_14113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27866__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27869__B (.DIODE(_13042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27870__B (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27877__B (.DIODE(_13633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27886__A (.DIODE(_02304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27905__B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__27907__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__27908__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__27908__C (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__27909__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__27910__C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__27911__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__27913__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__27913__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__27914__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__27915__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27918__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27920__A (.DIODE(_02203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27922__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__27923__C (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__27927__B1 (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27930__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__27934__A2 (.DIODE(_02162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27934__A3 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__27934__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27938__A_N (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__27939__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__27943__S (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27944__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27947__A (.DIODE(_02152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27948__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__27950__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__27953__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27957__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__27958__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__27960__C (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27962__A (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27963__A1 (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27963__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__27963__B1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27965__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__27965__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__27966__A (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27967__A2 (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27968__A (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27969__A1 (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27969__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__27971__A (.DIODE(_02155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27972__A (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27977__A (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27978__A (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27978__B (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27979__A2 (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27980__A (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27982__A2 (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27982__B1 (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27984__B (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27985__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__27986__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__27988__B (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27992__A (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27993__A (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27994__B (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27995__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__27997__A (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__27998__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__28004__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28006__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28006__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__28008__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28010__B1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28012__B (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28013__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__28014__B (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28017__A1 (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28017__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__28020__A (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28027__A2 (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28029__B (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28032__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28034__C (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28038__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28042__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28044__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28047__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__28052__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28053__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28053__C (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__28055__S (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28056__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28058__A (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28059__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__28065__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__28068__B (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28070__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28073__A (.DIODE(_04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28078__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28079__C (.DIODE(_04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28080__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28086__A2 (.DIODE(_04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28089__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28091__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28094__A (.DIODE(_04381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28100__A2 (.DIODE(_04381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28105__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28106__C (.DIODE(_04381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28107__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28109__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28114__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28117__A (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28123__A2 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28128__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28129__C (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28130__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28131__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28132__A (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28133__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28136__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28138__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28141__A (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28147__A2 (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28149__B (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28151__A (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28151__B (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28153__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28156__A (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28157__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28160__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28162__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28165__A (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28171__A2 (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28176__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28177__C (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28178__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28179__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28180__A (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28181__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28184__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28186__A (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28188__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__28190__A (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28195__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28196__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28196__C (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28199__A (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28200__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28204__A2 (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28206__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28207__B (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28212__A (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28217__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28218__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28218__C (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28222__A1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28222__B1 (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28226__A2 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28226__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28228__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28229__B (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28234__A (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28240__A2 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28242__B (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28244__A (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28244__B (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28246__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28249__A (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28250__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28253__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28258__A (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28263__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28264__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28264__C (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28266__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28267__A (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28268__A1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28268__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28272__A2 (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28275__B (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28280__A (.DIODE(_04578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28281__B (.DIODE(_04578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28284__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28285__A (.DIODE(_04578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28287__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28294__A1 (.DIODE(_04578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28294__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28297__A (.DIODE(_04578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28297__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28304__A (.DIODE(_04578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28304__C (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28305__A (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28309__A1 (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28309__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28309__B1 (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28311__A (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28312__A (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28314__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28315__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28316__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28316__B (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28317__A (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28318__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28321__A (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28321__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28326__A (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28327__A (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28328__B (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28331__A (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28332__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28336__B1 (.DIODE(_04270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28340__A1 (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28340__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28340__B1 (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28347__A (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28348__A (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28349__B (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28350__A (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28353__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28354__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28355__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28355__B (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28356__A (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28357__A1 (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28357__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28361__A1 (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28361__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__28361__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28364__A (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28364__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28369__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28374__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28375__C (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28376__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28378__A (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28378__B (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28383__A2 (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28385__B (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28395__A (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28396__C (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28397__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28404__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__28404__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28406__B (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28407__A1 (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28408__B (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28411__A (.DIODE(_04716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28416__A (.DIODE(_04183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28417__C (.DIODE(_04716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28418__C (.DIODE(_04262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28420__A (.DIODE(_04716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28425__A2 (.DIODE(_04716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28428__B (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28430__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__28438__A (.DIODE(_04258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28439__B (.DIODE(_04240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28440__A (.DIODE(_04192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28441__A (.DIODE(_04242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28442__B1 (.DIODE(_04212_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28448__B (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28449__B (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28452__A1 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28453__B (.DIODE(_04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28454__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28457__A (.DIODE(_04274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28458__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28458__C (.DIODE(_04649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28461__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28461__C (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28462__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28464__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28465__B (.DIODE(_04716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28470__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28476__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28476__C (.DIODE(_04603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28477__B (.DIODE(_04672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28479__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28480__A1 (.DIODE(_04381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28487__A (.DIODE(_04714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28495__B (.DIODE(_04457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28496__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28498__B (.DIODE(_04431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28499__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28502__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28503__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28505__B (.DIODE(_04381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28506__B (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28510__B (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28511__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28513__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__28514__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28517__B (.DIODE(_04303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28518__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28520__B (.DIODE(_04555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28521__B (.DIODE(_04766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28521__C (.DIODE(_04578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28526__A (.DIODE(_04222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28526__B (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28527__C (.DIODE(_04252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28531__B (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28532__A1 (.DIODE(_04205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28533__B (.DIODE(_04275_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28533__C (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__28536__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__28538__B (.DIODE(_04483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28539__B (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28554__A1 (.DIODE(_03296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28559__A (.DIODE(_02774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28559__B (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28560__A (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28560__B (.DIODE(_03106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28561__A (.DIODE(_03206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28561__B (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28562__A2 (.DIODE(_04876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28569__A (.DIODE(_11935_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28569__B (.DIODE(_08554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28569__C (.DIODE(_12495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28569__D (.DIODE(_09943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28570__D (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28571__B (.DIODE(_05386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28572__B (.DIODE(_05386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28574__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__28574__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__28574__C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__28574__D (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__28575__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__28575__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__28576__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__28576__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__28576__C (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__28576__D (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__28577__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__28580__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__28580__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__28580__C (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__28580__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__28582__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__28582__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__28582__C (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__28583__C (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28587__D (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28589__A (.DIODE(_05386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28590__B (.DIODE(_05386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28597__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__28597__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__28597__C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__28597__D (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__28598__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__28598__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__28598__C (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__28600__A (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28604__A (.DIODE(div_zero_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA__28608__C (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__28609__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__28610__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__28610__B (.DIODE(_04897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__28612__A (.DIODE(div_zero_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA__28613__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28613__D (.DIODE(\div1i.quot[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28613__RESET_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__28614__CLK (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28614__D (.DIODE(\div1i.quot[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28614__RESET_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__28615__CLK (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28615__D (.DIODE(\div1i.quot[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28615__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__28616__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28616__D (.DIODE(\div1i.quot[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28616__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__28617__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28617__D (.DIODE(\div1i.quot[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28617__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__28618__CLK (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28618__D (.DIODE(\div1i.quot[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28618__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__28619__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28619__D (.DIODE(\div1i.quot[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28619__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__28620__CLK (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28620__D (.DIODE(\div1i.quot[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28620__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__28621__CLK (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28621__D (.DIODE(\div1i.quot[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28621__RESET_B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__28622__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28622__D (.DIODE(\div1i.quot[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28622__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28623__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28623__D (.DIODE(\div1i.quot[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28623__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28624__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28624__D (.DIODE(\div1i.quot[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28624__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28625__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28625__D (.DIODE(\div1i.quot[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28625__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28626__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28626__D (.DIODE(\div1i.quot[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28626__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28627__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28627__D (.DIODE(\div1i.quot[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28627__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28628__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28628__D (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__28628__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28629__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28629__D (.DIODE(\div1i.quot[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28629__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28630__CLK (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28630__D (.DIODE(\div1i.quot[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28630__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28631__CLK (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28631__D (.DIODE(\div1i.quot[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28631__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__28632__CLK (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28632__D (.DIODE(\div1i.quot[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28632__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__28633__CLK (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28633__D (.DIODE(\div1i.quot[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28633__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__28634__CLK (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28634__D (.DIODE(\div1i.quot[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28634__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__28635__CLK (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28635__D (.DIODE(\div1i.quot[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28635__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__28636__CLK (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28636__D (.DIODE(\div1i.quot[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28636__RESET_B (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__28637__CLK (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28637__RESET_B (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__28638__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28639__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28639__RESET_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__28640__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28641__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28642__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28643__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28644__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28645__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28646__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28647__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28648__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28649__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28650__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28651__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28652__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28653__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28654__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28655__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28656__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28657__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28658__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28659__CLK (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28660__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28661__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28662__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28663__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28664__CLK (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28664__RESET_B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__28665__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28666__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28667__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28668__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28669__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28670__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28671__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28672__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28673__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28674__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28675__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28676__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28677__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28678__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28678__D (.DIODE(\out_f_c[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28679__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28679__D (.DIODE(\out_f_c[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__28680__CLK (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28681__CLK (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28681__D (.DIODE(div_zero_f_c));
 sky130_fd_sc_hd__diode_2 ANTENNA__28682__CLK (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__28682__D (.DIODE(forward_c));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold57_A (.DIODE(_04227_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold66_A (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold81_A (.DIODE(_04332_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold82_A (.DIODE(\M00r[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold96_A (.DIODE(\M00r[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_A (.DIODE(_06383_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer11_A (.DIODE(_07538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer12_A (.DIODE(_06383_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer16_A (.DIODE(_06385_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer41_A (.DIODE(_10009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_A (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer6_A (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer7_A (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer8_A (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer9_A (.DIODE(_06969_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split11_A (.DIODE(_01586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split14_A (.DIODE(_02112_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split1_A (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split22_A (.DIODE(\div1i.quot[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_split30_A (.DIODE(_13104_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split34_A (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split43_A (.DIODE(_07055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split5_A (.DIODE(_12974_));
 sky130_fd_sc_hd__diode_2 ANTENNA_split6_A (.DIODE(_07011_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire107_A (.DIODE(_02135_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_1551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_1514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_1466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_1319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_1519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_1435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_1443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_1550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_1486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_1456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_1445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_1512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_1229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_1507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_1432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_1508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_1552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1066 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1087 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_1529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_1541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1043 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1068 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_892 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_87 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_871 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_1363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1092 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_1238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_1322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1008 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_1341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_919 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_1287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_1549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1020 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_1553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1024 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_1383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_1516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_1364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_1500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_1520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_1495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_1503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_1506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_1522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_1545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1050 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1366 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1044 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_1334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_1442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_1498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_1544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_1298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_1488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_871 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1404 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_1541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1493 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1273 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_1407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_1524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_1532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_1499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_868 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_1532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_1519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1014 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_1509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_1521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_1497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_1522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_1508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1098 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_1521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1532 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_996 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_1354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_1513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1534 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_1503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_1525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_979 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__nor2_8 _14292_ (.A(net44),
    .B(net33),
    .Y(_05167_));
 sky130_fd_sc_hd__inv_6 _14293_ (.A(net58),
    .Y(_05178_));
 sky130_fd_sc_hd__inv_6 _14294_ (.A(net55),
    .Y(_05189_));
 sky130_fd_sc_hd__and3_4 _14295_ (.A(_05167_),
    .B(_05178_),
    .C(_05189_),
    .X(_05200_));
 sky130_fd_sc_hd__buf_6 _14296_ (.A(net60),
    .X(_05211_));
 sky130_fd_sc_hd__nor2_1 _14297_ (.A(_05211_),
    .B(net59),
    .Y(_05222_));
 sky130_fd_sc_hd__nand2_4 _14298_ (.A(_05200_),
    .B(_05222_),
    .Y(_05233_));
 sky130_fd_sc_hd__nor2_8 _14299_ (.A(net61),
    .B(_05233_),
    .Y(_05244_));
 sky130_fd_sc_hd__inv_6 _14300_ (.A(net62),
    .Y(_05255_));
 sky130_fd_sc_hd__and2_4 _14301_ (.A(_05244_),
    .B(_05255_),
    .X(_05266_));
 sky130_fd_sc_hd__buf_8 _14302_ (.A(_05266_),
    .X(_05277_));
 sky130_fd_sc_hd__clkinv_4 _14303_ (.A(net35),
    .Y(_05288_));
 sky130_fd_sc_hd__clkinv_4 _14304_ (.A(net34),
    .Y(_05299_));
 sky130_fd_sc_hd__inv_2 _14305_ (.A(net64),
    .Y(_05310_));
 sky130_fd_sc_hd__clkinv_4 _14306_ (.A(net63),
    .Y(_05321_));
 sky130_fd_sc_hd__and4_1 _14307_ (.A(_05288_),
    .B(_05299_),
    .C(_05310_),
    .D(_05321_),
    .X(_05332_));
 sky130_fd_sc_hd__nor2_1 _14308_ (.A(net37),
    .B(net36),
    .Y(_05342_));
 sky130_fd_sc_hd__nand3_4 _14309_ (.A(_05277_),
    .B(_05332_),
    .C(_05342_),
    .Y(_05353_));
 sky130_fd_sc_hd__nor2_8 _14310_ (.A(net38),
    .B(_05353_),
    .Y(_05364_));
 sky130_fd_sc_hd__inv_6 _14311_ (.A(net39),
    .Y(_05375_));
 sky130_fd_sc_hd__nand2_8 _14312_ (.A(_05364_),
    .B(_05375_),
    .Y(_05386_));
 sky130_fd_sc_hd__inv_6 _14313_ (.A(_05386_),
    .Y(_05397_));
 sky130_fd_sc_hd__clkinv_4 _14314_ (.A(net40),
    .Y(_05408_));
 sky130_fd_sc_hd__nand2_1 _14315_ (.A(_05397_),
    .B(_05408_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2_1 _14316_ (.A(_05386_),
    .B(net40),
    .Y(_05430_));
 sky130_fd_sc_hd__nand2_1 _14317_ (.A(_05419_),
    .B(_05430_),
    .Y(_05441_));
 sky130_fd_sc_hd__inv_2 _14318_ (.A(net12),
    .Y(_05452_));
 sky130_fd_sc_hd__nand2_1 _14319_ (.A(_05452_),
    .B(net44),
    .Y(_05463_));
 sky130_fd_sc_hd__inv_4 _14320_ (.A(net44),
    .Y(_05474_));
 sky130_fd_sc_hd__nand2_1 _14321_ (.A(_05474_),
    .B(net12),
    .Y(_05485_));
 sky130_fd_sc_hd__clkinv_4 _14322_ (.A(net33),
    .Y(_05496_));
 sky130_fd_sc_hd__nand2_1 _14323_ (.A(_05496_),
    .B(net1),
    .Y(_05507_));
 sky130_fd_sc_hd__nand3_1 _14324_ (.A(_05463_),
    .B(_05485_),
    .C(_05507_),
    .Y(_05518_));
 sky130_fd_sc_hd__nand2_1 _14325_ (.A(_05518_),
    .B(_05463_),
    .Y(_05529_));
 sky130_fd_sc_hd__inv_2 _14326_ (.A(net26),
    .Y(_05540_));
 sky130_fd_sc_hd__nand2_1 _14327_ (.A(_05540_),
    .B(net58),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_1 _14328_ (.A(_05178_),
    .B(net26),
    .Y(_05562_));
 sky130_fd_sc_hd__nand2_1 _14329_ (.A(_05551_),
    .B(_05562_),
    .Y(_05573_));
 sky130_fd_sc_hd__nand2_1 _14330_ (.A(_05189_),
    .B(net23),
    .Y(_05584_));
 sky130_fd_sc_hd__inv_2 _14331_ (.A(net23),
    .Y(_05595_));
 sky130_fd_sc_hd__nand2_1 _14332_ (.A(_05595_),
    .B(net55),
    .Y(_05606_));
 sky130_fd_sc_hd__nand2_1 _14333_ (.A(_05584_),
    .B(_05606_),
    .Y(_05617_));
 sky130_fd_sc_hd__nor2_1 _14334_ (.A(_05573_),
    .B(_05617_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_1 _14335_ (.A(_05529_),
    .B(_05628_),
    .Y(_05639_));
 sky130_fd_sc_hd__nor2_1 _14336_ (.A(net23),
    .B(_05189_),
    .Y(_05650_));
 sky130_fd_sc_hd__a21boi_1 _14337_ (.A1(_05650_),
    .A2(_05562_),
    .B1_N(_05551_),
    .Y(_05661_));
 sky130_fd_sc_hd__nand2_1 _14338_ (.A(_05639_),
    .B(_05661_),
    .Y(_05672_));
 sky130_fd_sc_hd__clkinvlp_2 _14339_ (.A(net27),
    .Y(_05683_));
 sky130_fd_sc_hd__nand2_1 _14340_ (.A(_05683_),
    .B(net59),
    .Y(_05694_));
 sky130_fd_sc_hd__clkinv_4 _14341_ (.A(net59),
    .Y(_05705_));
 sky130_fd_sc_hd__nand2_1 _14342_ (.A(_05705_),
    .B(net27),
    .Y(_05716_));
 sky130_fd_sc_hd__and2_1 _14343_ (.A(_05694_),
    .B(_05716_),
    .X(_05727_));
 sky130_fd_sc_hd__inv_6 _14344_ (.A(_05211_),
    .Y(_05738_));
 sky130_fd_sc_hd__nor2_1 _14345_ (.A(net28),
    .B(_05738_),
    .Y(_05749_));
 sky130_fd_sc_hd__inv_2 _14346_ (.A(net28),
    .Y(_05760_));
 sky130_fd_sc_hd__nor2_1 _14347_ (.A(_05211_),
    .B(_05760_),
    .Y(_05771_));
 sky130_fd_sc_hd__nor2_1 _14348_ (.A(_05749_),
    .B(_05771_),
    .Y(_05782_));
 sky130_fd_sc_hd__nand2_1 _14349_ (.A(_05727_),
    .B(_05782_),
    .Y(_05793_));
 sky130_fd_sc_hd__inv_2 _14350_ (.A(net30),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_1 _14351_ (.A(_05804_),
    .B(net62),
    .Y(_05815_));
 sky130_fd_sc_hd__nand2_1 _14352_ (.A(_05255_),
    .B(net30),
    .Y(_05826_));
 sky130_fd_sc_hd__nand2_1 _14353_ (.A(_05815_),
    .B(_05826_),
    .Y(_05836_));
 sky130_fd_sc_hd__inv_2 _14354_ (.A(net61),
    .Y(_05847_));
 sky130_fd_sc_hd__nand2_1 _14355_ (.A(_05847_),
    .B(net29),
    .Y(_05858_));
 sky130_fd_sc_hd__inv_2 _14356_ (.A(net29),
    .Y(_05869_));
 sky130_fd_sc_hd__nand2_1 _14357_ (.A(_05869_),
    .B(net61),
    .Y(_05880_));
 sky130_fd_sc_hd__nand2_1 _14358_ (.A(_05858_),
    .B(_05880_),
    .Y(_05891_));
 sky130_fd_sc_hd__nor2_2 _14359_ (.A(_05836_),
    .B(_05891_),
    .Y(_05902_));
 sky130_fd_sc_hd__inv_2 _14360_ (.A(_05902_),
    .Y(_05913_));
 sky130_fd_sc_hd__nor2_1 _14361_ (.A(_05793_),
    .B(_05913_),
    .Y(_05924_));
 sky130_fd_sc_hd__nand2_1 _14362_ (.A(_05672_),
    .B(_05924_),
    .Y(_05935_));
 sky130_fd_sc_hd__o21bai_1 _14363_ (.A1(_05694_),
    .A2(_05771_),
    .B1_N(_05749_),
    .Y(_05946_));
 sky130_fd_sc_hd__o21ai_1 _14364_ (.A1(_05880_),
    .A2(_05836_),
    .B1(_05815_),
    .Y(_05957_));
 sky130_fd_sc_hd__a21oi_1 _14365_ (.A1(_05946_),
    .A2(_05902_),
    .B1(_05957_),
    .Y(_05968_));
 sky130_fd_sc_hd__nand2_1 _14366_ (.A(_05935_),
    .B(_05968_),
    .Y(_05979_));
 sky130_fd_sc_hd__inv_2 _14367_ (.A(net4),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2_1 _14368_ (.A(_05990_),
    .B(net36),
    .Y(_06001_));
 sky130_fd_sc_hd__clkinv_4 _14369_ (.A(net36),
    .Y(_06012_));
 sky130_fd_sc_hd__nand2_1 _14370_ (.A(_06012_),
    .B(net4),
    .Y(_06023_));
 sky130_fd_sc_hd__and2_1 _14371_ (.A(_06001_),
    .B(_06023_),
    .X(_06034_));
 sky130_fd_sc_hd__clkinv_4 _14372_ (.A(net37),
    .Y(_06045_));
 sky130_fd_sc_hd__nor2_1 _14373_ (.A(net5),
    .B(_06045_),
    .Y(_06056_));
 sky130_fd_sc_hd__and2b_1 _14374_ (.A_N(net37),
    .B(net5),
    .X(_06067_));
 sky130_fd_sc_hd__nor2_1 _14375_ (.A(_06056_),
    .B(_06067_),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2_1 _14376_ (.A(_06034_),
    .B(_06078_),
    .Y(_06089_));
 sky130_fd_sc_hd__inv_2 _14377_ (.A(net7),
    .Y(_06100_));
 sky130_fd_sc_hd__nand2_1 _14378_ (.A(_06100_),
    .B(net39),
    .Y(_06111_));
 sky130_fd_sc_hd__nand2_1 _14379_ (.A(_05375_),
    .B(net7),
    .Y(_06122_));
 sky130_fd_sc_hd__nand2_1 _14380_ (.A(_06111_),
    .B(_06122_),
    .Y(_06133_));
 sky130_fd_sc_hd__nand2b_1 _14381_ (.A_N(net6),
    .B(net38),
    .Y(_06144_));
 sky130_fd_sc_hd__clkinv_4 _14382_ (.A(net38),
    .Y(_06155_));
 sky130_fd_sc_hd__nand2_1 _14383_ (.A(_06155_),
    .B(net6),
    .Y(_06166_));
 sky130_fd_sc_hd__nand2_1 _14384_ (.A(_06144_),
    .B(_06166_),
    .Y(_06177_));
 sky130_fd_sc_hd__nor2_1 _14385_ (.A(_06133_),
    .B(_06177_),
    .Y(_06188_));
 sky130_fd_sc_hd__nand2b_1 _14386_ (.A_N(_06089_),
    .B(_06188_),
    .Y(_06199_));
 sky130_fd_sc_hd__inv_2 _14387_ (.A(net32),
    .Y(_06210_));
 sky130_fd_sc_hd__nor2_1 _14388_ (.A(net64),
    .B(_06210_),
    .Y(_06221_));
 sky130_fd_sc_hd__inv_2 _14389_ (.A(net31),
    .Y(_06232_));
 sky130_fd_sc_hd__nand2_1 _14390_ (.A(_06232_),
    .B(net63),
    .Y(_06243_));
 sky130_fd_sc_hd__nand2_1 _14391_ (.A(_05321_),
    .B(net31),
    .Y(_06254_));
 sky130_fd_sc_hd__nand2_1 _14392_ (.A(_06243_),
    .B(_06254_),
    .Y(_06265_));
 sky130_fd_sc_hd__nand2_1 _14393_ (.A(_06210_),
    .B(net64),
    .Y(_06276_));
 sky130_fd_sc_hd__nor3b_1 _14394_ (.A(_06221_),
    .B(_06265_),
    .C_N(_06276_),
    .Y(_06287_));
 sky130_fd_sc_hd__inv_2 _14395_ (.A(net3),
    .Y(_06298_));
 sky130_fd_sc_hd__nand2_1 _14396_ (.A(_06298_),
    .B(net35),
    .Y(_06309_));
 sky130_fd_sc_hd__nand2_1 _14397_ (.A(_05288_),
    .B(net3),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_1 _14398_ (.A(_06309_),
    .B(_06320_),
    .Y(_06331_));
 sky130_fd_sc_hd__nand2_1 _14399_ (.A(_05299_),
    .B(net2),
    .Y(_06342_));
 sky130_fd_sc_hd__inv_2 _14400_ (.A(net2),
    .Y(_06353_));
 sky130_fd_sc_hd__nand2_1 _14401_ (.A(_06353_),
    .B(net34),
    .Y(_06364_));
 sky130_fd_sc_hd__nand2_1 _14402_ (.A(_06342_),
    .B(_06364_),
    .Y(_06375_));
 sky130_fd_sc_hd__nor2_1 _14403_ (.A(_06331_),
    .B(_06375_),
    .Y(_06386_));
 sky130_fd_sc_hd__nand2_1 _14404_ (.A(_06287_),
    .B(_06386_),
    .Y(_06396_));
 sky130_fd_sc_hd__nor2_2 _14405_ (.A(_06199_),
    .B(_06396_),
    .Y(_06407_));
 sky130_fd_sc_hd__nand2_1 _14406_ (.A(_05979_),
    .B(_06407_),
    .Y(_06418_));
 sky130_fd_sc_hd__o21a_1 _14407_ (.A1(_06364_),
    .A2(_06331_),
    .B1(_06309_),
    .X(_06429_));
 sky130_fd_sc_hd__o21ai_1 _14408_ (.A1(_06243_),
    .A2(_06221_),
    .B1(_06276_),
    .Y(_06440_));
 sky130_fd_sc_hd__nand2_1 _14409_ (.A(_06440_),
    .B(_06386_),
    .Y(_06451_));
 sky130_fd_sc_hd__nand2_1 _14410_ (.A(_06429_),
    .B(_06451_),
    .Y(_06462_));
 sky130_fd_sc_hd__nor2b_1 _14411_ (.A(_06089_),
    .B_N(_06188_),
    .Y(_06473_));
 sky130_fd_sc_hd__o21a_1 _14412_ (.A1(_06144_),
    .A2(_06133_),
    .B1(_06111_),
    .X(_06484_));
 sky130_fd_sc_hd__o21bai_1 _14413_ (.A1(_06001_),
    .A2(_06067_),
    .B1_N(_06056_),
    .Y(_06495_));
 sky130_fd_sc_hd__nand2_1 _14414_ (.A(_06495_),
    .B(_06188_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand2_1 _14415_ (.A(_06484_),
    .B(_06506_),
    .Y(_06517_));
 sky130_fd_sc_hd__a21oi_1 _14416_ (.A1(_06462_),
    .A2(_06473_),
    .B1(_06517_),
    .Y(_06528_));
 sky130_fd_sc_hd__nand2_1 _14417_ (.A(_06418_),
    .B(_06528_),
    .Y(_06539_));
 sky130_fd_sc_hd__clkinv_4 _14418_ (.A(net46),
    .Y(_06550_));
 sky130_fd_sc_hd__nor2_1 _14419_ (.A(net14),
    .B(_06550_),
    .Y(_06561_));
 sky130_fd_sc_hd__nand2_1 _14420_ (.A(_06550_),
    .B(net14),
    .Y(_06572_));
 sky130_fd_sc_hd__nor2b_1 _14421_ (.A(_06561_),
    .B_N(_06572_),
    .Y(_06583_));
 sky130_fd_sc_hd__clkinv_4 _14422_ (.A(net47),
    .Y(_06594_));
 sky130_fd_sc_hd__nor2_1 _14423_ (.A(net15),
    .B(_06594_),
    .Y(_06605_));
 sky130_fd_sc_hd__inv_2 _14424_ (.A(net15),
    .Y(_06616_));
 sky130_fd_sc_hd__nor2_1 _14425_ (.A(net47),
    .B(_06616_),
    .Y(_06627_));
 sky130_fd_sc_hd__nor2_1 _14426_ (.A(_06605_),
    .B(_06627_),
    .Y(_06638_));
 sky130_fd_sc_hd__buf_6 _14427_ (.A(net45),
    .X(_06649_));
 sky130_fd_sc_hd__xnor2_1 _14428_ (.A(_06649_),
    .B(net13),
    .Y(_06660_));
 sky130_fd_sc_hd__and3_1 _14429_ (.A(_06583_),
    .B(_06638_),
    .C(_06660_),
    .X(_06671_));
 sky130_fd_sc_hd__clkinvlp_2 _14430_ (.A(net11),
    .Y(_06682_));
 sky130_fd_sc_hd__nand2_1 _14431_ (.A(_06682_),
    .B(net43),
    .Y(_06693_));
 sky130_fd_sc_hd__clkinv_4 _14432_ (.A(net43),
    .Y(_06704_));
 sky130_fd_sc_hd__nand2_1 _14433_ (.A(_06704_),
    .B(net11),
    .Y(_06715_));
 sky130_fd_sc_hd__buf_6 _14434_ (.A(net42),
    .X(_06726_));
 sky130_fd_sc_hd__inv_6 _14435_ (.A(_06726_),
    .Y(_06737_));
 sky130_fd_sc_hd__nand2_1 _14436_ (.A(_06737_),
    .B(net10),
    .Y(_06748_));
 sky130_fd_sc_hd__clkinvlp_2 _14437_ (.A(net10),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_1 _14438_ (.A(_06759_),
    .B(_06726_),
    .Y(_06770_));
 sky130_fd_sc_hd__and4_1 _14439_ (.A(_06693_),
    .B(_06715_),
    .C(_06748_),
    .D(_06770_),
    .X(_06781_));
 sky130_fd_sc_hd__clkinvlp_2 _14440_ (.A(net9),
    .Y(_06792_));
 sky130_fd_sc_hd__nand2_1 _14441_ (.A(_06792_),
    .B(net41),
    .Y(_06803_));
 sky130_fd_sc_hd__clkinv_4 _14442_ (.A(net41),
    .Y(_06814_));
 sky130_fd_sc_hd__nand2_1 _14443_ (.A(_06814_),
    .B(net9),
    .Y(_06825_));
 sky130_fd_sc_hd__clkinvlp_2 _14444_ (.A(net8),
    .Y(_06836_));
 sky130_fd_sc_hd__nand2_1 _14445_ (.A(_06836_),
    .B(net40),
    .Y(_06847_));
 sky130_fd_sc_hd__nand2_1 _14446_ (.A(_05408_),
    .B(net8),
    .Y(_06858_));
 sky130_fd_sc_hd__and4_1 _14447_ (.A(_06803_),
    .B(_06825_),
    .C(_06847_),
    .D(_06858_),
    .X(_06869_));
 sky130_fd_sc_hd__and3_2 _14448_ (.A(_06671_),
    .B(_06781_),
    .C(_06869_),
    .X(_06880_));
 sky130_fd_sc_hd__nand2_1 _14449_ (.A(_06539_),
    .B(_06880_),
    .Y(_06891_));
 sky130_fd_sc_hd__nand2_1 _14450_ (.A(_06803_),
    .B(_06825_),
    .Y(_06902_));
 sky130_fd_sc_hd__o21ai_1 _14451_ (.A1(_06847_),
    .A2(_06902_),
    .B1(_06803_),
    .Y(_06913_));
 sky130_fd_sc_hd__nand2_1 _14452_ (.A(_06781_),
    .B(_06913_),
    .Y(_06924_));
 sky130_fd_sc_hd__nand2_1 _14453_ (.A(_06693_),
    .B(_06715_),
    .Y(_06935_));
 sky130_fd_sc_hd__o21a_1 _14454_ (.A1(_06770_),
    .A2(_06935_),
    .B1(_06693_),
    .X(_06946_));
 sky130_fd_sc_hd__nand2_1 _14455_ (.A(_06924_),
    .B(_06946_),
    .Y(_06957_));
 sky130_fd_sc_hd__inv_2 _14456_ (.A(net13),
    .Y(_06968_));
 sky130_fd_sc_hd__a31o_1 _14457_ (.A1(_06572_),
    .A2(_06649_),
    .A3(_06968_),
    .B1(_06561_),
    .X(_06978_));
 sky130_fd_sc_hd__a21o_1 _14458_ (.A1(_06978_),
    .A2(_06638_),
    .B1(_06605_),
    .X(_06989_));
 sky130_fd_sc_hd__a21oi_2 _14459_ (.A1(_06957_),
    .A2(_06671_),
    .B1(_06989_),
    .Y(_07000_));
 sky130_fd_sc_hd__nand2_4 _14460_ (.A(_06891_),
    .B(_07000_),
    .Y(_07011_));
 sky130_fd_sc_hd__clkinvlp_2 _14461_ (.A(net1),
    .Y(_07022_));
 sky130_fd_sc_hd__a21oi_1 _14462_ (.A1(net33),
    .A2(_07022_),
    .B1(_05518_),
    .Y(_07033_));
 sky130_fd_sc_hd__and3_1 _14463_ (.A(_05924_),
    .B(_05628_),
    .C(_07033_),
    .X(_07044_));
 sky130_fd_sc_hd__nand3_4 _14464_ (.A(_06880_),
    .B(_06407_),
    .C(_07044_),
    .Y(_07055_));
 sky130_fd_sc_hd__nand2_4 _14465_ (.A(_07011_),
    .B(_07055_),
    .Y(_07066_));
 sky130_fd_sc_hd__clkbuf_8 _14466_ (.A(_07066_),
    .X(_07077_));
 sky130_fd_sc_hd__inv_6 _14467_ (.A(_07077_),
    .Y(_07088_));
 sky130_fd_sc_hd__nor2_1 _14468_ (.A(_06836_),
    .B(_07088_),
    .Y(_07099_));
 sky130_fd_sc_hd__a21oi_1 _14469_ (.A1(net7),
    .A2(_07088_),
    .B1(_07099_),
    .Y(_07110_));
 sky130_fd_sc_hd__or2_2 _14470_ (.A(_05441_),
    .B(_07110_),
    .X(_07121_));
 sky130_fd_sc_hd__nand2_1 _14471_ (.A(_07110_),
    .B(_05441_),
    .Y(_07132_));
 sky130_fd_sc_hd__nand2_1 _14472_ (.A(_07121_),
    .B(_07132_),
    .Y(_07143_));
 sky130_fd_sc_hd__inv_2 _14473_ (.A(_07143_),
    .Y(_07154_));
 sky130_fd_sc_hd__nand2_1 _14474_ (.A(_07077_),
    .B(_05452_),
    .Y(_07165_));
 sky130_fd_sc_hd__buf_6 _14475_ (.A(_07011_),
    .X(_07176_));
 sky130_fd_sc_hd__clkbuf_4 _14476_ (.A(_07055_),
    .X(_07187_));
 sky130_fd_sc_hd__nand3_1 _14477_ (.A(_07176_),
    .B(_07022_),
    .C(_07187_),
    .Y(_07198_));
 sky130_fd_sc_hd__inv_2 _14478_ (.A(_05167_),
    .Y(_07209_));
 sky130_fd_sc_hd__nand2_1 _14479_ (.A(net44),
    .B(net33),
    .Y(_07220_));
 sky130_fd_sc_hd__nand2_2 _14480_ (.A(_07209_),
    .B(_07220_),
    .Y(_07231_));
 sky130_fd_sc_hd__inv_2 _14481_ (.A(_07231_),
    .Y(_07242_));
 sky130_fd_sc_hd__nand3_2 _14482_ (.A(_07165_),
    .B(_07198_),
    .C(_07242_),
    .Y(_07253_));
 sky130_fd_sc_hd__nand2_1 _14483_ (.A(_07077_),
    .B(net12),
    .Y(_07264_));
 sky130_fd_sc_hd__nand3_1 _14484_ (.A(_07176_),
    .B(net1),
    .C(_07187_),
    .Y(_07275_));
 sky130_fd_sc_hd__nand3_1 _14485_ (.A(_07264_),
    .B(_07275_),
    .C(_07231_),
    .Y(_07286_));
 sky130_fd_sc_hd__buf_6 _14486_ (.A(_07066_),
    .X(_07297_));
 sky130_fd_sc_hd__buf_6 _14487_ (.A(net33),
    .X(_07308_));
 sky130_fd_sc_hd__nand3_1 _14488_ (.A(_07297_),
    .B(_07308_),
    .C(net1),
    .Y(_07319_));
 sky130_fd_sc_hd__inv_2 _14489_ (.A(_07319_),
    .Y(_07330_));
 sky130_fd_sc_hd__nand3_1 _14490_ (.A(_07253_),
    .B(_07286_),
    .C(_07330_),
    .Y(_07341_));
 sky130_fd_sc_hd__nand2_1 _14491_ (.A(_07341_),
    .B(_07253_),
    .Y(_07352_));
 sky130_fd_sc_hd__nand2_1 _14492_ (.A(_07077_),
    .B(_05540_),
    .Y(_07363_));
 sky130_fd_sc_hd__nand3_1 _14493_ (.A(_07176_),
    .B(_05595_),
    .C(_07187_),
    .Y(_07374_));
 sky130_fd_sc_hd__nor2_2 _14494_ (.A(net55),
    .B(_07209_),
    .Y(_07385_));
 sky130_fd_sc_hd__or2_1 _14495_ (.A(_05178_),
    .B(_07385_),
    .X(_07396_));
 sky130_fd_sc_hd__inv_2 _14496_ (.A(_05200_),
    .Y(_07407_));
 sky130_fd_sc_hd__nand2_2 _14497_ (.A(_07396_),
    .B(_07407_),
    .Y(_07418_));
 sky130_fd_sc_hd__clkinvlp_2 _14498_ (.A(_07418_),
    .Y(_07429_));
 sky130_fd_sc_hd__nand3_1 _14499_ (.A(_07363_),
    .B(_07374_),
    .C(_07429_),
    .Y(_07440_));
 sky130_fd_sc_hd__nand2_1 _14500_ (.A(_07297_),
    .B(net26),
    .Y(_07451_));
 sky130_fd_sc_hd__nand3_1 _14501_ (.A(_07011_),
    .B(net23),
    .C(_07055_),
    .Y(_07462_));
 sky130_fd_sc_hd__nand3_1 _14502_ (.A(_07451_),
    .B(_07462_),
    .C(_07418_),
    .Y(_07473_));
 sky130_fd_sc_hd__nand2_1 _14503_ (.A(_07440_),
    .B(_07473_),
    .Y(_07484_));
 sky130_fd_sc_hd__nand2_1 _14504_ (.A(_07297_),
    .B(net23),
    .Y(_07495_));
 sky130_fd_sc_hd__nand3_1 _14505_ (.A(_07176_),
    .B(net12),
    .C(_07187_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand2_1 _14506_ (.A(_07495_),
    .B(_07506_),
    .Y(_07517_));
 sky130_fd_sc_hd__nor2_2 _14507_ (.A(_05189_),
    .B(_05167_),
    .Y(_07528_));
 sky130_fd_sc_hd__nor2_8 _14508_ (.A(_07528_),
    .B(_07385_),
    .Y(_07539_));
 sky130_fd_sc_hd__nand2_1 _14509_ (.A(_07517_),
    .B(_07539_),
    .Y(_07549_));
 sky130_fd_sc_hd__clkinv_4 _14510_ (.A(_07539_),
    .Y(_07560_));
 sky130_fd_sc_hd__nand3_1 _14511_ (.A(_07495_),
    .B(_07506_),
    .C(_07560_),
    .Y(_07571_));
 sky130_fd_sc_hd__nand2_1 _14512_ (.A(_07549_),
    .B(_07571_),
    .Y(_07582_));
 sky130_fd_sc_hd__nor2_1 _14513_ (.A(_07484_),
    .B(_07582_),
    .Y(_07593_));
 sky130_fd_sc_hd__nand2_1 _14514_ (.A(_07352_),
    .B(_07593_),
    .Y(_07604_));
 sky130_fd_sc_hd__inv_2 _14515_ (.A(_07473_),
    .Y(_07615_));
 sky130_fd_sc_hd__o21a_1 _14516_ (.A1(_07549_),
    .A2(_07615_),
    .B1(_07440_),
    .X(_07626_));
 sky130_fd_sc_hd__nand2_2 _14517_ (.A(_07604_),
    .B(_07626_),
    .Y(_07637_));
 sky130_fd_sc_hd__nand2_1 _14518_ (.A(_07066_),
    .B(_05683_),
    .Y(_07648_));
 sky130_fd_sc_hd__nand3_1 _14519_ (.A(net134),
    .B(_05540_),
    .C(net243),
    .Y(_07659_));
 sky130_fd_sc_hd__nand2_1 _14520_ (.A(_07648_),
    .B(_07659_),
    .Y(_07670_));
 sky130_fd_sc_hd__nand2_2 _14521_ (.A(_07407_),
    .B(net59),
    .Y(_07681_));
 sky130_fd_sc_hd__nand2_2 _14522_ (.A(_05200_),
    .B(_05705_),
    .Y(_07692_));
 sky130_fd_sc_hd__nand2_8 _14523_ (.A(_07681_),
    .B(_07692_),
    .Y(_07703_));
 sky130_fd_sc_hd__nand2_1 _14524_ (.A(_07670_),
    .B(_07703_),
    .Y(_07714_));
 sky130_fd_sc_hd__inv_12 _14525_ (.A(_07703_),
    .Y(_07725_));
 sky130_fd_sc_hd__nand3_2 _14526_ (.A(_07648_),
    .B(_07659_),
    .C(_07725_),
    .Y(_07736_));
 sky130_fd_sc_hd__nand2_1 _14527_ (.A(_07714_),
    .B(_07736_),
    .Y(_07747_));
 sky130_fd_sc_hd__inv_2 _14528_ (.A(_07747_),
    .Y(_07758_));
 sky130_fd_sc_hd__nand2_1 _14529_ (.A(_07066_),
    .B(net28),
    .Y(_07769_));
 sky130_fd_sc_hd__nand3_1 _14530_ (.A(net134),
    .B(net27),
    .C(_07055_),
    .Y(_07780_));
 sky130_fd_sc_hd__nand2_1 _14531_ (.A(_07769_),
    .B(_07780_),
    .Y(_07791_));
 sky130_fd_sc_hd__nand2_1 _14532_ (.A(_07692_),
    .B(_05211_),
    .Y(_07802_));
 sky130_fd_sc_hd__nand2_2 _14533_ (.A(_07802_),
    .B(_05233_),
    .Y(_07813_));
 sky130_fd_sc_hd__clkinvlp_2 _14534_ (.A(_07813_),
    .Y(_07824_));
 sky130_fd_sc_hd__nand2_1 _14535_ (.A(_07791_),
    .B(_07824_),
    .Y(_07835_));
 sky130_fd_sc_hd__nand3_1 _14536_ (.A(_07769_),
    .B(_07780_),
    .C(_07813_),
    .Y(_07846_));
 sky130_fd_sc_hd__nand2_1 _14537_ (.A(_07835_),
    .B(_07846_),
    .Y(_07857_));
 sky130_fd_sc_hd__inv_2 _14538_ (.A(_07857_),
    .Y(_07868_));
 sky130_fd_sc_hd__nand2_1 _14539_ (.A(_07758_),
    .B(_07868_),
    .Y(_07879_));
 sky130_fd_sc_hd__nand2_1 _14540_ (.A(_07066_),
    .B(_05804_),
    .Y(_07890_));
 sky130_fd_sc_hd__nor2_1 _14541_ (.A(_05255_),
    .B(_05244_),
    .Y(_07901_));
 sky130_fd_sc_hd__nor2_2 _14542_ (.A(_07901_),
    .B(_05277_),
    .Y(_07912_));
 sky130_fd_sc_hd__nand3_1 _14543_ (.A(_07011_),
    .B(_05869_),
    .C(net243),
    .Y(_07923_));
 sky130_fd_sc_hd__nand3_1 _14544_ (.A(_07890_),
    .B(_07912_),
    .C(_07923_),
    .Y(_07934_));
 sky130_fd_sc_hd__nand2_1 _14545_ (.A(_07297_),
    .B(net30),
    .Y(_07945_));
 sky130_fd_sc_hd__nand3_1 _14546_ (.A(net134),
    .B(net29),
    .C(net243),
    .Y(_07956_));
 sky130_fd_sc_hd__clkinvlp_2 _14547_ (.A(_07912_),
    .Y(_07967_));
 sky130_fd_sc_hd__nand3_1 _14548_ (.A(_07945_),
    .B(_07956_),
    .C(_07967_),
    .Y(_07978_));
 sky130_fd_sc_hd__nand2_1 _14549_ (.A(_07934_),
    .B(_07978_),
    .Y(_07989_));
 sky130_fd_sc_hd__nand2_1 _14550_ (.A(_07066_),
    .B(_05869_),
    .Y(_08000_));
 sky130_fd_sc_hd__nand3_1 _14551_ (.A(_07011_),
    .B(_05760_),
    .C(_07055_),
    .Y(_08011_));
 sky130_fd_sc_hd__nand2_1 _14552_ (.A(_08000_),
    .B(_08011_),
    .Y(_08022_));
 sky130_fd_sc_hd__nand2_1 _14553_ (.A(_05233_),
    .B(net61),
    .Y(_08033_));
 sky130_fd_sc_hd__inv_2 _14554_ (.A(_08033_),
    .Y(_08044_));
 sky130_fd_sc_hd__nor2_8 _14555_ (.A(_05244_),
    .B(_08044_),
    .Y(_08055_));
 sky130_fd_sc_hd__inv_6 _14556_ (.A(_08055_),
    .Y(_08066_));
 sky130_fd_sc_hd__nand2_1 _14557_ (.A(_08022_),
    .B(_08066_),
    .Y(_08077_));
 sky130_fd_sc_hd__nand3_2 _14558_ (.A(_08000_),
    .B(_08011_),
    .C(_08055_),
    .Y(_08088_));
 sky130_fd_sc_hd__nand2_1 _14559_ (.A(_08077_),
    .B(_08088_),
    .Y(_08099_));
 sky130_fd_sc_hd__nor2_1 _14560_ (.A(_07989_),
    .B(_08099_),
    .Y(_08109_));
 sky130_fd_sc_hd__inv_2 _14561_ (.A(_08109_),
    .Y(_08120_));
 sky130_fd_sc_hd__nor2_1 _14562_ (.A(_07879_),
    .B(_08120_),
    .Y(_08131_));
 sky130_fd_sc_hd__nand2_1 _14563_ (.A(_07637_),
    .B(_08131_),
    .Y(_08142_));
 sky130_fd_sc_hd__inv_2 _14564_ (.A(_07846_),
    .Y(_08153_));
 sky130_fd_sc_hd__o21ai_2 _14565_ (.A1(_07736_),
    .A2(_08153_),
    .B1(_07835_),
    .Y(_08164_));
 sky130_fd_sc_hd__o21ai_1 _14566_ (.A1(_08088_),
    .A2(_07989_),
    .B1(_07934_),
    .Y(_08175_));
 sky130_fd_sc_hd__a21oi_1 _14567_ (.A1(_08164_),
    .A2(_08109_),
    .B1(_08175_),
    .Y(_08186_));
 sky130_fd_sc_hd__nand2_4 _14568_ (.A(_08142_),
    .B(_08186_),
    .Y(_08197_));
 sky130_fd_sc_hd__nand2_1 _14569_ (.A(_07297_),
    .B(_05990_),
    .Y(_08208_));
 sky130_fd_sc_hd__nand3_1 _14570_ (.A(net134),
    .B(_06298_),
    .C(net243),
    .Y(_08219_));
 sky130_fd_sc_hd__nand2_1 _14571_ (.A(_08208_),
    .B(_08219_),
    .Y(_08230_));
 sky130_fd_sc_hd__nand2_4 _14572_ (.A(_05277_),
    .B(_05332_),
    .Y(_08241_));
 sky130_fd_sc_hd__or2_4 _14573_ (.A(net36),
    .B(_08241_),
    .X(_08252_));
 sky130_fd_sc_hd__nand2_1 _14574_ (.A(_08241_),
    .B(net36),
    .Y(_08263_));
 sky130_fd_sc_hd__nand2_4 _14575_ (.A(_08252_),
    .B(_08263_),
    .Y(_08274_));
 sky130_fd_sc_hd__nand2_1 _14576_ (.A(_08230_),
    .B(_08274_),
    .Y(_08285_));
 sky130_fd_sc_hd__clkinv_4 _14577_ (.A(_08274_),
    .Y(_08296_));
 sky130_fd_sc_hd__nand3_2 _14578_ (.A(_08208_),
    .B(_08219_),
    .C(_08296_),
    .Y(_08307_));
 sky130_fd_sc_hd__nand2_1 _14579_ (.A(_08285_),
    .B(_08307_),
    .Y(_08318_));
 sky130_fd_sc_hd__nand2_1 _14580_ (.A(_07297_),
    .B(net5),
    .Y(_08329_));
 sky130_fd_sc_hd__nand3_1 _14581_ (.A(_07176_),
    .B(net4),
    .C(_07187_),
    .Y(_08340_));
 sky130_fd_sc_hd__nand2_1 _14582_ (.A(_08329_),
    .B(_08340_),
    .Y(_08351_));
 sky130_fd_sc_hd__nand2_1 _14583_ (.A(_08252_),
    .B(net37),
    .Y(_08362_));
 sky130_fd_sc_hd__nand2_2 _14584_ (.A(_08362_),
    .B(_05353_),
    .Y(_08373_));
 sky130_fd_sc_hd__clkinv_4 _14585_ (.A(_08373_),
    .Y(_08384_));
 sky130_fd_sc_hd__nand2_1 _14586_ (.A(_08351_),
    .B(_08384_),
    .Y(_08395_));
 sky130_fd_sc_hd__buf_6 _14587_ (.A(_08373_),
    .X(_08406_));
 sky130_fd_sc_hd__nand3_1 _14588_ (.A(_08329_),
    .B(_08340_),
    .C(_08406_),
    .Y(_08417_));
 sky130_fd_sc_hd__nand2_2 _14589_ (.A(_08395_),
    .B(_08417_),
    .Y(_08428_));
 sky130_fd_sc_hd__nor2_1 _14590_ (.A(_08318_),
    .B(_08428_),
    .Y(_08439_));
 sky130_fd_sc_hd__nand2_1 _14591_ (.A(_07297_),
    .B(net6),
    .Y(_08450_));
 sky130_fd_sc_hd__nand3_1 _14592_ (.A(net134),
    .B(net5),
    .C(net243),
    .Y(_08461_));
 sky130_fd_sc_hd__nand2_1 _14593_ (.A(_08450_),
    .B(_08461_),
    .Y(_08472_));
 sky130_fd_sc_hd__nand2_1 _14594_ (.A(_05353_),
    .B(net38),
    .Y(_08483_));
 sky130_fd_sc_hd__inv_2 _14595_ (.A(_08483_),
    .Y(_08494_));
 sky130_fd_sc_hd__nor2_8 _14596_ (.A(_05364_),
    .B(_08494_),
    .Y(_08505_));
 sky130_fd_sc_hd__nand2_1 _14597_ (.A(_08472_),
    .B(_08505_),
    .Y(_08516_));
 sky130_fd_sc_hd__clkinv_4 _14598_ (.A(_08505_),
    .Y(_08527_));
 sky130_fd_sc_hd__nand3_1 _14599_ (.A(_08450_),
    .B(_08461_),
    .C(_08527_),
    .Y(_08538_));
 sky130_fd_sc_hd__nand2_1 _14600_ (.A(_08516_),
    .B(_08538_),
    .Y(_08549_));
 sky130_fd_sc_hd__nor2_1 _14601_ (.A(_05375_),
    .B(_05364_),
    .Y(_08560_));
 sky130_fd_sc_hd__nor2_4 _14602_ (.A(_08560_),
    .B(_05397_),
    .Y(_08571_));
 sky130_fd_sc_hd__inv_6 _14603_ (.A(_08571_),
    .Y(_08582_));
 sky130_fd_sc_hd__nand2_1 _14604_ (.A(_07297_),
    .B(net7),
    .Y(_08593_));
 sky130_fd_sc_hd__nand3_1 _14605_ (.A(_07176_),
    .B(net6),
    .C(_07187_),
    .Y(_08604_));
 sky130_fd_sc_hd__nand3_1 _14606_ (.A(_08582_),
    .B(_08593_),
    .C(_08604_),
    .Y(_08615_));
 sky130_fd_sc_hd__nand2_1 _14607_ (.A(_08593_),
    .B(_08604_),
    .Y(_08626_));
 sky130_fd_sc_hd__nand2_2 _14608_ (.A(_08626_),
    .B(_08571_),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_2 _14609_ (.A(_08615_),
    .B(_08637_),
    .Y(_08647_));
 sky130_fd_sc_hd__nor2_2 _14610_ (.A(_08549_),
    .B(_08647_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand2_1 _14611_ (.A(_08439_),
    .B(_08658_),
    .Y(_08669_));
 sky130_fd_sc_hd__nand2_1 _14612_ (.A(_07077_),
    .B(net32),
    .Y(_08680_));
 sky130_fd_sc_hd__nand3_1 _14613_ (.A(_07176_),
    .B(net31),
    .C(_07187_),
    .Y(_08691_));
 sky130_fd_sc_hd__nand2_2 _14614_ (.A(_05277_),
    .B(_05321_),
    .Y(_08702_));
 sky130_fd_sc_hd__inv_6 _14615_ (.A(_08702_),
    .Y(_08713_));
 sky130_fd_sc_hd__nand2_1 _14616_ (.A(_08713_),
    .B(_05310_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand2_1 _14617_ (.A(_08702_),
    .B(net64),
    .Y(_08735_));
 sky130_fd_sc_hd__nand2_4 _14618_ (.A(_08724_),
    .B(_08735_),
    .Y(_08746_));
 sky130_fd_sc_hd__a21o_1 _14619_ (.A1(_08680_),
    .A2(_08691_),
    .B1(_08746_),
    .X(_08757_));
 sky130_fd_sc_hd__nand3_1 _14620_ (.A(_08680_),
    .B(_08691_),
    .C(_08746_),
    .Y(_08768_));
 sky130_fd_sc_hd__nand2_1 _14621_ (.A(_08757_),
    .B(_08768_),
    .Y(_08779_));
 sky130_fd_sc_hd__buf_6 _14622_ (.A(_07297_),
    .X(_08790_));
 sky130_fd_sc_hd__nand2_1 _14623_ (.A(_08790_),
    .B(_06232_),
    .Y(_08801_));
 sky130_fd_sc_hd__nand3_1 _14624_ (.A(_07176_),
    .B(_05804_),
    .C(_07187_),
    .Y(_08812_));
 sky130_fd_sc_hd__nor2_2 _14625_ (.A(_05321_),
    .B(_05277_),
    .Y(_08823_));
 sky130_fd_sc_hd__nor2_8 _14626_ (.A(_08823_),
    .B(_08713_),
    .Y(_08834_));
 sky130_fd_sc_hd__a21o_1 _14627_ (.A1(_08801_),
    .A2(_08812_),
    .B1(_08834_),
    .X(_08845_));
 sky130_fd_sc_hd__nand3_2 _14628_ (.A(_08801_),
    .B(_08812_),
    .C(_08834_),
    .Y(_08856_));
 sky130_fd_sc_hd__nand2_1 _14629_ (.A(_08845_),
    .B(_08856_),
    .Y(_08867_));
 sky130_fd_sc_hd__nor2_1 _14630_ (.A(_08779_),
    .B(_08867_),
    .Y(_08878_));
 sky130_fd_sc_hd__nand2_1 _14631_ (.A(_07297_),
    .B(_06298_),
    .Y(_08889_));
 sky130_fd_sc_hd__nand3_1 _14632_ (.A(_07176_),
    .B(_06353_),
    .C(_07187_),
    .Y(_08900_));
 sky130_fd_sc_hd__nand2_1 _14633_ (.A(_08889_),
    .B(_08900_),
    .Y(_08911_));
 sky130_fd_sc_hd__nand3_2 _14634_ (.A(_08713_),
    .B(_05299_),
    .C(_05310_),
    .Y(_08922_));
 sky130_fd_sc_hd__nand2_4 _14635_ (.A(_08922_),
    .B(net35),
    .Y(_08933_));
 sky130_fd_sc_hd__nand2_8 _14636_ (.A(_08933_),
    .B(_08241_),
    .Y(_08944_));
 sky130_fd_sc_hd__nand2_1 _14637_ (.A(_08911_),
    .B(_08944_),
    .Y(_08955_));
 sky130_fd_sc_hd__inv_6 _14638_ (.A(_08944_),
    .Y(_08966_));
 sky130_fd_sc_hd__nand3_2 _14639_ (.A(_08889_),
    .B(_08966_),
    .C(_08900_),
    .Y(_08977_));
 sky130_fd_sc_hd__nand2_1 _14640_ (.A(_08955_),
    .B(_08977_),
    .Y(_08988_));
 sky130_fd_sc_hd__nand2_1 _14641_ (.A(_08790_),
    .B(_06353_),
    .Y(_08999_));
 sky130_fd_sc_hd__nand3_1 _14642_ (.A(_07176_),
    .B(_06210_),
    .C(_07187_),
    .Y(_09010_));
 sky130_fd_sc_hd__nand2_1 _14643_ (.A(_08999_),
    .B(_09010_),
    .Y(_09021_));
 sky130_fd_sc_hd__nand2_1 _14644_ (.A(_08724_),
    .B(net34),
    .Y(_09032_));
 sky130_fd_sc_hd__nand2_2 _14645_ (.A(_09032_),
    .B(_08922_),
    .Y(_09043_));
 sky130_fd_sc_hd__buf_6 _14646_ (.A(_09043_),
    .X(_09054_));
 sky130_fd_sc_hd__nand2_1 _14647_ (.A(_09021_),
    .B(_09054_),
    .Y(_09065_));
 sky130_fd_sc_hd__clkinv_4 _14648_ (.A(_09043_),
    .Y(_09076_));
 sky130_fd_sc_hd__nand3_4 _14649_ (.A(_08999_),
    .B(_09010_),
    .C(_09076_),
    .Y(_09087_));
 sky130_fd_sc_hd__nand2_2 _14650_ (.A(_09065_),
    .B(_09087_),
    .Y(_09098_));
 sky130_fd_sc_hd__nor2_1 _14651_ (.A(_08988_),
    .B(_09098_),
    .Y(_09109_));
 sky130_fd_sc_hd__nand2_1 _14652_ (.A(_08878_),
    .B(_09109_),
    .Y(_09120_));
 sky130_fd_sc_hd__nor2_1 _14653_ (.A(_08669_),
    .B(_09120_),
    .Y(_09131_));
 sky130_fd_sc_hd__nand2_1 _14654_ (.A(_08197_),
    .B(_09131_),
    .Y(_09142_));
 sky130_fd_sc_hd__inv_2 _14655_ (.A(_08768_),
    .Y(_09153_));
 sky130_fd_sc_hd__o21ai_2 _14656_ (.A1(_08856_),
    .A2(_09153_),
    .B1(_08757_),
    .Y(_09164_));
 sky130_fd_sc_hd__nand2_1 _14657_ (.A(_09164_),
    .B(_09109_),
    .Y(_09175_));
 sky130_fd_sc_hd__inv_2 _14658_ (.A(_08955_),
    .Y(_09186_));
 sky130_fd_sc_hd__o21a_1 _14659_ (.A1(_09087_),
    .A2(_09186_),
    .B1(_08977_),
    .X(_09197_));
 sky130_fd_sc_hd__nand2_1 _14660_ (.A(_09175_),
    .B(_09197_),
    .Y(_09207_));
 sky130_fd_sc_hd__inv_2 _14661_ (.A(_08669_),
    .Y(_09218_));
 sky130_fd_sc_hd__o21a_1 _14662_ (.A1(_08516_),
    .A2(_08647_),
    .B1(_08637_),
    .X(_09229_));
 sky130_fd_sc_hd__inv_2 _14663_ (.A(_08417_),
    .Y(_09240_));
 sky130_fd_sc_hd__o21ai_1 _14664_ (.A1(_08307_),
    .A2(_09240_),
    .B1(_08395_),
    .Y(_09251_));
 sky130_fd_sc_hd__nand2_1 _14665_ (.A(_09251_),
    .B(_08658_),
    .Y(_09262_));
 sky130_fd_sc_hd__nand2_1 _14666_ (.A(_09229_),
    .B(_09262_),
    .Y(_09273_));
 sky130_fd_sc_hd__a21oi_2 _14667_ (.A1(_09207_),
    .A2(_09218_),
    .B1(_09273_),
    .Y(_09284_));
 sky130_fd_sc_hd__nand2_2 _14668_ (.A(_09142_),
    .B(_09284_),
    .Y(_09295_));
 sky130_fd_sc_hd__or2_1 _14669_ (.A(_07154_),
    .B(_09295_),
    .X(_09306_));
 sky130_fd_sc_hd__nand2_1 _14670_ (.A(_09295_),
    .B(_07154_),
    .Y(_09317_));
 sky130_fd_sc_hd__nand2_1 _14671_ (.A(_09306_),
    .B(_09317_),
    .Y(_09328_));
 sky130_fd_sc_hd__nand2_2 _14672_ (.A(_05419_),
    .B(net41),
    .Y(_09339_));
 sky130_fd_sc_hd__nand3_4 _14673_ (.A(_05397_),
    .B(_06814_),
    .C(_05408_),
    .Y(_09350_));
 sky130_fd_sc_hd__nand2_8 _14674_ (.A(_09339_),
    .B(_09350_),
    .Y(_09361_));
 sky130_fd_sc_hd__nand2_1 _14675_ (.A(_09328_),
    .B(_09361_),
    .Y(_09372_));
 sky130_fd_sc_hd__inv_6 _14676_ (.A(_09361_),
    .Y(_09383_));
 sky130_fd_sc_hd__nand3_1 _14677_ (.A(_09306_),
    .B(_09383_),
    .C(_09317_),
    .Y(_09394_));
 sky130_fd_sc_hd__nand2_1 _14678_ (.A(_09372_),
    .B(_09394_),
    .Y(_09405_));
 sky130_fd_sc_hd__inv_2 _14679_ (.A(_09120_),
    .Y(_09416_));
 sky130_fd_sc_hd__nand2_1 _14680_ (.A(_08197_),
    .B(_09416_),
    .Y(_09427_));
 sky130_fd_sc_hd__inv_2 _14681_ (.A(_09207_),
    .Y(_09438_));
 sky130_fd_sc_hd__nand2_1 _14682_ (.A(_09427_),
    .B(_09438_),
    .Y(_09449_));
 sky130_fd_sc_hd__nand2_1 _14683_ (.A(_09449_),
    .B(_08439_),
    .Y(_09460_));
 sky130_fd_sc_hd__inv_2 _14684_ (.A(_09251_),
    .Y(_09471_));
 sky130_fd_sc_hd__nand2_1 _14685_ (.A(_09460_),
    .B(_09471_),
    .Y(_09482_));
 sky130_fd_sc_hd__clkinvlp_2 _14686_ (.A(_08549_),
    .Y(_09493_));
 sky130_fd_sc_hd__nand2_1 _14687_ (.A(_09482_),
    .B(_09493_),
    .Y(_09504_));
 sky130_fd_sc_hd__nand2_1 _14688_ (.A(_09504_),
    .B(_08516_),
    .Y(_09515_));
 sky130_fd_sc_hd__inv_2 _14689_ (.A(_08647_),
    .Y(_09526_));
 sky130_fd_sc_hd__nand2_1 _14690_ (.A(_09515_),
    .B(_09526_),
    .Y(_09537_));
 sky130_fd_sc_hd__buf_6 _14691_ (.A(_05441_),
    .X(_09548_));
 sky130_fd_sc_hd__inv_2 _14692_ (.A(_09548_),
    .Y(_09559_));
 sky130_fd_sc_hd__nand3_1 _14693_ (.A(_09504_),
    .B(_08647_),
    .C(_08516_),
    .Y(_09570_));
 sky130_fd_sc_hd__nand3_2 _14694_ (.A(_09537_),
    .B(_09559_),
    .C(_09570_),
    .Y(_09581_));
 sky130_fd_sc_hd__o21ai_1 _14695_ (.A1(_09405_),
    .A2(_09581_),
    .B1(_09394_),
    .Y(_09592_));
 sky130_fd_sc_hd__mux2_1 _14696_ (.A0(net8),
    .A1(net9),
    .S(_07077_),
    .X(_09603_));
 sky130_fd_sc_hd__nand2_1 _14697_ (.A(_09603_),
    .B(_09383_),
    .Y(_09614_));
 sky130_fd_sc_hd__mux2_1 _14698_ (.A0(_06836_),
    .A1(_06792_),
    .S(_07077_),
    .X(_09625_));
 sky130_fd_sc_hd__nand2_1 _14699_ (.A(_09625_),
    .B(_09361_),
    .Y(_09636_));
 sky130_fd_sc_hd__nand2_2 _14700_ (.A(_09614_),
    .B(_09636_),
    .Y(_09647_));
 sky130_fd_sc_hd__a21o_1 _14701_ (.A1(_09317_),
    .A2(_07121_),
    .B1(_09647_),
    .X(_09658_));
 sky130_fd_sc_hd__nand3_1 _14702_ (.A(_09317_),
    .B(_09647_),
    .C(_07121_),
    .Y(_09669_));
 sky130_fd_sc_hd__nand2_1 _14703_ (.A(_09658_),
    .B(_09669_),
    .Y(_09680_));
 sky130_fd_sc_hd__nor2_4 _14704_ (.A(_06726_),
    .B(_09350_),
    .Y(_09691_));
 sky130_fd_sc_hd__nand2_2 _14705_ (.A(_09350_),
    .B(_06726_),
    .Y(_09702_));
 sky130_fd_sc_hd__inv_2 _14706_ (.A(_09702_),
    .Y(_09713_));
 sky130_fd_sc_hd__nor2_8 _14707_ (.A(_09691_),
    .B(_09713_),
    .Y(_09724_));
 sky130_fd_sc_hd__inv_6 _14708_ (.A(_09724_),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_1 _14709_ (.A(_09680_),
    .B(_09735_),
    .Y(_09745_));
 sky130_fd_sc_hd__nand3_2 _14710_ (.A(_09658_),
    .B(_09724_),
    .C(_09669_),
    .Y(_09756_));
 sky130_fd_sc_hd__nand2_1 _14711_ (.A(_09745_),
    .B(_09756_),
    .Y(_09767_));
 sky130_fd_sc_hd__mux2_1 _14712_ (.A0(_06792_),
    .A1(_06759_),
    .S(_08790_),
    .X(_09778_));
 sky130_fd_sc_hd__nand2_1 _14713_ (.A(_09778_),
    .B(_09735_),
    .Y(_09789_));
 sky130_fd_sc_hd__mux2_1 _14714_ (.A0(net9),
    .A1(net10),
    .S(_07077_),
    .X(_09800_));
 sky130_fd_sc_hd__nand2_2 _14715_ (.A(_09800_),
    .B(_09724_),
    .Y(_09811_));
 sky130_fd_sc_hd__nand2_2 _14716_ (.A(_09789_),
    .B(_09811_),
    .Y(_09822_));
 sky130_fd_sc_hd__inv_2 _14717_ (.A(_09822_),
    .Y(_09833_));
 sky130_fd_sc_hd__nor2_1 _14718_ (.A(_07143_),
    .B(_09647_),
    .Y(_09844_));
 sky130_fd_sc_hd__nand2_1 _14719_ (.A(_09295_),
    .B(_09844_),
    .Y(_09855_));
 sky130_fd_sc_hd__o21ai_2 _14720_ (.A1(_07121_),
    .A2(_09647_),
    .B1(_09614_),
    .Y(_09866_));
 sky130_fd_sc_hd__inv_2 _14721_ (.A(_09866_),
    .Y(_09877_));
 sky130_fd_sc_hd__nand2_1 _14722_ (.A(_09855_),
    .B(_09877_),
    .Y(_09888_));
 sky130_fd_sc_hd__or2_4 _14723_ (.A(_09833_),
    .B(_09888_),
    .X(_09899_));
 sky130_fd_sc_hd__nand2_2 _14724_ (.A(_09888_),
    .B(_09833_),
    .Y(_09910_));
 sky130_fd_sc_hd__nand2_2 _14725_ (.A(_09899_),
    .B(_09910_),
    .Y(_09921_));
 sky130_fd_sc_hd__o21ai_2 _14726_ (.A1(_06726_),
    .A2(_09350_),
    .B1(net43),
    .Y(_09932_));
 sky130_fd_sc_hd__or4_4 _14727_ (.A(net43),
    .B(_06726_),
    .C(net41),
    .D(net40),
    .X(_09943_));
 sky130_fd_sc_hd__nor2_1 _14728_ (.A(_09943_),
    .B(_05386_),
    .Y(_09954_));
 sky130_fd_sc_hd__inv_4 _14729_ (.A(_09954_),
    .Y(_09965_));
 sky130_fd_sc_hd__nand2_2 _14730_ (.A(_09932_),
    .B(_09965_),
    .Y(_09976_));
 sky130_fd_sc_hd__buf_6 _14731_ (.A(_09976_),
    .X(_09987_));
 sky130_fd_sc_hd__nand2_1 _14732_ (.A(_09921_),
    .B(_09987_),
    .Y(_09998_));
 sky130_fd_sc_hd__inv_6 _14733_ (.A(_09976_),
    .Y(_10009_));
 sky130_fd_sc_hd__nand3_1 _14734_ (.A(_09899_),
    .B(_10009_),
    .C(_09910_),
    .Y(_10020_));
 sky130_fd_sc_hd__nand2_1 _14735_ (.A(_09998_),
    .B(_10020_),
    .Y(_10031_));
 sky130_fd_sc_hd__nor2_1 _14736_ (.A(_09767_),
    .B(_10031_),
    .Y(_10042_));
 sky130_fd_sc_hd__nand2_1 _14737_ (.A(_09592_),
    .B(_10042_),
    .Y(_10053_));
 sky130_fd_sc_hd__inv_2 _14738_ (.A(_09756_),
    .Y(_10064_));
 sky130_fd_sc_hd__a21boi_1 _14739_ (.A1(_09998_),
    .A2(_10064_),
    .B1_N(_10020_),
    .Y(_10075_));
 sky130_fd_sc_hd__nand2_1 _14740_ (.A(_10053_),
    .B(_10075_),
    .Y(_10086_));
 sky130_fd_sc_hd__nand2_1 _14741_ (.A(_09910_),
    .B(_09811_),
    .Y(_10097_));
 sky130_fd_sc_hd__mux2_1 _14742_ (.A0(net10),
    .A1(net11),
    .S(_07077_),
    .X(_10108_));
 sky130_fd_sc_hd__nand2_2 _14743_ (.A(_10108_),
    .B(_10009_),
    .Y(_10119_));
 sky130_fd_sc_hd__mux2_1 _14744_ (.A0(_06759_),
    .A1(_06682_),
    .S(_07077_),
    .X(_10130_));
 sky130_fd_sc_hd__nand2_1 _14745_ (.A(_10130_),
    .B(_09976_),
    .Y(_10141_));
 sky130_fd_sc_hd__nand2_4 _14746_ (.A(_10119_),
    .B(_10141_),
    .Y(_10152_));
 sky130_fd_sc_hd__inv_2 _14747_ (.A(_10152_),
    .Y(_10163_));
 sky130_fd_sc_hd__nand2_1 _14748_ (.A(_10097_),
    .B(_10163_),
    .Y(_10174_));
 sky130_fd_sc_hd__nand3_1 _14749_ (.A(_09910_),
    .B(_10152_),
    .C(_09811_),
    .Y(_10185_));
 sky130_fd_sc_hd__nand2_1 _14750_ (.A(_10174_),
    .B(_10185_),
    .Y(_10196_));
 sky130_fd_sc_hd__nor2_2 _14751_ (.A(_06649_),
    .B(_09965_),
    .Y(_10207_));
 sky130_fd_sc_hd__nand2_1 _14752_ (.A(_09965_),
    .B(_06649_),
    .Y(_10218_));
 sky130_fd_sc_hd__inv_2 _14753_ (.A(_10218_),
    .Y(_10229_));
 sky130_fd_sc_hd__nor2_4 _14754_ (.A(_10207_),
    .B(_10229_),
    .Y(_10240_));
 sky130_fd_sc_hd__inv_2 _14755_ (.A(_10240_),
    .Y(_10251_));
 sky130_fd_sc_hd__nand2_1 _14756_ (.A(_10196_),
    .B(_10251_),
    .Y(_10262_));
 sky130_fd_sc_hd__nor2_4 _14757_ (.A(_09822_),
    .B(_10152_),
    .Y(_10273_));
 sky130_fd_sc_hd__and2_1 _14758_ (.A(_10273_),
    .B(_09844_),
    .X(_10284_));
 sky130_fd_sc_hd__nand2_2 _14759_ (.A(_09295_),
    .B(_10284_),
    .Y(_10295_));
 sky130_fd_sc_hd__o21ai_1 _14760_ (.A1(_09811_),
    .A2(_10152_),
    .B1(_10119_),
    .Y(_10305_));
 sky130_fd_sc_hd__a21oi_2 _14761_ (.A1(_09866_),
    .A2(_10273_),
    .B1(_10305_),
    .Y(_10316_));
 sky130_fd_sc_hd__nand2_2 _14762_ (.A(_10295_),
    .B(_10316_),
    .Y(_10327_));
 sky130_fd_sc_hd__mux2_1 _14763_ (.A0(net11),
    .A1(net13),
    .S(_08790_),
    .X(_10338_));
 sky130_fd_sc_hd__or2_1 _14764_ (.A(_10240_),
    .B(_10338_),
    .X(_10349_));
 sky130_fd_sc_hd__nand2_2 _14765_ (.A(_10338_),
    .B(_10240_),
    .Y(_10360_));
 sky130_fd_sc_hd__nand2_1 _14766_ (.A(_10349_),
    .B(_10360_),
    .Y(_10371_));
 sky130_fd_sc_hd__clkinvlp_2 _14767_ (.A(_10371_),
    .Y(_10382_));
 sky130_fd_sc_hd__nand2_2 _14768_ (.A(_10327_),
    .B(_10382_),
    .Y(_10393_));
 sky130_fd_sc_hd__nand3_1 _14769_ (.A(_10295_),
    .B(_10316_),
    .C(_10371_),
    .Y(_10404_));
 sky130_fd_sc_hd__nand2_1 _14770_ (.A(_10393_),
    .B(_10404_),
    .Y(_10415_));
 sky130_fd_sc_hd__inv_2 _14771_ (.A(_06649_),
    .Y(_10426_));
 sky130_fd_sc_hd__nand2_1 _14772_ (.A(_10426_),
    .B(_06550_),
    .Y(_10437_));
 sky130_fd_sc_hd__nor2_2 _14773_ (.A(_10437_),
    .B(_09965_),
    .Y(_10448_));
 sky130_fd_sc_hd__nor2_1 _14774_ (.A(_06550_),
    .B(_10207_),
    .Y(_10459_));
 sky130_fd_sc_hd__nor2_4 _14775_ (.A(_10448_),
    .B(_10459_),
    .Y(_10470_));
 sky130_fd_sc_hd__inv_2 _14776_ (.A(_10470_),
    .Y(_10481_));
 sky130_fd_sc_hd__nand2_1 _14777_ (.A(_10415_),
    .B(_10481_),
    .Y(_10492_));
 sky130_fd_sc_hd__nand3_1 _14778_ (.A(_10393_),
    .B(_10470_),
    .C(_10404_),
    .Y(_10503_));
 sky130_fd_sc_hd__nand2_1 _14779_ (.A(_10492_),
    .B(_10503_),
    .Y(_10514_));
 sky130_fd_sc_hd__inv_2 _14780_ (.A(_10514_),
    .Y(_10525_));
 sky130_fd_sc_hd__nand3_2 _14781_ (.A(_10174_),
    .B(_10240_),
    .C(_10185_),
    .Y(_10536_));
 sky130_fd_sc_hd__nand3_2 _14782_ (.A(_10262_),
    .B(_10525_),
    .C(_10536_),
    .Y(_10547_));
 sky130_fd_sc_hd__nand2_1 _14783_ (.A(_10393_),
    .B(_10360_),
    .Y(_10558_));
 sky130_fd_sc_hd__mux2_1 _14784_ (.A0(net13),
    .A1(net14),
    .S(_08790_),
    .X(_10569_));
 sky130_fd_sc_hd__or2_1 _14785_ (.A(_10470_),
    .B(_10569_),
    .X(_10580_));
 sky130_fd_sc_hd__nand2_1 _14786_ (.A(_10569_),
    .B(_10470_),
    .Y(_10591_));
 sky130_fd_sc_hd__nand2_1 _14787_ (.A(_10580_),
    .B(_10591_),
    .Y(_10602_));
 sky130_fd_sc_hd__clkinvlp_2 _14788_ (.A(_10602_),
    .Y(_10613_));
 sky130_fd_sc_hd__nand2_1 _14789_ (.A(_10558_),
    .B(_10613_),
    .Y(_10624_));
 sky130_fd_sc_hd__nand3_2 _14790_ (.A(_10393_),
    .B(_10602_),
    .C(_10360_),
    .Y(_10635_));
 sky130_fd_sc_hd__nand2_1 _14791_ (.A(_10624_),
    .B(_10635_),
    .Y(_10646_));
 sky130_fd_sc_hd__nor2_1 _14792_ (.A(_06594_),
    .B(_10448_),
    .Y(_10657_));
 sky130_fd_sc_hd__nand2_2 _14793_ (.A(_10448_),
    .B(_06594_),
    .Y(_10668_));
 sky130_fd_sc_hd__inv_4 _14794_ (.A(_10668_),
    .Y(_10679_));
 sky130_fd_sc_hd__nor2_4 _14795_ (.A(_10657_),
    .B(_10679_),
    .Y(_10690_));
 sky130_fd_sc_hd__clkinv_4 _14796_ (.A(_10690_),
    .Y(_10701_));
 sky130_fd_sc_hd__nand2_1 _14797_ (.A(_10646_),
    .B(_10701_),
    .Y(_10712_));
 sky130_fd_sc_hd__nand3_2 _14798_ (.A(_10624_),
    .B(_10690_),
    .C(_10635_),
    .Y(_10723_));
 sky130_fd_sc_hd__nand2_2 _14799_ (.A(_10712_),
    .B(_10723_),
    .Y(_10734_));
 sky130_fd_sc_hd__inv_2 _14800_ (.A(_10734_),
    .Y(_10745_));
 sky130_fd_sc_hd__nor2_1 _14801_ (.A(_10371_),
    .B(_10602_),
    .Y(_10756_));
 sky130_fd_sc_hd__nand2_2 _14802_ (.A(_10327_),
    .B(_10756_),
    .Y(_10767_));
 sky130_fd_sc_hd__o21a_1 _14803_ (.A1(_10360_),
    .A2(_10602_),
    .B1(_10591_),
    .X(_10778_));
 sky130_fd_sc_hd__nand2_1 _14804_ (.A(_10767_),
    .B(_10778_),
    .Y(_10789_));
 sky130_fd_sc_hd__mux2_1 _14805_ (.A0(net14),
    .A1(net15),
    .S(_08790_),
    .X(_10800_));
 sky130_fd_sc_hd__or2_1 _14806_ (.A(_10690_),
    .B(_10800_),
    .X(_10811_));
 sky130_fd_sc_hd__nand2_1 _14807_ (.A(_10800_),
    .B(_10690_),
    .Y(_10822_));
 sky130_fd_sc_hd__nand2_1 _14808_ (.A(_10811_),
    .B(_10822_),
    .Y(_10833_));
 sky130_fd_sc_hd__inv_2 _14809_ (.A(_10833_),
    .Y(_10843_));
 sky130_fd_sc_hd__nand2_2 _14810_ (.A(_10789_),
    .B(_10843_),
    .Y(_10854_));
 sky130_fd_sc_hd__nand3_2 _14811_ (.A(_10767_),
    .B(_10833_),
    .C(_10778_),
    .Y(_10865_));
 sky130_fd_sc_hd__nand2_2 _14812_ (.A(_10854_),
    .B(_10865_),
    .Y(_10876_));
 sky130_fd_sc_hd__buf_6 _14813_ (.A(_10679_),
    .X(_10887_));
 sky130_fd_sc_hd__nand2_1 _14814_ (.A(_10876_),
    .B(_10887_),
    .Y(_10898_));
 sky130_fd_sc_hd__buf_6 _14815_ (.A(_10668_),
    .X(_10909_));
 sky130_fd_sc_hd__nand3_1 _14816_ (.A(_10854_),
    .B(_10909_),
    .C(_10865_),
    .Y(_10920_));
 sky130_fd_sc_hd__nand2_1 _14817_ (.A(_10898_),
    .B(_10920_),
    .Y(_10931_));
 sky130_fd_sc_hd__nand2_1 _14818_ (.A(_10745_),
    .B(_10931_),
    .Y(_10942_));
 sky130_fd_sc_hd__nor2_2 _14819_ (.A(_10547_),
    .B(_10942_),
    .Y(_10953_));
 sky130_fd_sc_hd__nand2_2 _14820_ (.A(_10953_),
    .B(_10086_),
    .Y(_10964_));
 sky130_fd_sc_hd__nand2_1 _14821_ (.A(_10876_),
    .B(_10909_),
    .Y(_10975_));
 sky130_fd_sc_hd__nand3_1 _14822_ (.A(_10854_),
    .B(_10679_),
    .C(_10865_),
    .Y(_10986_));
 sky130_fd_sc_hd__nand2_1 _14823_ (.A(_10975_),
    .B(_10986_),
    .Y(_10997_));
 sky130_fd_sc_hd__nor2_2 _14824_ (.A(_10997_),
    .B(_10734_),
    .Y(_11008_));
 sky130_fd_sc_hd__o21ai_1 _14825_ (.A1(_10514_),
    .A2(_10536_),
    .B1(_10503_),
    .Y(_11019_));
 sky130_fd_sc_hd__a21oi_1 _14826_ (.A1(_10854_),
    .A2(_10865_),
    .B1(_10887_),
    .Y(_11030_));
 sky130_fd_sc_hd__o21ai_1 _14827_ (.A1(_10723_),
    .A2(_11030_),
    .B1(_10986_),
    .Y(_11041_));
 sky130_fd_sc_hd__a21oi_2 _14828_ (.A1(_11008_),
    .A2(_11019_),
    .B1(_11041_),
    .Y(_11052_));
 sky130_fd_sc_hd__nand2_4 _14829_ (.A(_11052_),
    .B(_10964_),
    .Y(_11063_));
 sky130_fd_sc_hd__inv_2 _14830_ (.A(_11063_),
    .Y(_11074_));
 sky130_fd_sc_hd__inv_2 _14831_ (.A(_08867_),
    .Y(_11085_));
 sky130_fd_sc_hd__or2_1 _14832_ (.A(_11085_),
    .B(_08197_),
    .X(_11096_));
 sky130_fd_sc_hd__nand2_1 _14833_ (.A(_08197_),
    .B(_11085_),
    .Y(_11107_));
 sky130_fd_sc_hd__nand2_1 _14834_ (.A(_11096_),
    .B(_11107_),
    .Y(_11118_));
 sky130_fd_sc_hd__nand2_1 _14835_ (.A(_11118_),
    .B(_08746_),
    .Y(_11129_));
 sky130_fd_sc_hd__inv_2 _14836_ (.A(_08746_),
    .Y(_11140_));
 sky130_fd_sc_hd__nand3_1 _14837_ (.A(_11096_),
    .B(_11140_),
    .C(_11107_),
    .Y(_11151_));
 sky130_fd_sc_hd__nand2_2 _14838_ (.A(_11129_),
    .B(_11151_),
    .Y(_11162_));
 sky130_fd_sc_hd__inv_2 _14839_ (.A(_07879_),
    .Y(_11173_));
 sky130_fd_sc_hd__nand2_1 _14840_ (.A(_07637_),
    .B(_11173_),
    .Y(_11184_));
 sky130_fd_sc_hd__inv_2 _14841_ (.A(_08164_),
    .Y(_11195_));
 sky130_fd_sc_hd__nand2_1 _14842_ (.A(_11184_),
    .B(_11195_),
    .Y(_11206_));
 sky130_fd_sc_hd__clkinvlp_2 _14843_ (.A(_08099_),
    .Y(_11217_));
 sky130_fd_sc_hd__nand2_1 _14844_ (.A(_11206_),
    .B(_11217_),
    .Y(_11228_));
 sky130_fd_sc_hd__nand2_1 _14845_ (.A(_11228_),
    .B(_08088_),
    .Y(_11239_));
 sky130_fd_sc_hd__inv_2 _14846_ (.A(_07989_),
    .Y(_11250_));
 sky130_fd_sc_hd__nand2_1 _14847_ (.A(_11239_),
    .B(_11250_),
    .Y(_11261_));
 sky130_fd_sc_hd__nand3_1 _14848_ (.A(_11228_),
    .B(_07989_),
    .C(_08088_),
    .Y(_11272_));
 sky130_fd_sc_hd__nand2_1 _14849_ (.A(_11261_),
    .B(_11272_),
    .Y(_11283_));
 sky130_fd_sc_hd__inv_2 _14850_ (.A(_11283_),
    .Y(_11294_));
 sky130_fd_sc_hd__nand2_1 _14851_ (.A(_11294_),
    .B(_08834_),
    .Y(_11305_));
 sky130_fd_sc_hd__o21ai_1 _14852_ (.A1(_11162_),
    .A2(_11305_),
    .B1(_11151_),
    .Y(_11316_));
 sky130_fd_sc_hd__nand2_1 _14853_ (.A(_11107_),
    .B(_08856_),
    .Y(_11327_));
 sky130_fd_sc_hd__inv_2 _14854_ (.A(_08779_),
    .Y(_11338_));
 sky130_fd_sc_hd__nand2_1 _14855_ (.A(_11327_),
    .B(_11338_),
    .Y(_11349_));
 sky130_fd_sc_hd__nand3_1 _14856_ (.A(_11107_),
    .B(_08779_),
    .C(_08856_),
    .Y(_11360_));
 sky130_fd_sc_hd__nand2_1 _14857_ (.A(_11349_),
    .B(_11360_),
    .Y(_11371_));
 sky130_fd_sc_hd__nand2_1 _14858_ (.A(_11371_),
    .B(_09054_),
    .Y(_11382_));
 sky130_fd_sc_hd__nand3_1 _14859_ (.A(_11349_),
    .B(_09076_),
    .C(_11360_),
    .Y(_11393_));
 sky130_fd_sc_hd__nand2_1 _14860_ (.A(_11382_),
    .B(_11393_),
    .Y(_11403_));
 sky130_fd_sc_hd__nand2_1 _14861_ (.A(_08197_),
    .B(_08878_),
    .Y(_11414_));
 sky130_fd_sc_hd__inv_2 _14862_ (.A(_09164_),
    .Y(_11425_));
 sky130_fd_sc_hd__nand2_1 _14863_ (.A(_11414_),
    .B(_11425_),
    .Y(_11436_));
 sky130_fd_sc_hd__inv_2 _14864_ (.A(_09098_),
    .Y(_11447_));
 sky130_fd_sc_hd__nand2_1 _14865_ (.A(_11436_),
    .B(_11447_),
    .Y(_11458_));
 sky130_fd_sc_hd__nand3_1 _14866_ (.A(_11414_),
    .B(_09098_),
    .C(_11425_),
    .Y(_11469_));
 sky130_fd_sc_hd__nand2_1 _14867_ (.A(_11458_),
    .B(_11469_),
    .Y(_11480_));
 sky130_fd_sc_hd__nand2_1 _14868_ (.A(_11480_),
    .B(_08944_),
    .Y(_11491_));
 sky130_fd_sc_hd__nand3_1 _14869_ (.A(_11458_),
    .B(_11469_),
    .C(_08966_),
    .Y(_11502_));
 sky130_fd_sc_hd__nand2_2 _14870_ (.A(_11491_),
    .B(_11502_),
    .Y(_11513_));
 sky130_fd_sc_hd__nor2_1 _14871_ (.A(_11403_),
    .B(_11513_),
    .Y(_11524_));
 sky130_fd_sc_hd__o21ai_1 _14872_ (.A1(_11393_),
    .A2(_11513_),
    .B1(_11502_),
    .Y(_11535_));
 sky130_fd_sc_hd__a21oi_1 _14873_ (.A1(_11316_),
    .A2(_11524_),
    .B1(_11535_),
    .Y(_11546_));
 sky130_fd_sc_hd__nand3_1 _14874_ (.A(_11184_),
    .B(_08099_),
    .C(_11195_),
    .Y(_11557_));
 sky130_fd_sc_hd__nand2_1 _14875_ (.A(_11228_),
    .B(_11557_),
    .Y(_11568_));
 sky130_fd_sc_hd__buf_6 _14876_ (.A(_07967_),
    .X(_11579_));
 sky130_fd_sc_hd__nand2_1 _14877_ (.A(_11568_),
    .B(_11579_),
    .Y(_11590_));
 sky130_fd_sc_hd__nand3_1 _14878_ (.A(_11228_),
    .B(_07912_),
    .C(_11557_),
    .Y(_11601_));
 sky130_fd_sc_hd__nand2_1 _14879_ (.A(_11590_),
    .B(_11601_),
    .Y(_11612_));
 sky130_fd_sc_hd__nand2_1 _14880_ (.A(_07637_),
    .B(_07758_),
    .Y(_11623_));
 sky130_fd_sc_hd__nand2_1 _14881_ (.A(_11623_),
    .B(_07736_),
    .Y(_11634_));
 sky130_fd_sc_hd__nand2_1 _14882_ (.A(_11634_),
    .B(_07868_),
    .Y(_11645_));
 sky130_fd_sc_hd__nand3_1 _14883_ (.A(_11623_),
    .B(_07857_),
    .C(_07736_),
    .Y(_11656_));
 sky130_fd_sc_hd__nand2_2 _14884_ (.A(_11645_),
    .B(_11656_),
    .Y(_11667_));
 sky130_fd_sc_hd__inv_2 _14885_ (.A(_11667_),
    .Y(_11678_));
 sky130_fd_sc_hd__nand2_1 _14886_ (.A(_11678_),
    .B(_08055_),
    .Y(_11689_));
 sky130_fd_sc_hd__nand2_1 _14887_ (.A(_11667_),
    .B(_08066_),
    .Y(_11700_));
 sky130_fd_sc_hd__nand2_1 _14888_ (.A(_11689_),
    .B(_11700_),
    .Y(_11711_));
 sky130_fd_sc_hd__nor2_1 _14889_ (.A(_11612_),
    .B(_11711_),
    .Y(_11722_));
 sky130_fd_sc_hd__inv_2 _14890_ (.A(_07582_),
    .Y(_11733_));
 sky130_fd_sc_hd__or2_1 _14891_ (.A(_11733_),
    .B(_07352_),
    .X(_11744_));
 sky130_fd_sc_hd__nand2_1 _14892_ (.A(_07352_),
    .B(_11733_),
    .Y(_11755_));
 sky130_fd_sc_hd__nand2_1 _14893_ (.A(_11744_),
    .B(_11755_),
    .Y(_11766_));
 sky130_fd_sc_hd__buf_6 _14894_ (.A(_07429_),
    .X(_11777_));
 sky130_fd_sc_hd__nand2b_1 _14895_ (.A_N(_11766_),
    .B(_11777_),
    .Y(_11788_));
 sky130_fd_sc_hd__buf_8 _14896_ (.A(_07418_),
    .X(_11799_));
 sky130_fd_sc_hd__nand2_1 _14897_ (.A(_11766_),
    .B(_11799_),
    .Y(_11810_));
 sky130_fd_sc_hd__and2_1 _14898_ (.A(_11788_),
    .B(_11810_),
    .X(_11821_));
 sky130_fd_sc_hd__a21o_1 _14899_ (.A1(_08790_),
    .A2(net1),
    .B1(_07308_),
    .X(_11832_));
 sky130_fd_sc_hd__nand2_1 _14900_ (.A(_11832_),
    .B(_07319_),
    .Y(_11843_));
 sky130_fd_sc_hd__inv_2 _14901_ (.A(_11843_),
    .Y(_11854_));
 sky130_fd_sc_hd__nand2_1 _14902_ (.A(_11854_),
    .B(_07242_),
    .Y(_11865_));
 sky130_fd_sc_hd__clkinvlp_2 _14903_ (.A(_11865_),
    .Y(_11876_));
 sky130_fd_sc_hd__a21o_1 _14904_ (.A1(_07253_),
    .A2(_07286_),
    .B1(_07330_),
    .X(_11887_));
 sky130_fd_sc_hd__nand2_1 _14905_ (.A(_11887_),
    .B(_07341_),
    .Y(_11898_));
 sky130_fd_sc_hd__nor2_1 _14906_ (.A(_07560_),
    .B(_11898_),
    .Y(_11909_));
 sky130_fd_sc_hd__inv_2 _14907_ (.A(_11909_),
    .Y(_11920_));
 sky130_fd_sc_hd__nand2_1 _14908_ (.A(_11898_),
    .B(_07560_),
    .Y(_11931_));
 sky130_fd_sc_hd__nand2_1 _14909_ (.A(_11920_),
    .B(_11931_),
    .Y(_11942_));
 sky130_fd_sc_hd__inv_2 _14910_ (.A(_11942_),
    .Y(_11953_));
 sky130_fd_sc_hd__nand3_1 _14911_ (.A(_11821_),
    .B(_11876_),
    .C(_11953_),
    .Y(_11964_));
 sky130_fd_sc_hd__a21boi_1 _14912_ (.A1(_11810_),
    .A2(_11909_),
    .B1_N(_11788_),
    .Y(_11974_));
 sky130_fd_sc_hd__nand2_1 _14913_ (.A(_11964_),
    .B(_11974_),
    .Y(_11985_));
 sky130_fd_sc_hd__or2_1 _14914_ (.A(_07758_),
    .B(_07637_),
    .X(_11996_));
 sky130_fd_sc_hd__nand2_2 _14915_ (.A(_11996_),
    .B(_11623_),
    .Y(_12007_));
 sky130_fd_sc_hd__inv_2 _14916_ (.A(_12007_),
    .Y(_12018_));
 sky130_fd_sc_hd__buf_6 _14917_ (.A(_07824_),
    .X(_12029_));
 sky130_fd_sc_hd__nand2_1 _14918_ (.A(_12018_),
    .B(_12029_),
    .Y(_12040_));
 sky130_fd_sc_hd__buf_6 _14919_ (.A(_07813_),
    .X(_12051_));
 sky130_fd_sc_hd__nand2_1 _14920_ (.A(_12007_),
    .B(_12051_),
    .Y(_12062_));
 sky130_fd_sc_hd__nand2_1 _14921_ (.A(_12040_),
    .B(_12062_),
    .Y(_12073_));
 sky130_fd_sc_hd__inv_2 _14922_ (.A(_07484_),
    .Y(_12084_));
 sky130_fd_sc_hd__nand2_1 _14923_ (.A(_11755_),
    .B(_07549_),
    .Y(_12095_));
 sky130_fd_sc_hd__or2_1 _14924_ (.A(_12084_),
    .B(_12095_),
    .X(_12106_));
 sky130_fd_sc_hd__nand2_1 _14925_ (.A(_12095_),
    .B(_12084_),
    .Y(_12117_));
 sky130_fd_sc_hd__nand2_1 _14926_ (.A(_12106_),
    .B(_12117_),
    .Y(_12128_));
 sky130_fd_sc_hd__inv_2 _14927_ (.A(_12128_),
    .Y(_12139_));
 sky130_fd_sc_hd__nand2_1 _14928_ (.A(_12139_),
    .B(_07725_),
    .Y(_12150_));
 sky130_fd_sc_hd__nand2_1 _14929_ (.A(_12128_),
    .B(_07703_),
    .Y(_12161_));
 sky130_fd_sc_hd__nand2_1 _14930_ (.A(_12150_),
    .B(_12161_),
    .Y(_12172_));
 sky130_fd_sc_hd__nor2_1 _14931_ (.A(_12073_),
    .B(_12172_),
    .Y(_12183_));
 sky130_fd_sc_hd__nand3_1 _14932_ (.A(_11722_),
    .B(_11985_),
    .C(_12183_),
    .Y(_12194_));
 sky130_fd_sc_hd__o21ai_1 _14933_ (.A1(_12150_),
    .A2(_12073_),
    .B1(_12040_),
    .Y(_12205_));
 sky130_fd_sc_hd__nand2_1 _14934_ (.A(_12205_),
    .B(_11722_),
    .Y(_12216_));
 sky130_fd_sc_hd__o21a_1 _14935_ (.A1(_11689_),
    .A2(_11612_),
    .B1(_11601_),
    .X(_12227_));
 sky130_fd_sc_hd__nand3_2 _14936_ (.A(_12194_),
    .B(_12216_),
    .C(_12227_),
    .Y(_12238_));
 sky130_fd_sc_hd__inv_2 _14937_ (.A(_11162_),
    .Y(_12249_));
 sky130_fd_sc_hd__inv_2 _14938_ (.A(_08834_),
    .Y(_12260_));
 sky130_fd_sc_hd__nand2_1 _14939_ (.A(_11283_),
    .B(_12260_),
    .Y(_12271_));
 sky130_fd_sc_hd__nand3_1 _14940_ (.A(_12249_),
    .B(_11305_),
    .C(_12271_),
    .Y(_12282_));
 sky130_fd_sc_hd__inv_2 _14941_ (.A(_11513_),
    .Y(_12293_));
 sky130_fd_sc_hd__inv_2 _14942_ (.A(_11403_),
    .Y(_12304_));
 sky130_fd_sc_hd__nand2_1 _14943_ (.A(_12293_),
    .B(_12304_),
    .Y(_12315_));
 sky130_fd_sc_hd__nor2_1 _14944_ (.A(_12282_),
    .B(_12315_),
    .Y(_12326_));
 sky130_fd_sc_hd__nand2_1 _14945_ (.A(_12238_),
    .B(_12326_),
    .Y(_12337_));
 sky130_fd_sc_hd__nand2_2 _14946_ (.A(_11546_),
    .B(_12337_),
    .Y(_12348_));
 sky130_fd_sc_hd__nand2_1 _14947_ (.A(_11458_),
    .B(_09087_),
    .Y(_12359_));
 sky130_fd_sc_hd__nand3_1 _14948_ (.A(_12359_),
    .B(_08977_),
    .C(_08955_),
    .Y(_12370_));
 sky130_fd_sc_hd__nand3_1 _14949_ (.A(_11458_),
    .B(_08988_),
    .C(_09087_),
    .Y(_12381_));
 sky130_fd_sc_hd__nand2_1 _14950_ (.A(_12370_),
    .B(_12381_),
    .Y(_12392_));
 sky130_fd_sc_hd__nand2_1 _14951_ (.A(_12392_),
    .B(_08274_),
    .Y(_12403_));
 sky130_fd_sc_hd__inv_2 _14952_ (.A(_08318_),
    .Y(_12414_));
 sky130_fd_sc_hd__nand2_1 _14953_ (.A(_09449_),
    .B(_12414_),
    .Y(_12425_));
 sky130_fd_sc_hd__nand3_1 _14954_ (.A(_09427_),
    .B(_08318_),
    .C(_09438_),
    .Y(_12436_));
 sky130_fd_sc_hd__nand2_1 _14955_ (.A(_12425_),
    .B(_12436_),
    .Y(_12447_));
 sky130_fd_sc_hd__nand2_1 _14956_ (.A(_12447_),
    .B(_08406_),
    .Y(_12458_));
 sky130_fd_sc_hd__nand3_1 _14957_ (.A(_12425_),
    .B(_08384_),
    .C(_12436_),
    .Y(_12469_));
 sky130_fd_sc_hd__nand2_1 _14958_ (.A(_12458_),
    .B(_12469_),
    .Y(_12480_));
 sky130_fd_sc_hd__inv_2 _14959_ (.A(_12480_),
    .Y(_12491_));
 sky130_fd_sc_hd__nand3_2 _14960_ (.A(_12370_),
    .B(_08296_),
    .C(_12381_),
    .Y(_12502_));
 sky130_fd_sc_hd__nand3_1 _14961_ (.A(_12403_),
    .B(_12491_),
    .C(_12502_),
    .Y(_12513_));
 sky130_fd_sc_hd__nand3_1 _14962_ (.A(_09460_),
    .B(_08549_),
    .C(_09471_),
    .Y(_12524_));
 sky130_fd_sc_hd__nand2_1 _14963_ (.A(_09504_),
    .B(_12524_),
    .Y(_12535_));
 sky130_fd_sc_hd__nand2_1 _14964_ (.A(_12535_),
    .B(_08582_),
    .Y(_12546_));
 sky130_fd_sc_hd__nand3_1 _14965_ (.A(_09504_),
    .B(_08571_),
    .C(_12524_),
    .Y(_12556_));
 sky130_fd_sc_hd__nand2_1 _14966_ (.A(_12546_),
    .B(_12556_),
    .Y(_12567_));
 sky130_fd_sc_hd__inv_2 _14967_ (.A(_12567_),
    .Y(_12578_));
 sky130_fd_sc_hd__nand2_1 _14968_ (.A(_12425_),
    .B(_08307_),
    .Y(_12589_));
 sky130_fd_sc_hd__inv_2 _14969_ (.A(_08428_),
    .Y(_12600_));
 sky130_fd_sc_hd__nand2_1 _14970_ (.A(_12589_),
    .B(_12600_),
    .Y(_12611_));
 sky130_fd_sc_hd__nand3_1 _14971_ (.A(_12425_),
    .B(_08428_),
    .C(_08307_),
    .Y(_12622_));
 sky130_fd_sc_hd__nand2_1 _14972_ (.A(_12611_),
    .B(_12622_),
    .Y(_12633_));
 sky130_fd_sc_hd__nand2_1 _14973_ (.A(_12633_),
    .B(_08527_),
    .Y(_12644_));
 sky130_fd_sc_hd__nand3_2 _14974_ (.A(_12611_),
    .B(_08505_),
    .C(_12622_),
    .Y(_12655_));
 sky130_fd_sc_hd__nand2_1 _14975_ (.A(_12644_),
    .B(_12655_),
    .Y(_12666_));
 sky130_fd_sc_hd__inv_2 _14976_ (.A(_12666_),
    .Y(_12677_));
 sky130_fd_sc_hd__nand2_1 _14977_ (.A(_12578_),
    .B(_12677_),
    .Y(_12688_));
 sky130_fd_sc_hd__nor2_1 _14978_ (.A(_12513_),
    .B(_12688_),
    .Y(_12699_));
 sky130_fd_sc_hd__nand2_1 _14979_ (.A(_12348_),
    .B(_12699_),
    .Y(_12710_));
 sky130_fd_sc_hd__o21ai_1 _14980_ (.A1(_12480_),
    .A2(_12502_),
    .B1(_12469_),
    .Y(_12721_));
 sky130_fd_sc_hd__nor2_1 _14981_ (.A(_12567_),
    .B(_12666_),
    .Y(_12732_));
 sky130_fd_sc_hd__nand2_1 _14982_ (.A(_12721_),
    .B(_12732_),
    .Y(_12743_));
 sky130_fd_sc_hd__inv_2 _14983_ (.A(_12655_),
    .Y(_12754_));
 sky130_fd_sc_hd__a21boi_1 _14984_ (.A1(_12754_),
    .A2(_12546_),
    .B1_N(_12556_),
    .Y(_12765_));
 sky130_fd_sc_hd__nand2_1 _14985_ (.A(_12743_),
    .B(_12765_),
    .Y(_12776_));
 sky130_fd_sc_hd__inv_2 _14986_ (.A(_12776_),
    .Y(_12787_));
 sky130_fd_sc_hd__nand2_2 _14987_ (.A(_12710_),
    .B(_12787_),
    .Y(_12798_));
 sky130_fd_sc_hd__inv_2 _14988_ (.A(_09767_),
    .Y(_12809_));
 sky130_fd_sc_hd__nand2_1 _14989_ (.A(_09921_),
    .B(_10009_),
    .Y(_12820_));
 sky130_fd_sc_hd__nand3_1 _14990_ (.A(_09899_),
    .B(_09987_),
    .C(_09910_),
    .Y(_12831_));
 sky130_fd_sc_hd__nand2_1 _14991_ (.A(_12820_),
    .B(_12831_),
    .Y(_12842_));
 sky130_fd_sc_hd__nand2_1 _14992_ (.A(_12809_),
    .B(_12842_),
    .Y(_12853_));
 sky130_fd_sc_hd__nand2_1 _14993_ (.A(_09537_),
    .B(_09570_),
    .Y(_12864_));
 sky130_fd_sc_hd__nand2_1 _14994_ (.A(_12864_),
    .B(_09548_),
    .Y(_12875_));
 sky130_fd_sc_hd__inv_2 _14995_ (.A(_09405_),
    .Y(_12886_));
 sky130_fd_sc_hd__nand3_1 _14996_ (.A(_12875_),
    .B(_12886_),
    .C(_09581_),
    .Y(_12897_));
 sky130_fd_sc_hd__nor2_2 _14997_ (.A(_12853_),
    .B(_12897_),
    .Y(_12908_));
 sky130_fd_sc_hd__nand3_2 _14998_ (.A(_12798_),
    .B(_10953_),
    .C(_12908_),
    .Y(_12919_));
 sky130_fd_sc_hd__o21ai_4 _14999_ (.A1(net15),
    .A2(_08790_),
    .B1(_10909_),
    .Y(_12930_));
 sky130_fd_sc_hd__nand2_2 _15000_ (.A(_10854_),
    .B(_10822_),
    .Y(_12941_));
 sky130_fd_sc_hd__xor2_4 _15001_ (.A(_12930_),
    .B(_12941_),
    .X(_12952_));
 sky130_fd_sc_hd__nand3_2 _15002_ (.A(_11074_),
    .B(_12919_),
    .C(_12952_),
    .Y(_12963_));
 sky130_fd_sc_hd__buf_6 _15003_ (.A(_12963_),
    .X(_12974_));
 sky130_fd_sc_hd__buf_8 _15004_ (.A(_12974_),
    .X(\div1i.quot[23] ));
 sky130_fd_sc_hd__nand2_1 _15005_ (.A(_11843_),
    .B(_07231_),
    .Y(_12995_));
 sky130_fd_sc_hd__nand2_1 _15006_ (.A(_11865_),
    .B(_12995_),
    .Y(_13006_));
 sky130_fd_sc_hd__nand2_1 _15007_ (.A(_12974_),
    .B(_13006_),
    .Y(_13017_));
 sky130_fd_sc_hd__inv_2 _15008_ (.A(_10547_),
    .Y(_13028_));
 sky130_fd_sc_hd__nand3_2 _15009_ (.A(_12908_),
    .B(_11008_),
    .C(_13028_),
    .Y(_13039_));
 sky130_fd_sc_hd__a21oi_1 _15010_ (.A1(_12348_),
    .A2(_12699_),
    .B1(_12776_),
    .Y(_13050_));
 sky130_fd_sc_hd__nor2_4 _15011_ (.A(_13039_),
    .B(_13050_),
    .Y(_13061_));
 sky130_fd_sc_hd__nor2_8 _15012_ (.A(_11063_),
    .B(_13061_),
    .Y(_13072_));
 sky130_fd_sc_hd__nand3_1 _15013_ (.A(_13072_),
    .B(_11843_),
    .C(_12952_),
    .Y(_13083_));
 sky130_fd_sc_hd__nand3_1 _15014_ (.A(_13017_),
    .B(_13083_),
    .C(_07539_),
    .Y(_13094_));
 sky130_fd_sc_hd__buf_8 _15015_ (.A(_12974_),
    .X(_13104_));
 sky130_fd_sc_hd__inv_2 _15016_ (.A(_13006_),
    .Y(_13115_));
 sky130_fd_sc_hd__nand2_1 _15017_ (.A(net230),
    .B(_13115_),
    .Y(_13126_));
 sky130_fd_sc_hd__buf_6 _15018_ (.A(_13072_),
    .X(_13137_));
 sky130_fd_sc_hd__clkbuf_4 _15019_ (.A(_12952_),
    .X(_13148_));
 sky130_fd_sc_hd__nand3_1 _15020_ (.A(_13137_),
    .B(_11854_),
    .C(_13148_),
    .Y(_13159_));
 sky130_fd_sc_hd__nand3_1 _15021_ (.A(_13126_),
    .B(_13159_),
    .C(_07560_),
    .Y(_13170_));
 sky130_fd_sc_hd__nand2_2 _15022_ (.A(_13094_),
    .B(_13170_),
    .Y(_13181_));
 sky130_fd_sc_hd__inv_2 _15023_ (.A(_13181_),
    .Y(_13192_));
 sky130_fd_sc_hd__nand2_1 _15024_ (.A(net133),
    .B(_07308_),
    .Y(_13203_));
 sky130_fd_sc_hd__inv_2 _15025_ (.A(_13203_),
    .Y(_13214_));
 sky130_fd_sc_hd__nand2_2 _15026_ (.A(_13214_),
    .B(_07242_),
    .Y(_13225_));
 sky130_fd_sc_hd__inv_4 _15027_ (.A(_13225_),
    .Y(_13236_));
 sky130_fd_sc_hd__xor2_1 _15028_ (.A(_11876_),
    .B(_11942_),
    .X(_13247_));
 sky130_fd_sc_hd__nand2_1 _15029_ (.A(_13104_),
    .B(_13247_),
    .Y(_13258_));
 sky130_fd_sc_hd__nand3_1 _15030_ (.A(_13137_),
    .B(_11898_),
    .C(_13148_),
    .Y(_13269_));
 sky130_fd_sc_hd__nand2_2 _15031_ (.A(_13258_),
    .B(_13269_),
    .Y(_13280_));
 sky130_fd_sc_hd__nand2_1 _15032_ (.A(_13280_),
    .B(_11777_),
    .Y(_13291_));
 sky130_fd_sc_hd__nand3_1 _15033_ (.A(_13258_),
    .B(_13269_),
    .C(_11799_),
    .Y(_13302_));
 sky130_fd_sc_hd__nand2_1 _15034_ (.A(_13291_),
    .B(_13302_),
    .Y(_13313_));
 sky130_fd_sc_hd__nand3_1 _15035_ (.A(_13192_),
    .B(_13236_),
    .C(_13313_),
    .Y(_13324_));
 sky130_fd_sc_hd__clkinvlp_2 _15036_ (.A(_13094_),
    .Y(_13335_));
 sky130_fd_sc_hd__nand2_1 _15037_ (.A(_13280_),
    .B(_11799_),
    .Y(_13346_));
 sky130_fd_sc_hd__nor2_1 _15038_ (.A(_11799_),
    .B(_13280_),
    .Y(_13357_));
 sky130_fd_sc_hd__a21oi_2 _15039_ (.A1(_13335_),
    .A2(_13346_),
    .B1(_13357_),
    .Y(_13368_));
 sky130_fd_sc_hd__nand2_2 _15040_ (.A(_13324_),
    .B(_13368_),
    .Y(_13379_));
 sky130_fd_sc_hd__a21bo_1 _15041_ (.A1(_11985_),
    .A2(_12161_),
    .B1_N(_12150_),
    .X(_13390_));
 sky130_fd_sc_hd__xor2_1 _15042_ (.A(_12073_),
    .B(_13390_),
    .X(_13401_));
 sky130_fd_sc_hd__nand2_2 _15043_ (.A(net133),
    .B(_13401_),
    .Y(_13412_));
 sky130_fd_sc_hd__nand3_1 _15044_ (.A(_13072_),
    .B(_12007_),
    .C(_12952_),
    .Y(_13423_));
 sky130_fd_sc_hd__nand3_4 _15045_ (.A(_13412_),
    .B(_13423_),
    .C(_08055_),
    .Y(_13434_));
 sky130_fd_sc_hd__clkinvlp_2 _15046_ (.A(_13401_),
    .Y(_13445_));
 sky130_fd_sc_hd__nand2_1 _15047_ (.A(net133),
    .B(_13445_),
    .Y(_13456_));
 sky130_fd_sc_hd__nand3_1 _15048_ (.A(_13072_),
    .B(_12018_),
    .C(_12952_),
    .Y(_13467_));
 sky130_fd_sc_hd__nand3_1 _15049_ (.A(_13456_),
    .B(_13467_),
    .C(_08066_),
    .Y(_13478_));
 sky130_fd_sc_hd__nand2_2 _15050_ (.A(_13434_),
    .B(_13478_),
    .Y(_13489_));
 sky130_fd_sc_hd__clkinvlp_2 _15051_ (.A(_13489_),
    .Y(_13500_));
 sky130_fd_sc_hd__a21o_1 _15052_ (.A1(_11985_),
    .A2(_12183_),
    .B1(_12205_),
    .X(_13511_));
 sky130_fd_sc_hd__xor2_1 _15053_ (.A(_11711_),
    .B(_13511_),
    .X(_13522_));
 sky130_fd_sc_hd__inv_2 _15054_ (.A(_13522_),
    .Y(_13533_));
 sky130_fd_sc_hd__nand2_2 _15055_ (.A(net230),
    .B(_13533_),
    .Y(_13544_));
 sky130_fd_sc_hd__nand3_1 _15056_ (.A(_13137_),
    .B(_11678_),
    .C(_13148_),
    .Y(_13555_));
 sky130_fd_sc_hd__nand2_2 _15057_ (.A(_13544_),
    .B(_13555_),
    .Y(_13566_));
 sky130_fd_sc_hd__nand2_1 _15058_ (.A(_13566_),
    .B(_11579_),
    .Y(_13577_));
 sky130_fd_sc_hd__buf_6 _15059_ (.A(_07912_),
    .X(_13588_));
 sky130_fd_sc_hd__nand3_1 _15060_ (.A(_13544_),
    .B(_13555_),
    .C(_13588_),
    .Y(_13599_));
 sky130_fd_sc_hd__nand2_1 _15061_ (.A(_13577_),
    .B(_13599_),
    .Y(_13610_));
 sky130_fd_sc_hd__nand2_1 _15062_ (.A(_13500_),
    .B(_13610_),
    .Y(_13621_));
 sky130_fd_sc_hd__a21oi_1 _15063_ (.A1(_11931_),
    .A2(_11876_),
    .B1(_11909_),
    .Y(_13632_));
 sky130_fd_sc_hd__xor2_1 _15064_ (.A(_13632_),
    .B(_11821_),
    .X(_13643_));
 sky130_fd_sc_hd__nand2_1 _15065_ (.A(net133),
    .B(_13643_),
    .Y(_13654_));
 sky130_fd_sc_hd__nand3_1 _15066_ (.A(_13072_),
    .B(_11766_),
    .C(_12952_),
    .Y(_13665_));
 sky130_fd_sc_hd__nand2_2 _15067_ (.A(_13654_),
    .B(_13665_),
    .Y(_13675_));
 sky130_fd_sc_hd__nand2_1 _15068_ (.A(_13675_),
    .B(_07703_),
    .Y(_13686_));
 sky130_fd_sc_hd__nand3_1 _15069_ (.A(_13654_),
    .B(_13665_),
    .C(_07725_),
    .Y(_13697_));
 sky130_fd_sc_hd__nand2_1 _15070_ (.A(_13686_),
    .B(_13697_),
    .Y(_13708_));
 sky130_fd_sc_hd__inv_2 _15071_ (.A(_13708_),
    .Y(_13719_));
 sky130_fd_sc_hd__xor2_1 _15072_ (.A(_12172_),
    .B(_11985_),
    .X(_13730_));
 sky130_fd_sc_hd__inv_2 _15073_ (.A(_13730_),
    .Y(_13741_));
 sky130_fd_sc_hd__nand2_1 _15074_ (.A(_13104_),
    .B(_13741_),
    .Y(_13752_));
 sky130_fd_sc_hd__nand3_1 _15075_ (.A(_13137_),
    .B(_12139_),
    .C(_13148_),
    .Y(_13763_));
 sky130_fd_sc_hd__nand2_1 _15076_ (.A(_13752_),
    .B(_13763_),
    .Y(_13774_));
 sky130_fd_sc_hd__nand2_1 _15077_ (.A(_13774_),
    .B(_12051_),
    .Y(_13785_));
 sky130_fd_sc_hd__nand3_1 _15078_ (.A(_13752_),
    .B(_13763_),
    .C(_12029_),
    .Y(_13796_));
 sky130_fd_sc_hd__nand2_1 _15079_ (.A(_13785_),
    .B(_13796_),
    .Y(_13807_));
 sky130_fd_sc_hd__nand2_1 _15080_ (.A(_13719_),
    .B(_13807_),
    .Y(_13818_));
 sky130_fd_sc_hd__nor2_1 _15081_ (.A(_13621_),
    .B(_13818_),
    .Y(_13829_));
 sky130_fd_sc_hd__nand2_2 _15082_ (.A(_13829_),
    .B(_13379_),
    .Y(_13840_));
 sky130_fd_sc_hd__nor2_1 _15083_ (.A(_12029_),
    .B(_13774_),
    .Y(_13851_));
 sky130_fd_sc_hd__nand2_1 _15084_ (.A(_13774_),
    .B(_12029_),
    .Y(_13862_));
 sky130_fd_sc_hd__o21ai_1 _15085_ (.A1(_13697_),
    .A2(_13851_),
    .B1(_13862_),
    .Y(_13873_));
 sky130_fd_sc_hd__nand2_1 _15086_ (.A(\div1i.quot[23] ),
    .B(_13522_),
    .Y(_13884_));
 sky130_fd_sc_hd__nand3_1 _15087_ (.A(_13137_),
    .B(_11667_),
    .C(_13148_),
    .Y(_13895_));
 sky130_fd_sc_hd__nand3_1 _15088_ (.A(_13884_),
    .B(_13895_),
    .C(_13588_),
    .Y(_13906_));
 sky130_fd_sc_hd__nand3_1 _15089_ (.A(_13544_),
    .B(_13555_),
    .C(_11579_),
    .Y(_13917_));
 sky130_fd_sc_hd__nand2_1 _15090_ (.A(_13906_),
    .B(_13917_),
    .Y(_13928_));
 sky130_fd_sc_hd__nor2_1 _15091_ (.A(_13928_),
    .B(_13489_),
    .Y(_13939_));
 sky130_fd_sc_hd__nor2_1 _15092_ (.A(_13588_),
    .B(_13566_),
    .Y(_13950_));
 sky130_fd_sc_hd__o21ai_1 _15093_ (.A1(_13434_),
    .A2(_13950_),
    .B1(_13906_),
    .Y(_13961_));
 sky130_fd_sc_hd__a21oi_2 _15094_ (.A1(_13873_),
    .A2(_13939_),
    .B1(_13961_),
    .Y(_13972_));
 sky130_fd_sc_hd__nand2_4 _15095_ (.A(_13840_),
    .B(_13972_),
    .Y(_13983_));
 sky130_fd_sc_hd__inv_2 _15096_ (.A(_12282_),
    .Y(_13994_));
 sky130_fd_sc_hd__a21o_1 _15097_ (.A1(_12238_),
    .A2(_13994_),
    .B1(_11316_),
    .X(_14005_));
 sky130_fd_sc_hd__nand2_1 _15098_ (.A(_14005_),
    .B(_12304_),
    .Y(_14016_));
 sky130_fd_sc_hd__nand2_1 _15099_ (.A(_14016_),
    .B(_11393_),
    .Y(_14027_));
 sky130_fd_sc_hd__xor2_1 _15100_ (.A(_11513_),
    .B(_14027_),
    .X(_14038_));
 sky130_fd_sc_hd__nand2_1 _15101_ (.A(net133),
    .B(_14038_),
    .Y(_14049_));
 sky130_fd_sc_hd__nand3_1 _15102_ (.A(_13072_),
    .B(_11480_),
    .C(_12952_),
    .Y(_14060_));
 sky130_fd_sc_hd__nand2_1 _15103_ (.A(_14049_),
    .B(_14060_),
    .Y(_14071_));
 sky130_fd_sc_hd__nand2_1 _15104_ (.A(_14071_),
    .B(_08274_),
    .Y(_14082_));
 sky130_fd_sc_hd__nand3_2 _15105_ (.A(_14049_),
    .B(_14060_),
    .C(_08296_),
    .Y(_14093_));
 sky130_fd_sc_hd__nand2_1 _15106_ (.A(_14082_),
    .B(_14093_),
    .Y(_14104_));
 sky130_fd_sc_hd__inv_2 _15107_ (.A(_14104_),
    .Y(_14115_));
 sky130_fd_sc_hd__a21o_1 _15108_ (.A1(_12502_),
    .A2(_12403_),
    .B1(_12348_),
    .X(_14126_));
 sky130_fd_sc_hd__nand3_1 _15109_ (.A(_12348_),
    .B(_12502_),
    .C(_12403_),
    .Y(_14137_));
 sky130_fd_sc_hd__nand2_1 _15110_ (.A(_14126_),
    .B(_14137_),
    .Y(_14148_));
 sky130_fd_sc_hd__nand2_1 _15111_ (.A(_12963_),
    .B(_14148_),
    .Y(_14159_));
 sky130_fd_sc_hd__nand3_1 _15112_ (.A(_13072_),
    .B(_12392_),
    .C(_12952_),
    .Y(_14170_));
 sky130_fd_sc_hd__nand2_1 _15113_ (.A(_14159_),
    .B(_14170_),
    .Y(_14181_));
 sky130_fd_sc_hd__nand2_1 _15114_ (.A(_14181_),
    .B(_08406_),
    .Y(_14192_));
 sky130_fd_sc_hd__nand3_1 _15115_ (.A(_14159_),
    .B(_14170_),
    .C(_08384_),
    .Y(_14203_));
 sky130_fd_sc_hd__nand2_1 _15116_ (.A(_14192_),
    .B(_14203_),
    .Y(_14213_));
 sky130_fd_sc_hd__inv_2 _15117_ (.A(_14213_),
    .Y(_14224_));
 sky130_fd_sc_hd__nand2_1 _15118_ (.A(_14115_),
    .B(_14224_),
    .Y(_14235_));
 sky130_fd_sc_hd__inv_2 _15119_ (.A(_14235_),
    .Y(_14246_));
 sky130_fd_sc_hd__inv_2 _15120_ (.A(_12513_),
    .Y(_14257_));
 sky130_fd_sc_hd__nand2_1 _15121_ (.A(_12348_),
    .B(_14257_),
    .Y(_14268_));
 sky130_fd_sc_hd__inv_2 _15122_ (.A(_12721_),
    .Y(_14279_));
 sky130_fd_sc_hd__nand2_1 _15123_ (.A(_14268_),
    .B(_14279_),
    .Y(_14290_));
 sky130_fd_sc_hd__or2_1 _15124_ (.A(_12677_),
    .B(_14290_),
    .X(_00047_));
 sky130_fd_sc_hd__nand2_1 _15125_ (.A(_14290_),
    .B(_12677_),
    .Y(_00058_));
 sky130_fd_sc_hd__nand2_1 _15126_ (.A(_00047_),
    .B(_00058_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_1 _15127_ (.A(net230),
    .B(_00069_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand3_1 _15128_ (.A(_13137_),
    .B(_12633_),
    .C(_13148_),
    .Y(_00091_));
 sky130_fd_sc_hd__nand2_1 _15129_ (.A(_00080_),
    .B(_00091_),
    .Y(_00102_));
 sky130_fd_sc_hd__nand2_1 _15130_ (.A(_00102_),
    .B(_08582_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand3_1 _15131_ (.A(_00080_),
    .B(_00091_),
    .C(_08571_),
    .Y(_00124_));
 sky130_fd_sc_hd__nand2_2 _15132_ (.A(_00113_),
    .B(_00124_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand2_1 _15133_ (.A(_14137_),
    .B(_12502_),
    .Y(_00146_));
 sky130_fd_sc_hd__xor2_1 _15134_ (.A(_12480_),
    .B(_00146_),
    .X(_00157_));
 sky130_fd_sc_hd__nand2_2 _15135_ (.A(net230),
    .B(_00157_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand3_1 _15136_ (.A(_13137_),
    .B(_12447_),
    .C(_13148_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_2 _15137_ (.A(_00168_),
    .B(_00179_),
    .Y(_00190_));
 sky130_fd_sc_hd__nand2_1 _15138_ (.A(_00190_),
    .B(_08527_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand3_2 _15139_ (.A(_00168_),
    .B(_00179_),
    .C(_08505_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_2 _15140_ (.A(_00201_),
    .B(_00212_),
    .Y(_00223_));
 sky130_fd_sc_hd__nor2_2 _15141_ (.A(_00223_),
    .B(_00135_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _15142_ (.A(_14246_),
    .B(_00234_),
    .Y(_00245_));
 sky130_fd_sc_hd__a21bo_1 _15143_ (.A1(_13511_),
    .A2(_11700_),
    .B1_N(_11689_),
    .X(_00256_));
 sky130_fd_sc_hd__xor2_1 _15144_ (.A(_11612_),
    .B(_00256_),
    .X(_00267_));
 sky130_fd_sc_hd__nand2_1 _15145_ (.A(\div1i.quot[23] ),
    .B(_00267_),
    .Y(_00278_));
 sky130_fd_sc_hd__nand3_1 _15146_ (.A(_13137_),
    .B(_11568_),
    .C(_13148_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _15147_ (.A(_00278_),
    .B(_00289_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _15148_ (.A(_00300_),
    .B(_12260_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand3_1 _15149_ (.A(_00278_),
    .B(_00289_),
    .C(_08834_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _15150_ (.A(_00311_),
    .B(_00322_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _15151_ (.A(_11305_),
    .B(_12271_),
    .Y(_00344_));
 sky130_fd_sc_hd__xor2_1 _15152_ (.A(_00344_),
    .B(_12238_),
    .X(_00355_));
 sky130_fd_sc_hd__clkinvlp_2 _15153_ (.A(_00355_),
    .Y(_00366_));
 sky130_fd_sc_hd__nand2_1 _15154_ (.A(_12974_),
    .B(_00366_),
    .Y(_00377_));
 sky130_fd_sc_hd__nand3_1 _15155_ (.A(_13072_),
    .B(_11294_),
    .C(_12952_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _15156_ (.A(_00377_),
    .B(_00388_),
    .Y(_00399_));
 sky130_fd_sc_hd__nor2_1 _15157_ (.A(_00399_),
    .B(_11140_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _15158_ (.A(_00399_),
    .B(_11140_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2b_1 _15159_ (.A_N(_00410_),
    .B(_00421_),
    .Y(_00432_));
 sky130_fd_sc_hd__nor2_1 _15160_ (.A(_00432_),
    .B(_00333_),
    .Y(_00443_));
 sky130_fd_sc_hd__or2_1 _15161_ (.A(_12304_),
    .B(_14005_),
    .X(_00454_));
 sky130_fd_sc_hd__nand2_1 _15162_ (.A(_00454_),
    .B(_14016_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _15163_ (.A(\div1i.quot[23] ),
    .B(_00465_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand3_1 _15164_ (.A(_13137_),
    .B(_11371_),
    .C(_13148_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _15165_ (.A(_00476_),
    .B(_00487_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _15166_ (.A(_00498_),
    .B(_08944_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand3_1 _15167_ (.A(_00476_),
    .B(_00487_),
    .C(_08966_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_2 _15168_ (.A(_00508_),
    .B(_00519_),
    .Y(_00530_));
 sky130_fd_sc_hd__a21bo_1 _15169_ (.A1(_12238_),
    .A2(_12271_),
    .B1_N(_11305_),
    .X(_00541_));
 sky130_fd_sc_hd__xor2_1 _15170_ (.A(_11162_),
    .B(_00541_),
    .X(_00552_));
 sky130_fd_sc_hd__nand2_2 _15171_ (.A(net230),
    .B(_00552_),
    .Y(_00563_));
 sky130_fd_sc_hd__nand3_1 _15172_ (.A(_13137_),
    .B(_11118_),
    .C(_13148_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _15173_ (.A(_00563_),
    .B(_00574_),
    .Y(_00585_));
 sky130_fd_sc_hd__nand2_1 _15174_ (.A(_00585_),
    .B(_09054_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand3_4 _15175_ (.A(_00563_),
    .B(_00574_),
    .C(_09076_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_2 _15176_ (.A(_00596_),
    .B(_00607_),
    .Y(_00618_));
 sky130_fd_sc_hd__nor2_2 _15177_ (.A(_00530_),
    .B(_00618_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_2 _15178_ (.A(_00629_),
    .B(_00443_),
    .Y(_00640_));
 sky130_fd_sc_hd__nor2_2 _15179_ (.A(_00640_),
    .B(_00245_),
    .Y(_00651_));
 sky130_fd_sc_hd__nand2_2 _15180_ (.A(_13983_),
    .B(_00651_),
    .Y(_00662_));
 sky130_fd_sc_hd__o21ai_1 _15181_ (.A1(_00322_),
    .A2(_00410_),
    .B1(_00421_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand2_1 _15182_ (.A(_00673_),
    .B(_00629_),
    .Y(_00684_));
 sky130_fd_sc_hd__inv_2 _15183_ (.A(_00607_),
    .Y(_00695_));
 sky130_fd_sc_hd__a21boi_1 _15184_ (.A1(_00695_),
    .A2(_00508_),
    .B1_N(_00519_),
    .Y(_00706_));
 sky130_fd_sc_hd__nand2_2 _15185_ (.A(_00684_),
    .B(_00706_),
    .Y(_00717_));
 sky130_fd_sc_hd__inv_2 _15186_ (.A(_00135_),
    .Y(_00728_));
 sky130_fd_sc_hd__inv_2 _15187_ (.A(_00223_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _15188_ (.A(_00728_),
    .B(_00739_),
    .Y(_00750_));
 sky130_fd_sc_hd__nor2_2 _15189_ (.A(_00750_),
    .B(_14235_),
    .Y(_00761_));
 sky130_fd_sc_hd__inv_2 _15190_ (.A(_14093_),
    .Y(_00772_));
 sky130_fd_sc_hd__nand3_1 _15191_ (.A(_00772_),
    .B(_14192_),
    .C(_14203_),
    .Y(_00783_));
 sky130_fd_sc_hd__nand2_1 _15192_ (.A(_00783_),
    .B(_14203_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand2_1 _15193_ (.A(_00794_),
    .B(_00234_),
    .Y(_00805_));
 sky130_fd_sc_hd__and2_1 _15194_ (.A(_00102_),
    .B(_08582_),
    .X(_00816_));
 sky130_fd_sc_hd__o21a_1 _15195_ (.A1(_00212_),
    .A2(_00816_),
    .B1(_00124_),
    .X(_00827_));
 sky130_fd_sc_hd__nand2_1 _15196_ (.A(_00805_),
    .B(_00827_),
    .Y(_00838_));
 sky130_fd_sc_hd__a21oi_4 _15197_ (.A1(_00717_),
    .A2(_00761_),
    .B1(_00838_),
    .Y(_00849_));
 sky130_fd_sc_hd__nand2_4 _15198_ (.A(_00849_),
    .B(_00662_),
    .Y(_00860_));
 sky130_fd_sc_hd__inv_2 _15199_ (.A(_12535_),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_1 _15200_ (.A(_00058_),
    .B(_12655_),
    .Y(_00882_));
 sky130_fd_sc_hd__nand2_1 _15201_ (.A(_00882_),
    .B(_12578_),
    .Y(_00893_));
 sky130_fd_sc_hd__nand3_1 _15202_ (.A(_00058_),
    .B(_12567_),
    .C(_12655_),
    .Y(_00904_));
 sky130_fd_sc_hd__nand2_1 _15203_ (.A(_00893_),
    .B(_00904_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand2_1 _15204_ (.A(_00915_),
    .B(_13104_),
    .Y(_00926_));
 sky130_fd_sc_hd__o21ai_1 _15205_ (.A1(_00871_),
    .A2(\div1i.quot[23] ),
    .B1(_00926_),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2_1 _15206_ (.A(_09548_),
    .B(_00937_),
    .Y(_00948_));
 sky130_fd_sc_hd__inv_2 _15207_ (.A(_00948_),
    .Y(_00959_));
 sky130_fd_sc_hd__nand2_1 _15208_ (.A(_00937_),
    .B(_09548_),
    .Y(_00970_));
 sky130_fd_sc_hd__nand2_1 _15209_ (.A(_00959_),
    .B(_00970_),
    .Y(_00981_));
 sky130_fd_sc_hd__inv_6 _15210_ (.A(_12974_),
    .Y(_00992_));
 sky130_fd_sc_hd__nand2_1 _15211_ (.A(_00992_),
    .B(_12864_),
    .Y(_01003_));
 sky130_fd_sc_hd__nand2_1 _15212_ (.A(_12875_),
    .B(_09581_),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _15213_ (.A(_13050_),
    .B(_01014_),
    .Y(_01025_));
 sky130_fd_sc_hd__inv_2 _15214_ (.A(_01014_),
    .Y(_01036_));
 sky130_fd_sc_hd__nand2_1 _15215_ (.A(_12798_),
    .B(_01036_),
    .Y(_01046_));
 sky130_fd_sc_hd__nand2_1 _15216_ (.A(_01025_),
    .B(_01046_),
    .Y(_01057_));
 sky130_fd_sc_hd__nand2_1 _15217_ (.A(_13104_),
    .B(_01057_),
    .Y(_01068_));
 sky130_fd_sc_hd__nand2_1 _15218_ (.A(_01003_),
    .B(_01068_),
    .Y(_01079_));
 sky130_fd_sc_hd__nor2_1 _15219_ (.A(_09361_),
    .B(_01079_),
    .Y(_01090_));
 sky130_fd_sc_hd__nand2_1 _15220_ (.A(_01079_),
    .B(_09361_),
    .Y(_01101_));
 sky130_fd_sc_hd__nand2b_1 _15221_ (.A_N(_01090_),
    .B(_01101_),
    .Y(_01112_));
 sky130_fd_sc_hd__nor2_1 _15222_ (.A(_00981_),
    .B(_01112_),
    .Y(_01123_));
 sky130_fd_sc_hd__nand2_1 _15223_ (.A(_00992_),
    .B(_09680_),
    .Y(_01134_));
 sky130_fd_sc_hd__inv_2 _15224_ (.A(_12897_),
    .Y(_01145_));
 sky130_fd_sc_hd__nand2_1 _15225_ (.A(_12798_),
    .B(_01145_),
    .Y(_01156_));
 sky130_fd_sc_hd__inv_2 _15226_ (.A(_09592_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand2_1 _15227_ (.A(_01156_),
    .B(_01167_),
    .Y(_01178_));
 sky130_fd_sc_hd__nand2_1 _15228_ (.A(_01178_),
    .B(_12809_),
    .Y(_01189_));
 sky130_fd_sc_hd__nand3_1 _15229_ (.A(_01156_),
    .B(_09767_),
    .C(_01167_),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_1 _15230_ (.A(_01189_),
    .B(_01200_),
    .Y(_01211_));
 sky130_fd_sc_hd__nand2_1 _15231_ (.A(_01211_),
    .B(\div1i.quot[23] ),
    .Y(_01222_));
 sky130_fd_sc_hd__nand2_1 _15232_ (.A(_01134_),
    .B(_01222_),
    .Y(_01233_));
 sky130_fd_sc_hd__nand2_1 _15233_ (.A(_01233_),
    .B(_09987_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand3_1 _15234_ (.A(_01134_),
    .B(_01222_),
    .C(_10009_),
    .Y(_01255_));
 sky130_fd_sc_hd__nand2_1 _15235_ (.A(_01244_),
    .B(_01255_),
    .Y(_01266_));
 sky130_fd_sc_hd__nand2_1 _15236_ (.A(_01046_),
    .B(_09581_),
    .Y(_01277_));
 sky130_fd_sc_hd__xor2_1 _15237_ (.A(_09405_),
    .B(_01277_),
    .X(_01288_));
 sky130_fd_sc_hd__nand2_1 _15238_ (.A(_01288_),
    .B(\div1i.quot[23] ),
    .Y(_01299_));
 sky130_fd_sc_hd__nand2_1 _15239_ (.A(_00992_),
    .B(_09328_),
    .Y(_01310_));
 sky130_fd_sc_hd__nand2_1 _15240_ (.A(_01299_),
    .B(_01310_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_1 _15241_ (.A(_01321_),
    .B(_09735_),
    .Y(_01332_));
 sky130_fd_sc_hd__nand3_2 _15242_ (.A(_01299_),
    .B(_01310_),
    .C(_09724_),
    .Y(_01343_));
 sky130_fd_sc_hd__nand2_1 _15243_ (.A(_01332_),
    .B(_01343_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor2_2 _15244_ (.A(_01266_),
    .B(_01354_),
    .Y(_01365_));
 sky130_fd_sc_hd__nand2_1 _15245_ (.A(_01123_),
    .B(_01365_),
    .Y(_01376_));
 sky130_fd_sc_hd__nand2_1 _15246_ (.A(_12798_),
    .B(_12908_),
    .Y(_01387_));
 sky130_fd_sc_hd__inv_2 _15247_ (.A(_10086_),
    .Y(_01398_));
 sky130_fd_sc_hd__nand2_1 _15248_ (.A(_01387_),
    .B(_01398_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2_1 _15249_ (.A(_01409_),
    .B(_13028_),
    .Y(_01420_));
 sky130_fd_sc_hd__inv_2 _15250_ (.A(_11019_),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_1 _15251_ (.A(_01420_),
    .B(_01431_),
    .Y(_01442_));
 sky130_fd_sc_hd__nand2_1 _15252_ (.A(_01442_),
    .B(_10745_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand3_1 _15253_ (.A(_01420_),
    .B(_10734_),
    .C(_01431_),
    .Y(_01464_));
 sky130_fd_sc_hd__nand2_1 _15254_ (.A(_01453_),
    .B(_01464_),
    .Y(_01475_));
 sky130_fd_sc_hd__nand2_1 _15255_ (.A(_01475_),
    .B(\div1i.quot[23] ),
    .Y(_01486_));
 sky130_fd_sc_hd__nand2_1 _15256_ (.A(_00992_),
    .B(_10646_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand2_1 _15257_ (.A(_01486_),
    .B(_01497_),
    .Y(_01508_));
 sky130_fd_sc_hd__nand2_1 _15258_ (.A(_01508_),
    .B(_10909_),
    .Y(_01519_));
 sky130_fd_sc_hd__nand3_1 _15259_ (.A(_01486_),
    .B(_10887_),
    .C(_01497_),
    .Y(_01530_));
 sky130_fd_sc_hd__nand2_1 _15260_ (.A(_01519_),
    .B(_01530_),
    .Y(_01541_));
 sky130_fd_sc_hd__nand3_1 _15261_ (.A(_01409_),
    .B(_10536_),
    .C(_10262_),
    .Y(_01552_));
 sky130_fd_sc_hd__nand2_1 _15262_ (.A(_01552_),
    .B(_10536_),
    .Y(_01563_));
 sky130_fd_sc_hd__nand2_1 _15263_ (.A(_01563_),
    .B(_10525_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand3_1 _15264_ (.A(_01552_),
    .B(_10514_),
    .C(_10536_),
    .Y(_01585_));
 sky130_fd_sc_hd__nand2_1 _15265_ (.A(_01574_),
    .B(_01585_),
    .Y(_01595_));
 sky130_fd_sc_hd__nand2_1 _15266_ (.A(_01595_),
    .B(\div1i.quot[23] ),
    .Y(_01606_));
 sky130_fd_sc_hd__nand2_1 _15267_ (.A(_00992_),
    .B(_10415_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand2_1 _15268_ (.A(_01606_),
    .B(_01617_),
    .Y(_01628_));
 sky130_fd_sc_hd__nand2_1 _15269_ (.A(_01628_),
    .B(_10701_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand3_1 _15270_ (.A(_01606_),
    .B(_10690_),
    .C(_01617_),
    .Y(_01650_));
 sky130_fd_sc_hd__nand2_1 _15271_ (.A(_01639_),
    .B(_01650_),
    .Y(_01661_));
 sky130_fd_sc_hd__nor2_2 _15272_ (.A(_01541_),
    .B(_01661_),
    .Y(_01672_));
 sky130_fd_sc_hd__nand2_1 _15273_ (.A(_10262_),
    .B(_10536_),
    .Y(_01683_));
 sky130_fd_sc_hd__nand2b_1 _15274_ (.A_N(_01409_),
    .B(_01683_),
    .Y(_01694_));
 sky130_fd_sc_hd__nand2_1 _15275_ (.A(_01694_),
    .B(_01552_),
    .Y(_01705_));
 sky130_fd_sc_hd__nand2_1 _15276_ (.A(_01705_),
    .B(_13104_),
    .Y(_01716_));
 sky130_fd_sc_hd__nand2_1 _15277_ (.A(_00992_),
    .B(_10196_),
    .Y(_01727_));
 sky130_fd_sc_hd__nand2_1 _15278_ (.A(_01716_),
    .B(_01727_),
    .Y(_01738_));
 sky130_fd_sc_hd__inv_2 _15279_ (.A(_01738_),
    .Y(_01749_));
 sky130_fd_sc_hd__nand2_1 _15280_ (.A(_01749_),
    .B(_10470_),
    .Y(_01760_));
 sky130_fd_sc_hd__nand2_1 _15281_ (.A(_01738_),
    .B(_10481_),
    .Y(_01771_));
 sky130_fd_sc_hd__nand2_1 _15282_ (.A(_01760_),
    .B(_01771_),
    .Y(_01782_));
 sky130_fd_sc_hd__nand2_1 _15283_ (.A(_01189_),
    .B(_09756_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand2_1 _15284_ (.A(_01793_),
    .B(_12842_),
    .Y(_01804_));
 sky130_fd_sc_hd__nand3_1 _15285_ (.A(_01189_),
    .B(_10031_),
    .C(_09756_),
    .Y(_01815_));
 sky130_fd_sc_hd__nand2_1 _15286_ (.A(_01804_),
    .B(_01815_),
    .Y(_01826_));
 sky130_fd_sc_hd__nand2_1 _15287_ (.A(_01826_),
    .B(\div1i.quot[23] ),
    .Y(_01837_));
 sky130_fd_sc_hd__nand2_1 _15288_ (.A(_00992_),
    .B(_09921_),
    .Y(_01848_));
 sky130_fd_sc_hd__nand2_1 _15289_ (.A(_01837_),
    .B(_01848_),
    .Y(_01859_));
 sky130_fd_sc_hd__nand2_1 _15290_ (.A(_01859_),
    .B(_10251_),
    .Y(_01870_));
 sky130_fd_sc_hd__nand3_2 _15291_ (.A(_01837_),
    .B(_10240_),
    .C(_01848_),
    .Y(_01881_));
 sky130_fd_sc_hd__nand2_1 _15292_ (.A(_01870_),
    .B(_01881_),
    .Y(_01892_));
 sky130_fd_sc_hd__nor2_1 _15293_ (.A(_01782_),
    .B(_01892_),
    .Y(_01903_));
 sky130_fd_sc_hd__nand2_1 _15294_ (.A(_01672_),
    .B(_01903_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_4 _15295_ (.A(_01376_),
    .B(_01914_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2_2 _15296_ (.A(_00860_),
    .B(_01925_),
    .Y(_01936_));
 sky130_fd_sc_hd__o21ai_1 _15297_ (.A1(_01650_),
    .A2(_01541_),
    .B1(_01530_),
    .Y(_01947_));
 sky130_fd_sc_hd__inv_2 _15298_ (.A(_01947_),
    .Y(_01958_));
 sky130_fd_sc_hd__inv_2 _15299_ (.A(_01771_),
    .Y(_01969_));
 sky130_fd_sc_hd__o21ai_2 _15300_ (.A1(_01881_),
    .A2(_01969_),
    .B1(_01760_),
    .Y(_01980_));
 sky130_fd_sc_hd__nand2_1 _15301_ (.A(_01672_),
    .B(_01980_),
    .Y(_01991_));
 sky130_fd_sc_hd__nand2_1 _15302_ (.A(_01958_),
    .B(_01991_),
    .Y(_02002_));
 sky130_fd_sc_hd__a21o_1 _15303_ (.A1(_00948_),
    .A2(_01101_),
    .B1(_01090_),
    .X(_02013_));
 sky130_fd_sc_hd__o21ai_1 _15304_ (.A1(_01343_),
    .A2(_01266_),
    .B1(_01255_),
    .Y(_02024_));
 sky130_fd_sc_hd__a21oi_2 _15305_ (.A1(_02013_),
    .A2(_01365_),
    .B1(_02024_),
    .Y(_02035_));
 sky130_fd_sc_hd__nor2_1 _15306_ (.A(_01914_),
    .B(_02035_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_2 _15307_ (.A(_02002_),
    .B(_02046_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_1 _15308_ (.A(_01453_),
    .B(_10723_),
    .Y(_02068_));
 sky130_fd_sc_hd__xor2_1 _15309_ (.A(_10997_),
    .B(_02068_),
    .X(_02079_));
 sky130_fd_sc_hd__mux2_4 _15310_ (.A0(_02079_),
    .A1(_10876_),
    .S(_00992_),
    .X(_02090_));
 sky130_fd_sc_hd__nand3_4 _15311_ (.A(_01936_),
    .B(_02057_),
    .C(_02090_),
    .Y(_02101_));
 sky130_fd_sc_hd__buf_8 _15312_ (.A(_02101_),
    .X(_02112_));
 sky130_fd_sc_hd__buf_12 _15313_ (.A(_02112_),
    .X(\div1i.quot[22] ));
 sky130_fd_sc_hd__inv_4 _15314_ (.A(_02101_),
    .Y(_02133_));
 sky130_fd_sc_hd__buf_6 _15315_ (.A(_02133_),
    .X(_02142_));
 sky130_fd_sc_hd__nand2_1 _15316_ (.A(_02142_),
    .B(_00937_),
    .Y(_02153_));
 sky130_fd_sc_hd__inv_2 _15317_ (.A(_00981_),
    .Y(_02164_));
 sky130_fd_sc_hd__or2_1 _15318_ (.A(_02164_),
    .B(_00860_),
    .X(_02175_));
 sky130_fd_sc_hd__nand2_1 _15319_ (.A(_00860_),
    .B(_02164_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand2_1 _15320_ (.A(_02175_),
    .B(_02186_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _15321_ (.A(_02197_),
    .B(net132),
    .Y(_02208_));
 sky130_fd_sc_hd__nand2_1 _15322_ (.A(_02153_),
    .B(_02208_),
    .Y(_02219_));
 sky130_fd_sc_hd__nand2_1 _15323_ (.A(_02219_),
    .B(_09361_),
    .Y(_02230_));
 sky130_fd_sc_hd__nand3_1 _15324_ (.A(_02153_),
    .B(_02208_),
    .C(_09383_),
    .Y(_02241_));
 sky130_fd_sc_hd__nand2_1 _15325_ (.A(_02230_),
    .B(_02241_),
    .Y(_02252_));
 sky130_fd_sc_hd__inv_2 _15326_ (.A(_00640_),
    .Y(_02263_));
 sky130_fd_sc_hd__nand2_1 _15327_ (.A(_13983_),
    .B(_02263_),
    .Y(_02274_));
 sky130_fd_sc_hd__inv_2 _15328_ (.A(_00717_),
    .Y(_02285_));
 sky130_fd_sc_hd__nand2_1 _15329_ (.A(_02274_),
    .B(_02285_),
    .Y(_02296_));
 sky130_fd_sc_hd__nand2_1 _15330_ (.A(_02296_),
    .B(_14246_),
    .Y(_02307_));
 sky130_fd_sc_hd__inv_2 _15331_ (.A(_00794_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _15332_ (.A(_02307_),
    .B(_02318_),
    .Y(_02329_));
 sky130_fd_sc_hd__nand2_1 _15333_ (.A(_02329_),
    .B(_00739_),
    .Y(_02340_));
 sky130_fd_sc_hd__nand2_1 _15334_ (.A(_02340_),
    .B(_00212_),
    .Y(_02351_));
 sky130_fd_sc_hd__nand2_1 _15335_ (.A(_02351_),
    .B(_00728_),
    .Y(_02362_));
 sky130_fd_sc_hd__nand3_1 _15336_ (.A(_02340_),
    .B(_00135_),
    .C(_00212_),
    .Y(_02373_));
 sky130_fd_sc_hd__nand2_1 _15337_ (.A(_02362_),
    .B(_02373_),
    .Y(_02384_));
 sky130_fd_sc_hd__nand2_1 _15338_ (.A(_02384_),
    .B(\div1i.quot[22] ),
    .Y(_02395_));
 sky130_fd_sc_hd__buf_4 _15339_ (.A(_02133_),
    .X(_02406_));
 sky130_fd_sc_hd__nand2_1 _15340_ (.A(_02406_),
    .B(_00102_),
    .Y(_02417_));
 sky130_fd_sc_hd__nand3_2 _15341_ (.A(_02395_),
    .B(_09559_),
    .C(_02417_),
    .Y(_02428_));
 sky130_fd_sc_hd__o21ai_2 _15342_ (.A1(_02252_),
    .A2(_02428_),
    .B1(_02241_),
    .Y(_02439_));
 sky130_fd_sc_hd__nand2_1 _15343_ (.A(_02186_),
    .B(_00959_),
    .Y(_02450_));
 sky130_fd_sc_hd__xor2_1 _15344_ (.A(_01112_),
    .B(_02450_),
    .X(_02461_));
 sky130_fd_sc_hd__buf_8 _15345_ (.A(_02112_),
    .X(_02472_));
 sky130_fd_sc_hd__nand2_1 _15346_ (.A(_02461_),
    .B(_02472_),
    .Y(_02483_));
 sky130_fd_sc_hd__nand2_1 _15347_ (.A(_02142_),
    .B(_01079_),
    .Y(_02494_));
 sky130_fd_sc_hd__nand2_1 _15348_ (.A(_02483_),
    .B(_02494_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_1 _15349_ (.A(_02505_),
    .B(_09735_),
    .Y(_02516_));
 sky130_fd_sc_hd__nand3_2 _15350_ (.A(_02483_),
    .B(_09724_),
    .C(_02494_),
    .Y(_02527_));
 sky130_fd_sc_hd__nand2_1 _15351_ (.A(_02516_),
    .B(_02527_),
    .Y(_02538_));
 sky130_fd_sc_hd__inv_2 _15352_ (.A(_01354_),
    .Y(_02549_));
 sky130_fd_sc_hd__nand2_1 _15353_ (.A(_00860_),
    .B(_01123_),
    .Y(_02560_));
 sky130_fd_sc_hd__clkinvlp_2 _15354_ (.A(_02013_),
    .Y(_02571_));
 sky130_fd_sc_hd__nand2_1 _15355_ (.A(_02560_),
    .B(_02571_),
    .Y(_02582_));
 sky130_fd_sc_hd__or2_1 _15356_ (.A(_02549_),
    .B(_02582_),
    .X(_02593_));
 sky130_fd_sc_hd__nand2_1 _15357_ (.A(_02582_),
    .B(_02549_),
    .Y(_02604_));
 sky130_fd_sc_hd__nand2_1 _15358_ (.A(_02593_),
    .B(_02604_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _15359_ (.A(_02615_),
    .B(_02472_),
    .Y(_02626_));
 sky130_fd_sc_hd__nand2_1 _15360_ (.A(_02406_),
    .B(_01321_),
    .Y(_02637_));
 sky130_fd_sc_hd__nand2_1 _15361_ (.A(_02626_),
    .B(_02637_),
    .Y(_02648_));
 sky130_fd_sc_hd__nand2_1 _15362_ (.A(_02648_),
    .B(_09987_),
    .Y(_02658_));
 sky130_fd_sc_hd__nand3_1 _15363_ (.A(_02626_),
    .B(_10009_),
    .C(_02637_),
    .Y(_02669_));
 sky130_fd_sc_hd__nand2_1 _15364_ (.A(_02658_),
    .B(_02669_),
    .Y(_02680_));
 sky130_fd_sc_hd__nor2_2 _15365_ (.A(_02680_),
    .B(_02538_),
    .Y(_02691_));
 sky130_fd_sc_hd__nand2_1 _15366_ (.A(_02439_),
    .B(_02691_),
    .Y(_02702_));
 sky130_fd_sc_hd__inv_2 _15367_ (.A(_02527_),
    .Y(_02713_));
 sky130_fd_sc_hd__a21boi_2 _15368_ (.A1(_02713_),
    .A2(_02658_),
    .B1_N(_02669_),
    .Y(_02724_));
 sky130_fd_sc_hd__nand2_1 _15369_ (.A(_02702_),
    .B(_02724_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand2_1 _15370_ (.A(_02604_),
    .B(_01343_),
    .Y(_02746_));
 sky130_fd_sc_hd__inv_2 _15371_ (.A(_01266_),
    .Y(_02757_));
 sky130_fd_sc_hd__nand2_1 _15372_ (.A(_02746_),
    .B(_02757_),
    .Y(_02767_));
 sky130_fd_sc_hd__nand3_1 _15373_ (.A(_02604_),
    .B(_01266_),
    .C(_01343_),
    .Y(_02778_));
 sky130_fd_sc_hd__nand2_1 _15374_ (.A(_02767_),
    .B(_02778_),
    .Y(_02789_));
 sky130_fd_sc_hd__nand2_1 _15375_ (.A(_02789_),
    .B(\div1i.quot[22] ),
    .Y(_02800_));
 sky130_fd_sc_hd__nand2_1 _15376_ (.A(_02406_),
    .B(_01233_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand2_1 _15377_ (.A(_02800_),
    .B(_02811_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _15378_ (.A(_02822_),
    .B(_10251_),
    .Y(_02833_));
 sky130_fd_sc_hd__inv_2 _15379_ (.A(_01376_),
    .Y(_02844_));
 sky130_fd_sc_hd__nand2_1 _15380_ (.A(_00860_),
    .B(_02844_),
    .Y(_02855_));
 sky130_fd_sc_hd__nand2_1 _15381_ (.A(_02855_),
    .B(_02035_),
    .Y(_02866_));
 sky130_fd_sc_hd__inv_2 _15382_ (.A(_01892_),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_1 _15383_ (.A(_02866_),
    .B(_02876_),
    .Y(_02887_));
 sky130_fd_sc_hd__nand3_1 _15384_ (.A(_02855_),
    .B(_01892_),
    .C(_02035_),
    .Y(_02898_));
 sky130_fd_sc_hd__nand2_1 _15385_ (.A(_02887_),
    .B(_02898_),
    .Y(_02909_));
 sky130_fd_sc_hd__nand2_1 _15386_ (.A(_02909_),
    .B(net132),
    .Y(_02920_));
 sky130_fd_sc_hd__nand2_1 _15387_ (.A(_02142_),
    .B(_01859_),
    .Y(_02931_));
 sky130_fd_sc_hd__nand2_1 _15388_ (.A(_02920_),
    .B(_02931_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2_1 _15389_ (.A(_02942_),
    .B(_10481_),
    .Y(_02953_));
 sky130_fd_sc_hd__nand3_1 _15390_ (.A(_02920_),
    .B(_10470_),
    .C(_02931_),
    .Y(_02964_));
 sky130_fd_sc_hd__nand2_1 _15391_ (.A(_02953_),
    .B(_02964_),
    .Y(_02974_));
 sky130_fd_sc_hd__inv_2 _15392_ (.A(_02974_),
    .Y(_02985_));
 sky130_fd_sc_hd__nand3_2 _15393_ (.A(_02800_),
    .B(_10240_),
    .C(_02811_),
    .Y(_02996_));
 sky130_fd_sc_hd__nand3_2 _15394_ (.A(_02833_),
    .B(_02985_),
    .C(_02996_),
    .Y(_03007_));
 sky130_fd_sc_hd__nand2_1 _15395_ (.A(_02887_),
    .B(_01881_),
    .Y(_03018_));
 sky130_fd_sc_hd__inv_2 _15396_ (.A(_01782_),
    .Y(_03029_));
 sky130_fd_sc_hd__nand2_1 _15397_ (.A(_03018_),
    .B(_03029_),
    .Y(_03040_));
 sky130_fd_sc_hd__nand3_1 _15398_ (.A(_02887_),
    .B(_01782_),
    .C(_01881_),
    .Y(_03051_));
 sky130_fd_sc_hd__nand2_1 _15399_ (.A(_03040_),
    .B(_03051_),
    .Y(_03062_));
 sky130_fd_sc_hd__nand2_1 _15400_ (.A(_03062_),
    .B(_02472_),
    .Y(_03073_));
 sky130_fd_sc_hd__nand2_1 _15401_ (.A(_02142_),
    .B(_01738_),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2_1 _15402_ (.A(_03073_),
    .B(_03084_),
    .Y(_03094_));
 sky130_fd_sc_hd__nand2_1 _15403_ (.A(_03094_),
    .B(_10701_),
    .Y(_03105_));
 sky130_fd_sc_hd__nand3_1 _15404_ (.A(_03073_),
    .B(_10690_),
    .C(_03084_),
    .Y(_03116_));
 sky130_fd_sc_hd__nand2_1 _15405_ (.A(_03105_),
    .B(_03116_),
    .Y(_03127_));
 sky130_fd_sc_hd__inv_2 _15406_ (.A(_03127_),
    .Y(_03138_));
 sky130_fd_sc_hd__nand2_1 _15407_ (.A(_02866_),
    .B(_01903_),
    .Y(_03149_));
 sky130_fd_sc_hd__inv_2 _15408_ (.A(_01980_),
    .Y(_03160_));
 sky130_fd_sc_hd__nand2_1 _15409_ (.A(_03149_),
    .B(_03160_),
    .Y(_03171_));
 sky130_fd_sc_hd__clkinvlp_2 _15410_ (.A(_01661_),
    .Y(_03182_));
 sky130_fd_sc_hd__nand2_1 _15411_ (.A(_03171_),
    .B(_03182_),
    .Y(_03192_));
 sky130_fd_sc_hd__nand3_1 _15412_ (.A(_03149_),
    .B(_01661_),
    .C(_03160_),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2_1 _15413_ (.A(_03192_),
    .B(_03203_),
    .Y(_03214_));
 sky130_fd_sc_hd__nand2_1 _15414_ (.A(_03214_),
    .B(\div1i.quot[22] ),
    .Y(_03225_));
 sky130_fd_sc_hd__nand2_1 _15415_ (.A(_02406_),
    .B(_01628_),
    .Y(_03236_));
 sky130_fd_sc_hd__nand2_1 _15416_ (.A(_03225_),
    .B(_03236_),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _15417_ (.A(_03247_),
    .B(_10887_),
    .Y(_03258_));
 sky130_fd_sc_hd__nand3_1 _15418_ (.A(_03225_),
    .B(_10909_),
    .C(_03236_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand2_1 _15419_ (.A(_03258_),
    .B(_03269_),
    .Y(_03280_));
 sky130_fd_sc_hd__nand2_1 _15420_ (.A(_03138_),
    .B(_03280_),
    .Y(_03290_));
 sky130_fd_sc_hd__nor2_1 _15421_ (.A(_03007_),
    .B(_03290_),
    .Y(_03301_));
 sky130_fd_sc_hd__nand2_1 _15422_ (.A(_02735_),
    .B(_03301_),
    .Y(_03312_));
 sky130_fd_sc_hd__nand2_1 _15423_ (.A(_03247_),
    .B(_10909_),
    .Y(_03323_));
 sky130_fd_sc_hd__nand3_1 _15424_ (.A(_03225_),
    .B(_10887_),
    .C(_03236_),
    .Y(_03333_));
 sky130_fd_sc_hd__nand2_1 _15425_ (.A(_03323_),
    .B(_03333_),
    .Y(_03344_));
 sky130_fd_sc_hd__nor2_1 _15426_ (.A(_03344_),
    .B(_03127_),
    .Y(_03355_));
 sky130_fd_sc_hd__o21ai_1 _15427_ (.A1(_02974_),
    .A2(_02996_),
    .B1(_02964_),
    .Y(_03366_));
 sky130_fd_sc_hd__a21oi_1 _15428_ (.A1(_03225_),
    .A2(_03236_),
    .B1(_10887_),
    .Y(_03377_));
 sky130_fd_sc_hd__o21ai_1 _15429_ (.A1(_03116_),
    .A2(_03377_),
    .B1(_03333_),
    .Y(_03388_));
 sky130_fd_sc_hd__a21oi_1 _15430_ (.A1(_03355_),
    .A2(_03366_),
    .B1(_03388_),
    .Y(_03399_));
 sky130_fd_sc_hd__nand2_2 _15431_ (.A(_03312_),
    .B(_03399_),
    .Y(_03410_));
 sky130_fd_sc_hd__inv_1 _15432_ (.A(_03410_),
    .Y(_03421_));
 sky130_fd_sc_hd__nand3_1 _15433_ (.A(_02307_),
    .B(_00223_),
    .C(_02318_),
    .Y(_03432_));
 sky130_fd_sc_hd__nand2_1 _15434_ (.A(_02340_),
    .B(_03432_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand2_1 _15435_ (.A(_03443_),
    .B(net132),
    .Y(_03454_));
 sky130_fd_sc_hd__nand2_1 _15436_ (.A(_02142_),
    .B(_00190_),
    .Y(_03465_));
 sky130_fd_sc_hd__nand2_1 _15437_ (.A(_03454_),
    .B(_03465_),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _15438_ (.A(_03476_),
    .B(_08582_),
    .Y(_03487_));
 sky130_fd_sc_hd__nand3_1 _15439_ (.A(_03454_),
    .B(_08571_),
    .C(_03465_),
    .Y(_03498_));
 sky130_fd_sc_hd__nand2_1 _15440_ (.A(_03487_),
    .B(_03498_),
    .Y(_03509_));
 sky130_fd_sc_hd__nand2_1 _15441_ (.A(_02296_),
    .B(_14115_),
    .Y(_03520_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(_03520_),
    .B(_14093_),
    .Y(_03531_));
 sky130_fd_sc_hd__nand2_1 _15443_ (.A(_03531_),
    .B(_14224_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand3_1 _15444_ (.A(_03520_),
    .B(_14213_),
    .C(_14093_),
    .Y(_03553_));
 sky130_fd_sc_hd__nand2_1 _15445_ (.A(_03542_),
    .B(_03553_),
    .Y(_03564_));
 sky130_fd_sc_hd__nand2_1 _15446_ (.A(_03564_),
    .B(_02472_),
    .Y(_03575_));
 sky130_fd_sc_hd__nand2_1 _15447_ (.A(_02406_),
    .B(_14181_),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_1 _15448_ (.A(_03575_),
    .B(_03586_),
    .Y(_03597_));
 sky130_fd_sc_hd__nand2_1 _15449_ (.A(_03597_),
    .B(_08527_),
    .Y(_03608_));
 sky130_fd_sc_hd__nand3_2 _15450_ (.A(_03575_),
    .B(_08505_),
    .C(_03586_),
    .Y(_03619_));
 sky130_fd_sc_hd__nand2_1 _15451_ (.A(_03608_),
    .B(_03619_),
    .Y(_03630_));
 sky130_fd_sc_hd__nor2_1 _15452_ (.A(_03509_),
    .B(_03630_),
    .Y(_03641_));
 sky130_fd_sc_hd__a21oi_1 _15453_ (.A1(_01672_),
    .A2(_01980_),
    .B1(_01947_),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2_1 _15454_ (.A(_02013_),
    .B(_01365_),
    .Y(_03663_));
 sky130_fd_sc_hd__inv_2 _15455_ (.A(_02024_),
    .Y(_03674_));
 sky130_fd_sc_hd__nand2_1 _15456_ (.A(_03663_),
    .B(_03674_),
    .Y(_03685_));
 sky130_fd_sc_hd__nand3_1 _15457_ (.A(_03685_),
    .B(_01672_),
    .C(_01903_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand2_1 _15458_ (.A(_03652_),
    .B(_03696_),
    .Y(_03707_));
 sky130_fd_sc_hd__a21oi_4 _15459_ (.A1(_00860_),
    .A2(_01925_),
    .B1(_03707_),
    .Y(_03718_));
 sky130_fd_sc_hd__nand3_1 _15460_ (.A(_03718_),
    .B(_14071_),
    .C(_02090_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand3_1 _15461_ (.A(_02274_),
    .B(_02285_),
    .C(_14104_),
    .Y(_03740_));
 sky130_fd_sc_hd__nand2_1 _15462_ (.A(_03520_),
    .B(_03740_),
    .Y(_03751_));
 sky130_fd_sc_hd__nand2_1 _15463_ (.A(_02112_),
    .B(_03751_),
    .Y(_03762_));
 sky130_fd_sc_hd__nand2_1 _15464_ (.A(_03729_),
    .B(_03762_),
    .Y(_03773_));
 sky130_fd_sc_hd__nand2_1 _15465_ (.A(_03773_),
    .B(_08384_),
    .Y(_03784_));
 sky130_fd_sc_hd__nand3_1 _15466_ (.A(_03729_),
    .B(_08406_),
    .C(_03762_),
    .Y(_03795_));
 sky130_fd_sc_hd__nand2_1 _15467_ (.A(_03784_),
    .B(_03795_),
    .Y(_03806_));
 sky130_fd_sc_hd__inv_4 _15468_ (.A(_03806_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand2_1 _15469_ (.A(_13983_),
    .B(_00443_),
    .Y(_03828_));
 sky130_fd_sc_hd__inv_2 _15470_ (.A(_00673_),
    .Y(_03839_));
 sky130_fd_sc_hd__nand2_1 _15471_ (.A(_03828_),
    .B(_03839_),
    .Y(_03850_));
 sky130_fd_sc_hd__inv_2 _15472_ (.A(_00618_),
    .Y(_03861_));
 sky130_fd_sc_hd__nand2_1 _15473_ (.A(_03850_),
    .B(_03861_),
    .Y(_03872_));
 sky130_fd_sc_hd__nand2_1 _15474_ (.A(_03872_),
    .B(_00607_),
    .Y(_03883_));
 sky130_fd_sc_hd__clkinvlp_2 _15475_ (.A(_00530_),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _15476_ (.A(_03883_),
    .B(_03894_),
    .Y(_03905_));
 sky130_fd_sc_hd__nand3_1 _15477_ (.A(_03872_),
    .B(_00530_),
    .C(_00607_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2_1 _15478_ (.A(_03905_),
    .B(_03916_),
    .Y(_03927_));
 sky130_fd_sc_hd__nand2_1 _15479_ (.A(_03927_),
    .B(_02472_),
    .Y(_03938_));
 sky130_fd_sc_hd__nand2_1 _15480_ (.A(_02142_),
    .B(_00498_),
    .Y(_03949_));
 sky130_fd_sc_hd__nand2_1 _15481_ (.A(_03938_),
    .B(_03949_),
    .Y(_03960_));
 sky130_fd_sc_hd__nand2_1 _15482_ (.A(_03960_),
    .B(_08274_),
    .Y(_03971_));
 sky130_fd_sc_hd__nand3_2 _15483_ (.A(_03938_),
    .B(_08296_),
    .C(_03949_),
    .Y(_03982_));
 sky130_fd_sc_hd__nand2_2 _15484_ (.A(_03971_),
    .B(_03982_),
    .Y(_03993_));
 sky130_fd_sc_hd__nor2_1 _15485_ (.A(_03817_),
    .B(_03993_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2_1 _15486_ (.A(_03641_),
    .B(_04004_),
    .Y(_04015_));
 sky130_fd_sc_hd__clkinv_1 _15487_ (.A(_04015_),
    .Y(_04026_));
 sky130_fd_sc_hd__nand3b_1 _15488_ (.A_N(_13566_),
    .B(_03718_),
    .C(_02090_),
    .Y(_04037_));
 sky130_fd_sc_hd__inv_2 _15489_ (.A(_13379_),
    .Y(_04048_));
 sky130_fd_sc_hd__o21bai_1 _15490_ (.A1(_13818_),
    .A2(_04048_),
    .B1_N(_13873_),
    .Y(_04059_));
 sky130_fd_sc_hd__nand2_1 _15491_ (.A(_04059_),
    .B(_13500_),
    .Y(_04070_));
 sky130_fd_sc_hd__nand2_1 _15492_ (.A(_04070_),
    .B(_13434_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand2_1 _15493_ (.A(_04081_),
    .B(_13610_),
    .Y(_04092_));
 sky130_fd_sc_hd__nand3_1 _15494_ (.A(_04070_),
    .B(_13928_),
    .C(_13434_),
    .Y(_04103_));
 sky130_fd_sc_hd__nand2_1 _15495_ (.A(_04092_),
    .B(_04103_),
    .Y(_04114_));
 sky130_fd_sc_hd__nand2_1 _15496_ (.A(_04114_),
    .B(\div1i.quot[22] ),
    .Y(_04125_));
 sky130_fd_sc_hd__nand3_1 _15497_ (.A(_04037_),
    .B(_08834_),
    .C(_04125_),
    .Y(_04136_));
 sky130_fd_sc_hd__clkinvlp_2 _15498_ (.A(_00300_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand3_1 _15499_ (.A(_03718_),
    .B(_04147_),
    .C(_02090_),
    .Y(_04158_));
 sky130_fd_sc_hd__inv_2 _15500_ (.A(_00333_),
    .Y(_04169_));
 sky130_fd_sc_hd__or2_1 _15501_ (.A(_04169_),
    .B(_13983_),
    .X(_04180_));
 sky130_fd_sc_hd__nand2_1 _15502_ (.A(_13983_),
    .B(_04169_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2_1 _15503_ (.A(_04180_),
    .B(_04191_),
    .Y(_04202_));
 sky130_fd_sc_hd__clkinvlp_2 _15504_ (.A(_04202_),
    .Y(_04213_));
 sky130_fd_sc_hd__nand2_1 _15505_ (.A(_02472_),
    .B(_04213_),
    .Y(_04224_));
 sky130_fd_sc_hd__nand3_2 _15506_ (.A(_04158_),
    .B(_08746_),
    .C(_04224_),
    .Y(_04234_));
 sky130_fd_sc_hd__inv_2 _15507_ (.A(_04234_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2_1 _15508_ (.A(_04158_),
    .B(_04224_),
    .Y(_04255_));
 sky130_fd_sc_hd__nand2_1 _15509_ (.A(_04255_),
    .B(_11140_),
    .Y(_04266_));
 sky130_fd_sc_hd__o21ai_1 _15510_ (.A1(_04136_),
    .A2(_04245_),
    .B1(_04266_),
    .Y(_04277_));
 sky130_fd_sc_hd__nand3_1 _15511_ (.A(_03718_),
    .B(_00585_),
    .C(_02090_),
    .Y(_04287_));
 sky130_fd_sc_hd__or2b_1 _15512_ (.A(_03850_),
    .B_N(_00618_),
    .X(_04298_));
 sky130_fd_sc_hd__nand2_1 _15513_ (.A(_04298_),
    .B(_03872_),
    .Y(_04308_));
 sky130_fd_sc_hd__nand2_1 _15514_ (.A(_04308_),
    .B(_02472_),
    .Y(_04319_));
 sky130_fd_sc_hd__nand2_1 _15515_ (.A(_04287_),
    .B(_04319_),
    .Y(_04330_));
 sky130_fd_sc_hd__nand2_2 _15516_ (.A(_04330_),
    .B(_08944_),
    .Y(_04340_));
 sky130_fd_sc_hd__nand3_1 _15517_ (.A(_04287_),
    .B(_04319_),
    .C(_08966_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2_2 _15518_ (.A(_04340_),
    .B(_04351_),
    .Y(_04361_));
 sky130_fd_sc_hd__inv_2 _15519_ (.A(_00399_),
    .Y(_04372_));
 sky130_fd_sc_hd__nand2_1 _15520_ (.A(_02406_),
    .B(_04372_),
    .Y(_04382_));
 sky130_fd_sc_hd__nand2_1 _15521_ (.A(_04191_),
    .B(_00322_),
    .Y(_04393_));
 sky130_fd_sc_hd__xor2_1 _15522_ (.A(_00432_),
    .B(_04393_),
    .X(_04404_));
 sky130_fd_sc_hd__nand2_1 _15523_ (.A(_04404_),
    .B(\div1i.quot[22] ),
    .Y(_04414_));
 sky130_fd_sc_hd__nand2_1 _15524_ (.A(_04382_),
    .B(_04414_),
    .Y(_04425_));
 sky130_fd_sc_hd__nand2_1 _15525_ (.A(_04425_),
    .B(_09054_),
    .Y(_04435_));
 sky130_fd_sc_hd__nand3_2 _15526_ (.A(_04382_),
    .B(_04414_),
    .C(_09076_),
    .Y(_04446_));
 sky130_fd_sc_hd__nand2_1 _15527_ (.A(_04435_),
    .B(_04446_),
    .Y(_04456_));
 sky130_fd_sc_hd__nor2_2 _15528_ (.A(_04361_),
    .B(_04456_),
    .Y(_04467_));
 sky130_fd_sc_hd__nand2_1 _15529_ (.A(_04277_),
    .B(_04467_),
    .Y(_04478_));
 sky130_fd_sc_hd__inv_2 _15530_ (.A(_04446_),
    .Y(_04488_));
 sky130_fd_sc_hd__a21boi_2 _15531_ (.A1(_04488_),
    .A2(_04340_),
    .B1_N(_04351_),
    .Y(_04499_));
 sky130_fd_sc_hd__nand2_2 _15532_ (.A(_04478_),
    .B(_04499_),
    .Y(_04509_));
 sky130_fd_sc_hd__a21oi_1 _15533_ (.A1(_03729_),
    .A2(_03762_),
    .B1(_08384_),
    .Y(_04520_));
 sky130_fd_sc_hd__or2_1 _15534_ (.A(_08406_),
    .B(_03773_),
    .X(_04530_));
 sky130_fd_sc_hd__o21ai_1 _15535_ (.A1(_04520_),
    .A2(_03982_),
    .B1(_04530_),
    .Y(_04541_));
 sky130_fd_sc_hd__nand2_1 _15536_ (.A(_03641_),
    .B(_04541_),
    .Y(_04552_));
 sky130_fd_sc_hd__inv_2 _15537_ (.A(_03619_),
    .Y(_04562_));
 sky130_fd_sc_hd__a21boi_1 _15538_ (.A1(_04562_),
    .A2(_03487_),
    .B1_N(_03498_),
    .Y(_04573_));
 sky130_fd_sc_hd__nand2_1 _15539_ (.A(_04552_),
    .B(_04573_),
    .Y(_04583_));
 sky130_fd_sc_hd__a21oi_2 _15540_ (.A1(_04026_),
    .A2(_04509_),
    .B1(_04583_),
    .Y(_04594_));
 sky130_fd_sc_hd__nand2_1 _15541_ (.A(_02133_),
    .B(_13280_),
    .Y(_04604_));
 sky130_fd_sc_hd__nand2_1 _15542_ (.A(_13192_),
    .B(_13236_),
    .Y(_04615_));
 sky130_fd_sc_hd__nand2_1 _15543_ (.A(_04615_),
    .B(_13094_),
    .Y(_04626_));
 sky130_fd_sc_hd__xor2_1 _15544_ (.A(_13313_),
    .B(_04626_),
    .X(_04636_));
 sky130_fd_sc_hd__inv_2 _15545_ (.A(_04636_),
    .Y(_04647_));
 sky130_fd_sc_hd__nand2_1 _15546_ (.A(_02112_),
    .B(_04647_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand3_1 _15547_ (.A(_04604_),
    .B(_07725_),
    .C(_04657_),
    .Y(_04668_));
 sky130_fd_sc_hd__inv_2 _15548_ (.A(_13675_),
    .Y(_04678_));
 sky130_fd_sc_hd__nand2_1 _15549_ (.A(_02406_),
    .B(_04678_),
    .Y(_04689_));
 sky130_fd_sc_hd__nand2_1 _15550_ (.A(_04048_),
    .B(_13708_),
    .Y(_04699_));
 sky130_fd_sc_hd__nand2_1 _15551_ (.A(_13379_),
    .B(_13719_),
    .Y(_04710_));
 sky130_fd_sc_hd__nand2_1 _15552_ (.A(_04699_),
    .B(_04710_),
    .Y(_04720_));
 sky130_fd_sc_hd__inv_2 _15553_ (.A(_04720_),
    .Y(_04731_));
 sky130_fd_sc_hd__nand2_1 _15554_ (.A(_02472_),
    .B(_04731_),
    .Y(_04741_));
 sky130_fd_sc_hd__nand3_1 _15555_ (.A(_04689_),
    .B(_04741_),
    .C(_12051_),
    .Y(_04752_));
 sky130_fd_sc_hd__inv_2 _15556_ (.A(_04752_),
    .Y(_04762_));
 sky130_fd_sc_hd__nand2_1 _15557_ (.A(_04689_),
    .B(_04741_),
    .Y(_04773_));
 sky130_fd_sc_hd__nand2_1 _15558_ (.A(_04773_),
    .B(_12029_),
    .Y(_04784_));
 sky130_fd_sc_hd__o21ai_1 _15559_ (.A1(_04668_),
    .A2(_04762_),
    .B1(_04784_),
    .Y(_04795_));
 sky130_fd_sc_hd__nand2_1 _15560_ (.A(_13412_),
    .B(_13423_),
    .Y(_04806_));
 sky130_fd_sc_hd__nand3b_1 _15561_ (.A_N(_04806_),
    .B(_03718_),
    .C(_02090_),
    .Y(_04817_));
 sky130_fd_sc_hd__or2_1 _15562_ (.A(_13500_),
    .B(_04059_),
    .X(_04828_));
 sky130_fd_sc_hd__nand2_1 _15563_ (.A(_04828_),
    .B(_04070_),
    .Y(_04839_));
 sky130_fd_sc_hd__inv_2 _15564_ (.A(_04839_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _15565_ (.A(_04850_),
    .B(_02472_),
    .Y(_04861_));
 sky130_fd_sc_hd__nand3_1 _15566_ (.A(_04817_),
    .B(_11579_),
    .C(_04861_),
    .Y(_04869_));
 sky130_fd_sc_hd__nand2_1 _15567_ (.A(_02406_),
    .B(_04806_),
    .Y(_04878_));
 sky130_fd_sc_hd__nand2_1 _15568_ (.A(\div1i.quot[22] ),
    .B(_04839_),
    .Y(_04889_));
 sky130_fd_sc_hd__nand3_1 _15569_ (.A(_04878_),
    .B(_13588_),
    .C(_04889_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2_1 _15570_ (.A(_04869_),
    .B(_04900_),
    .Y(_04911_));
 sky130_fd_sc_hd__inv_2 _15571_ (.A(_13774_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_1 _15572_ (.A(_02406_),
    .B(_04921_),
    .Y(_04926_));
 sky130_fd_sc_hd__nand2_1 _15573_ (.A(_04710_),
    .B(_13697_),
    .Y(_04927_));
 sky130_fd_sc_hd__xnor2_1 _15574_ (.A(_13807_),
    .B(_04927_),
    .Y(_04928_));
 sky130_fd_sc_hd__nand2_1 _15575_ (.A(\div1i.quot[22] ),
    .B(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_2 _15576_ (.A(_04926_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__nand2_1 _15577_ (.A(_04930_),
    .B(_08066_),
    .Y(_04931_));
 sky130_fd_sc_hd__nand3_2 _15578_ (.A(_04926_),
    .B(_08055_),
    .C(_04929_),
    .Y(_04932_));
 sky130_fd_sc_hd__nand2_2 _15579_ (.A(_04931_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__nor2_1 _15580_ (.A(_04911_),
    .B(_04933_),
    .Y(_04934_));
 sky130_fd_sc_hd__inv_2 _15581_ (.A(_04869_),
    .Y(_04935_));
 sky130_fd_sc_hd__o21ai_1 _15582_ (.A1(_04932_),
    .A2(_04935_),
    .B1(_04900_),
    .Y(_04936_));
 sky130_fd_sc_hd__a21oi_2 _15583_ (.A1(_04795_),
    .A2(_04934_),
    .B1(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__nand2_1 _15584_ (.A(_02142_),
    .B(_13203_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_1 _15585_ (.A(_13203_),
    .B(_07231_),
    .Y(_04939_));
 sky130_fd_sc_hd__nand2_1 _15586_ (.A(_13225_),
    .B(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__nand2_1 _15587_ (.A(_02112_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__nand3_2 _15588_ (.A(_04938_),
    .B(_07539_),
    .C(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hd__nand2_1 _15589_ (.A(_02142_),
    .B(_13214_),
    .Y(_04943_));
 sky130_fd_sc_hd__inv_2 _15590_ (.A(_04940_),
    .Y(_04944_));
 sky130_fd_sc_hd__nand2_1 _15591_ (.A(net132),
    .B(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hd__nand3_1 _15592_ (.A(_04943_),
    .B(_07560_),
    .C(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__nand2_1 _15593_ (.A(_04942_),
    .B(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__inv_2 _15594_ (.A(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__nand2_1 _15595_ (.A(_13017_),
    .B(_13083_),
    .Y(_04949_));
 sky130_fd_sc_hd__nand2_1 _15596_ (.A(_02142_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__nand2_1 _15597_ (.A(_13181_),
    .B(_13225_),
    .Y(_04951_));
 sky130_fd_sc_hd__nand2_1 _15598_ (.A(_04615_),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__nand2_2 _15599_ (.A(_02472_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__nand2_2 _15600_ (.A(_04950_),
    .B(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hd__nand2_1 _15601_ (.A(_04954_),
    .B(_11777_),
    .Y(_04955_));
 sky130_fd_sc_hd__nand3_1 _15602_ (.A(_04950_),
    .B(_11799_),
    .C(_04953_),
    .Y(_04956_));
 sky130_fd_sc_hd__nand2_1 _15603_ (.A(_04955_),
    .B(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__nand2_1 _15604_ (.A(_02101_),
    .B(_07308_),
    .Y(_04958_));
 sky130_fd_sc_hd__inv_2 _15605_ (.A(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__nand2_1 _15606_ (.A(_04959_),
    .B(_07242_),
    .Y(_04960_));
 sky130_fd_sc_hd__inv_2 _15607_ (.A(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand3_2 _15608_ (.A(_04948_),
    .B(_04957_),
    .C(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__clkinvlp_2 _15609_ (.A(_04942_),
    .Y(_04963_));
 sky130_fd_sc_hd__nand2_1 _15610_ (.A(_04954_),
    .B(_11799_),
    .Y(_04964_));
 sky130_fd_sc_hd__nand3_1 _15611_ (.A(_04950_),
    .B(_11777_),
    .C(_04953_),
    .Y(_04965_));
 sky130_fd_sc_hd__a21boi_1 _15612_ (.A1(_04963_),
    .A2(_04964_),
    .B1_N(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__nand2_2 _15613_ (.A(_04962_),
    .B(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__inv_2 _15614_ (.A(_13280_),
    .Y(_04968_));
 sky130_fd_sc_hd__nand2_1 _15615_ (.A(_02142_),
    .B(_04968_),
    .Y(_04969_));
 sky130_fd_sc_hd__nand2_1 _15616_ (.A(net132),
    .B(_04636_),
    .Y(_04970_));
 sky130_fd_sc_hd__nand3_1 _15617_ (.A(_04969_),
    .B(_07703_),
    .C(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__nand2_1 _15618_ (.A(_04668_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__inv_2 _15619_ (.A(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__nand2_1 _15620_ (.A(_04773_),
    .B(_12051_),
    .Y(_04974_));
 sky130_fd_sc_hd__nand2_1 _15621_ (.A(\div1i.quot[22] ),
    .B(_04720_),
    .Y(_04975_));
 sky130_fd_sc_hd__o21ai_2 _15622_ (.A1(_04678_),
    .A2(\div1i.quot[22] ),
    .B1(_04975_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2_1 _15623_ (.A(_04976_),
    .B(_12029_),
    .Y(_04977_));
 sky130_fd_sc_hd__nand2_1 _15624_ (.A(_04974_),
    .B(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__nand2_1 _15625_ (.A(_04973_),
    .B(_04978_),
    .Y(_04979_));
 sky130_fd_sc_hd__nand3_1 _15626_ (.A(_04817_),
    .B(_13588_),
    .C(_04861_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand3_1 _15627_ (.A(_04878_),
    .B(_11579_),
    .C(_04889_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2_1 _15628_ (.A(_04980_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__nand3_1 _15629_ (.A(_04982_),
    .B(_04932_),
    .C(_04931_),
    .Y(_04983_));
 sky130_fd_sc_hd__nor2_1 _15630_ (.A(_04979_),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__nand2_2 _15631_ (.A(_04967_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__nand2_4 _15632_ (.A(_04937_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__nand2_2 _15633_ (.A(_04266_),
    .B(_04234_),
    .Y(_04987_));
 sky130_fd_sc_hd__nand2_1 _15634_ (.A(_04037_),
    .B(_04125_),
    .Y(_04988_));
 sky130_fd_sc_hd__nand2_1 _15635_ (.A(_04988_),
    .B(_12260_),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_1 _15636_ (.A(_04989_),
    .B(_04136_),
    .Y(_04990_));
 sky130_fd_sc_hd__nor2_4 _15637_ (.A(_04987_),
    .B(_04990_),
    .Y(_04991_));
 sky130_fd_sc_hd__nand2_1 _15638_ (.A(_04467_),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__nor2_2 _15639_ (.A(_04015_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__nand2_4 _15640_ (.A(_04986_),
    .B(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__nand2_4 _15641_ (.A(_04594_),
    .B(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__nand2_1 _15642_ (.A(_02395_),
    .B(_02417_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand2_1 _15643_ (.A(_04996_),
    .B(_09548_),
    .Y(_04997_));
 sky130_fd_sc_hd__inv_2 _15644_ (.A(_02252_),
    .Y(_04998_));
 sky130_fd_sc_hd__nand3_2 _15645_ (.A(_04997_),
    .B(_04998_),
    .C(_02428_),
    .Y(_04999_));
 sky130_fd_sc_hd__inv_4 _15646_ (.A(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_1 _15647_ (.A(_05000_),
    .B(_02691_),
    .Y(_05001_));
 sky130_fd_sc_hd__inv_2 _15648_ (.A(_03007_),
    .Y(_05002_));
 sky130_fd_sc_hd__nand2_1 _15649_ (.A(_03355_),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hd__nor2_4 _15650_ (.A(_05001_),
    .B(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__nand2_2 _15651_ (.A(_04995_),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__nand2_1 _15652_ (.A(_03192_),
    .B(_01650_),
    .Y(_05006_));
 sky130_fd_sc_hd__xor2_1 _15653_ (.A(_01541_),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__mux2_4 _15654_ (.A0(_05007_),
    .A1(_01508_),
    .S(_02406_),
    .X(_05008_));
 sky130_fd_sc_hd__nand3_4 _15655_ (.A(_03421_),
    .B(_05005_),
    .C(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__buf_8 _15656_ (.A(_05009_),
    .X(_05010_));
 sky130_fd_sc_hd__buf_8 _15657_ (.A(_05010_),
    .X(\div1i.quot[21] ));
 sky130_fd_sc_hd__nand2_1 _15658_ (.A(_04995_),
    .B(_05000_),
    .Y(_05011_));
 sky130_fd_sc_hd__inv_2 _15659_ (.A(_02439_),
    .Y(_05012_));
 sky130_fd_sc_hd__nand2_1 _15660_ (.A(_05011_),
    .B(_05012_),
    .Y(_05013_));
 sky130_fd_sc_hd__nand2_1 _15661_ (.A(_05013_),
    .B(_02691_),
    .Y(_05014_));
 sky130_fd_sc_hd__nand2_1 _15662_ (.A(_05014_),
    .B(_02724_),
    .Y(_05015_));
 sky130_fd_sc_hd__nand2_1 _15663_ (.A(_05015_),
    .B(_05002_),
    .Y(_05016_));
 sky130_fd_sc_hd__inv_2 _15664_ (.A(_03366_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_1 _15665_ (.A(_05016_),
    .B(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__nand2_1 _15666_ (.A(_05018_),
    .B(_03138_),
    .Y(_05019_));
 sky130_fd_sc_hd__nand3_1 _15667_ (.A(_05016_),
    .B(_03127_),
    .C(_05017_),
    .Y(_05020_));
 sky130_fd_sc_hd__nand2_1 _15668_ (.A(_05019_),
    .B(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_1 _15669_ (.A(_05021_),
    .B(\div1i.quot[21] ),
    .Y(_05022_));
 sky130_fd_sc_hd__inv_6 _15670_ (.A(_05009_),
    .Y(_05023_));
 sky130_fd_sc_hd__buf_6 _15671_ (.A(_05023_),
    .X(_05024_));
 sky130_fd_sc_hd__nand2_1 _15672_ (.A(_05024_),
    .B(_03094_),
    .Y(_05025_));
 sky130_fd_sc_hd__nand2_1 _15673_ (.A(_05022_),
    .B(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hd__nand2_1 _15674_ (.A(_05026_),
    .B(_10909_),
    .Y(_05027_));
 sky130_fd_sc_hd__nand3_1 _15675_ (.A(_05022_),
    .B(_10887_),
    .C(_05025_),
    .Y(_05028_));
 sky130_fd_sc_hd__nand2_2 _15676_ (.A(_05027_),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hd__and3_1 _15677_ (.A(_04995_),
    .B(_02691_),
    .C(_05000_),
    .X(_05030_));
 sky130_fd_sc_hd__nand2_1 _15678_ (.A(_02833_),
    .B(_02996_),
    .Y(_05031_));
 sky130_fd_sc_hd__o21bai_2 _15679_ (.A1(_02735_),
    .A2(_05030_),
    .B1_N(_05031_),
    .Y(_05032_));
 sky130_fd_sc_hd__nand2_1 _15680_ (.A(_05032_),
    .B(_02996_),
    .Y(_05033_));
 sky130_fd_sc_hd__nand2_1 _15681_ (.A(_05033_),
    .B(_02985_),
    .Y(_05034_));
 sky130_fd_sc_hd__nand3_1 _15682_ (.A(_05032_),
    .B(_02974_),
    .C(_02996_),
    .Y(_05035_));
 sky130_fd_sc_hd__nand2_1 _15683_ (.A(_05034_),
    .B(_05035_),
    .Y(_05036_));
 sky130_fd_sc_hd__nand2_1 _15684_ (.A(_05036_),
    .B(\div1i.quot[21] ),
    .Y(_05037_));
 sky130_fd_sc_hd__nand2_1 _15685_ (.A(_05024_),
    .B(_02942_),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _15686_ (.A(_05037_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_1 _15687_ (.A(_05039_),
    .B(_10701_),
    .Y(_05040_));
 sky130_fd_sc_hd__nand3_2 _15688_ (.A(_05037_),
    .B(_10690_),
    .C(_05038_),
    .Y(_05041_));
 sky130_fd_sc_hd__nand2_1 _15689_ (.A(_05040_),
    .B(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__nor2_1 _15690_ (.A(_05029_),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__inv_2 _15691_ (.A(_02538_),
    .Y(_05044_));
 sky130_fd_sc_hd__nand2_1 _15692_ (.A(_05013_),
    .B(_05044_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_1 _15693_ (.A(_05045_),
    .B(_02527_),
    .Y(_05046_));
 sky130_fd_sc_hd__xor2_1 _15694_ (.A(_02680_),
    .B(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__nand2_1 _15695_ (.A(_05047_),
    .B(_05010_),
    .Y(_05048_));
 sky130_fd_sc_hd__nand2_1 _15696_ (.A(_05023_),
    .B(_02648_),
    .Y(_05049_));
 sky130_fd_sc_hd__nand2_1 _15697_ (.A(_05048_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__or2_1 _15698_ (.A(_10251_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__nand3_1 _15699_ (.A(_05014_),
    .B(_05031_),
    .C(_02724_),
    .Y(_05052_));
 sky130_fd_sc_hd__nand2_1 _15700_ (.A(_05032_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__nand2_1 _15701_ (.A(_05053_),
    .B(net234),
    .Y(_05054_));
 sky130_fd_sc_hd__nand2_1 _15702_ (.A(_05023_),
    .B(_02822_),
    .Y(_05055_));
 sky130_fd_sc_hd__nand2_1 _15703_ (.A(_05054_),
    .B(_05055_),
    .Y(_05056_));
 sky130_fd_sc_hd__nand2_1 _15704_ (.A(_05056_),
    .B(_10481_),
    .Y(_05057_));
 sky130_fd_sc_hd__nand3_1 _15705_ (.A(_05054_),
    .B(_10470_),
    .C(_05055_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand2_2 _15706_ (.A(_05057_),
    .B(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__inv_2 _15707_ (.A(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_1 _15708_ (.A(_05050_),
    .B(_10251_),
    .Y(_05061_));
 sky130_fd_sc_hd__nand3_1 _15709_ (.A(_05051_),
    .B(_05060_),
    .C(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__inv_2 _15710_ (.A(_05062_),
    .Y(_05063_));
 sky130_fd_sc_hd__nand2_1 _15711_ (.A(_05043_),
    .B(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__clkinv_1 _15712_ (.A(_05064_),
    .Y(_05065_));
 sky130_fd_sc_hd__nand3_1 _15713_ (.A(_04986_),
    .B(_04467_),
    .C(_04991_),
    .Y(_05066_));
 sky130_fd_sc_hd__inv_2 _15714_ (.A(_04509_),
    .Y(_05067_));
 sky130_fd_sc_hd__nand2_1 _15715_ (.A(_05066_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hd__nand2_1 _15716_ (.A(_05068_),
    .B(_04004_),
    .Y(_05069_));
 sky130_fd_sc_hd__inv_2 _15717_ (.A(_04541_),
    .Y(_05070_));
 sky130_fd_sc_hd__nand2_1 _15718_ (.A(_05069_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__inv_2 _15719_ (.A(_03630_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_1 _15720_ (.A(_05071_),
    .B(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand2_1 _15721_ (.A(_05073_),
    .B(_03619_),
    .Y(_05074_));
 sky130_fd_sc_hd__xor2_1 _15722_ (.A(_03509_),
    .B(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__nand2_1 _15723_ (.A(_05075_),
    .B(\div1i.quot[21] ),
    .Y(_05076_));
 sky130_fd_sc_hd__nand2_1 _15724_ (.A(_05024_),
    .B(_03476_),
    .Y(_05077_));
 sky130_fd_sc_hd__nand3_2 _15725_ (.A(_05076_),
    .B(_09559_),
    .C(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hd__nand2_1 _15726_ (.A(_04997_),
    .B(_02428_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2b_1 _15727_ (.A_N(_05079_),
    .B(_04995_),
    .Y(_05080_));
 sky130_fd_sc_hd__or2b_1 _15728_ (.A(_04995_),
    .B_N(_05079_),
    .X(_05081_));
 sky130_fd_sc_hd__a21o_1 _15729_ (.A1(_05080_),
    .A2(_05081_),
    .B1(_05023_),
    .X(_05082_));
 sky130_fd_sc_hd__nand2_1 _15730_ (.A(_05023_),
    .B(_04996_),
    .Y(_05083_));
 sky130_fd_sc_hd__nand2_1 _15731_ (.A(_05082_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__nand2b_1 _15732_ (.A_N(_05084_),
    .B(_09383_),
    .Y(_05085_));
 sky130_fd_sc_hd__nand2_1 _15733_ (.A(_05084_),
    .B(_09361_),
    .Y(_05086_));
 sky130_fd_sc_hd__nand2_1 _15734_ (.A(_05085_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__o21ai_1 _15735_ (.A1(_05078_),
    .A2(_05087_),
    .B1(_05085_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(_05080_),
    .B(_02428_),
    .Y(_05089_));
 sky130_fd_sc_hd__or2_1 _15737_ (.A(_04998_),
    .B(_05089_),
    .X(_05090_));
 sky130_fd_sc_hd__nand2_1 _15738_ (.A(_05089_),
    .B(_04998_),
    .Y(_05091_));
 sky130_fd_sc_hd__a21o_1 _15739_ (.A1(_05090_),
    .A2(_05091_),
    .B1(_05024_),
    .X(_05092_));
 sky130_fd_sc_hd__nand2_1 _15740_ (.A(_05024_),
    .B(_02219_),
    .Y(_05093_));
 sky130_fd_sc_hd__nand2_1 _15741_ (.A(_05092_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__nand2_1 _15742_ (.A(_05094_),
    .B(_09735_),
    .Y(_05095_));
 sky130_fd_sc_hd__nand3_2 _15743_ (.A(_05092_),
    .B(net120),
    .C(_05093_),
    .Y(_05096_));
 sky130_fd_sc_hd__nand2_1 _15744_ (.A(_05095_),
    .B(_05096_),
    .Y(_05097_));
 sky130_fd_sc_hd__or2_1 _15745_ (.A(_05044_),
    .B(_05013_),
    .X(_05098_));
 sky130_fd_sc_hd__a21o_1 _15746_ (.A1(_05098_),
    .A2(_05045_),
    .B1(_05023_),
    .X(_05099_));
 sky130_fd_sc_hd__nand2_1 _15747_ (.A(_05024_),
    .B(_02505_),
    .Y(_05100_));
 sky130_fd_sc_hd__nand2_1 _15748_ (.A(_05099_),
    .B(_05100_),
    .Y(_05101_));
 sky130_fd_sc_hd__or2_1 _15749_ (.A(_09987_),
    .B(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__nand2_1 _15750_ (.A(_05101_),
    .B(_09987_),
    .Y(_05103_));
 sky130_fd_sc_hd__nand2_1 _15751_ (.A(_05102_),
    .B(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hd__nor2_1 _15752_ (.A(_05097_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__nand2_1 _15753_ (.A(_05088_),
    .B(_05105_),
    .Y(_05106_));
 sky130_fd_sc_hd__and2_1 _15754_ (.A(_05101_),
    .B(_09987_),
    .X(_05107_));
 sky130_fd_sc_hd__o21a_1 _15755_ (.A1(_05096_),
    .A2(_05107_),
    .B1(_05102_),
    .X(_05108_));
 sky130_fd_sc_hd__nand2_1 _15756_ (.A(_05106_),
    .B(_05108_),
    .Y(_05109_));
 sky130_fd_sc_hd__o21ai_1 _15757_ (.A1(_05059_),
    .A2(_05051_),
    .B1(_05058_),
    .Y(_05110_));
 sky130_fd_sc_hd__nand2_1 _15758_ (.A(_05110_),
    .B(_05043_),
    .Y(_05111_));
 sky130_fd_sc_hd__inv_2 _15759_ (.A(_05027_),
    .Y(_05112_));
 sky130_fd_sc_hd__o21a_1 _15760_ (.A1(_05041_),
    .A2(_05112_),
    .B1(_05028_),
    .X(_05113_));
 sky130_fd_sc_hd__nand2_1 _15761_ (.A(_05111_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hd__a21oi_4 _15762_ (.A1(_05065_),
    .A2(_05109_),
    .B1(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__or2_1 _15763_ (.A(_04255_),
    .B(_05010_),
    .X(_05116_));
 sky130_fd_sc_hd__nand2b_1 _15764_ (.A_N(_04990_),
    .B(_04986_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_1 _15765_ (.A(_05117_),
    .B(_04136_),
    .Y(_05118_));
 sky130_fd_sc_hd__xor2_1 _15766_ (.A(_04987_),
    .B(_05118_),
    .X(_05119_));
 sky130_fd_sc_hd__buf_6 _15767_ (.A(_05010_),
    .X(_05120_));
 sky130_fd_sc_hd__nand2_1 _15768_ (.A(_05119_),
    .B(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand2_1 _15769_ (.A(_05116_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__or2_4 _15770_ (.A(_09054_),
    .B(_05122_),
    .X(_05123_));
 sky130_fd_sc_hd__nand2_1 _15771_ (.A(_04986_),
    .B(_04991_),
    .Y(_05124_));
 sky130_fd_sc_hd__inv_2 _15772_ (.A(_04277_),
    .Y(_05125_));
 sky130_fd_sc_hd__nand2_1 _15773_ (.A(_05124_),
    .B(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__inv_2 _15774_ (.A(_04456_),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _15775_ (.A(_05126_),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__or2_1 _15776_ (.A(_05127_),
    .B(_05126_),
    .X(_05129_));
 sky130_fd_sc_hd__a21o_1 _15777_ (.A1(_05128_),
    .A2(_05129_),
    .B1(_05023_),
    .X(_05130_));
 sky130_fd_sc_hd__nand2_1 _15778_ (.A(_05024_),
    .B(_04425_),
    .Y(_05131_));
 sky130_fd_sc_hd__nand2_1 _15779_ (.A(_05130_),
    .B(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand2_1 _15780_ (.A(_05132_),
    .B(_08944_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand3_1 _15781_ (.A(_05130_),
    .B(_08966_),
    .C(_05131_),
    .Y(_05134_));
 sky130_fd_sc_hd__nand2_2 _15782_ (.A(_05133_),
    .B(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hd__o21a_1 _15783_ (.A1(_05123_),
    .A2(_05135_),
    .B1(_05134_),
    .X(_05136_));
 sky130_fd_sc_hd__nand2_1 _15784_ (.A(_05122_),
    .B(_09054_),
    .Y(_05137_));
 sky130_fd_sc_hd__nand2_2 _15785_ (.A(_05123_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__nor2_1 _15786_ (.A(_05135_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__inv_2 _15787_ (.A(_04967_),
    .Y(_05140_));
 sky130_fd_sc_hd__o21bai_1 _15788_ (.A1(_04979_),
    .A2(_05140_),
    .B1_N(_04795_),
    .Y(_05141_));
 sky130_fd_sc_hd__nand2b_1 _15789_ (.A_N(_04933_),
    .B(_05141_),
    .Y(_05142_));
 sky130_fd_sc_hd__nand2_1 _15790_ (.A(_05142_),
    .B(_04932_),
    .Y(_05143_));
 sky130_fd_sc_hd__xor2_1 _15791_ (.A(_04911_),
    .B(_05143_),
    .X(_05144_));
 sky130_fd_sc_hd__nand2_1 _15792_ (.A(_05144_),
    .B(\div1i.quot[21] ),
    .Y(_05145_));
 sky130_fd_sc_hd__a21o_1 _15793_ (.A1(_04878_),
    .A2(_04889_),
    .B1(_05120_),
    .X(_05146_));
 sky130_fd_sc_hd__nand3_2 _15794_ (.A(_05145_),
    .B(_05146_),
    .C(_08834_),
    .Y(_05147_));
 sky130_fd_sc_hd__nand2_1 _15795_ (.A(_05023_),
    .B(_04988_),
    .Y(_05148_));
 sky130_fd_sc_hd__or2b_1 _15796_ (.A(_04986_),
    .B_N(_04990_),
    .X(_05149_));
 sky130_fd_sc_hd__nand2_1 _15797_ (.A(_05149_),
    .B(_05117_),
    .Y(_05150_));
 sky130_fd_sc_hd__nand2_1 _15798_ (.A(_05120_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__a21o_1 _15799_ (.A1(_05148_),
    .A2(_05151_),
    .B1(_11140_),
    .X(_05152_));
 sky130_fd_sc_hd__inv_2 _15800_ (.A(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__and2_1 _15801_ (.A(_05148_),
    .B(_05151_),
    .X(_05154_));
 sky130_fd_sc_hd__nand2_1 _15802_ (.A(_05154_),
    .B(_11140_),
    .Y(_05155_));
 sky130_fd_sc_hd__o21ai_1 _15803_ (.A1(_05147_),
    .A2(_05153_),
    .B1(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__nand2_1 _15804_ (.A(_05139_),
    .B(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__nand2_1 _15805_ (.A(_05136_),
    .B(_05157_),
    .Y(_05158_));
 sky130_fd_sc_hd__clkinvlp_2 _15806_ (.A(_03993_),
    .Y(_05159_));
 sky130_fd_sc_hd__or2_1 _15807_ (.A(_05159_),
    .B(_05068_),
    .X(_05160_));
 sky130_fd_sc_hd__nand2_1 _15808_ (.A(_05068_),
    .B(_05159_),
    .Y(_05161_));
 sky130_fd_sc_hd__nand2_1 _15809_ (.A(_05160_),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_1 _15810_ (.A(_05162_),
    .B(_05120_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand2_1 _15811_ (.A(_05023_),
    .B(_03960_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand2_2 _15812_ (.A(_05163_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__or2_4 _15813_ (.A(_08406_),
    .B(_05165_),
    .X(_05166_));
 sky130_fd_sc_hd__nand2_1 _15814_ (.A(_05165_),
    .B(_08406_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand2_1 _15815_ (.A(_05166_),
    .B(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_1 _15816_ (.A(_05128_),
    .B(_04446_),
    .Y(_05170_));
 sky130_fd_sc_hd__xor2_1 _15817_ (.A(_04361_),
    .B(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nand2_1 _15818_ (.A(_05171_),
    .B(\div1i.quot[21] ),
    .Y(_05172_));
 sky130_fd_sc_hd__nand2_1 _15819_ (.A(_05024_),
    .B(_04330_),
    .Y(_05173_));
 sky130_fd_sc_hd__a21o_1 _15820_ (.A1(_05172_),
    .A2(_05173_),
    .B1(_08296_),
    .X(_05174_));
 sky130_fd_sc_hd__nand3_1 _15821_ (.A(_05172_),
    .B(_08296_),
    .C(_05173_),
    .Y(_05175_));
 sky130_fd_sc_hd__nand2_1 _15822_ (.A(_05174_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__nor2_1 _15823_ (.A(_05169_),
    .B(_05176_),
    .Y(_05177_));
 sky130_fd_sc_hd__nand2_1 _15824_ (.A(_05161_),
    .B(_03982_),
    .Y(_05179_));
 sky130_fd_sc_hd__xor2_1 _15825_ (.A(_03817_),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__nand2_1 _15826_ (.A(_05180_),
    .B(_05120_),
    .Y(_05181_));
 sky130_fd_sc_hd__nand2_1 _15827_ (.A(_05023_),
    .B(_03773_),
    .Y(_05182_));
 sky130_fd_sc_hd__nand2_1 _15828_ (.A(_05181_),
    .B(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__nand2_1 _15829_ (.A(_05183_),
    .B(_08527_),
    .Y(_05184_));
 sky130_fd_sc_hd__nand3_2 _15830_ (.A(_05181_),
    .B(_08505_),
    .C(_05182_),
    .Y(_05185_));
 sky130_fd_sc_hd__nand2_1 _15831_ (.A(_05184_),
    .B(_05185_),
    .Y(_05186_));
 sky130_fd_sc_hd__or2_1 _15832_ (.A(_05072_),
    .B(_05071_),
    .X(_05187_));
 sky130_fd_sc_hd__nand2_1 _15833_ (.A(_05187_),
    .B(_05073_),
    .Y(_05188_));
 sky130_fd_sc_hd__nand2_1 _15834_ (.A(_05188_),
    .B(\div1i.quot[21] ),
    .Y(_05190_));
 sky130_fd_sc_hd__nand2_1 _15835_ (.A(_05024_),
    .B(_03597_),
    .Y(_05191_));
 sky130_fd_sc_hd__nand2_1 _15836_ (.A(_05190_),
    .B(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__nand2_1 _15837_ (.A(_05192_),
    .B(net137),
    .Y(_05193_));
 sky130_fd_sc_hd__nand3_1 _15838_ (.A(_05190_),
    .B(net121),
    .C(_05191_),
    .Y(_05194_));
 sky130_fd_sc_hd__nand2_2 _15839_ (.A(_05193_),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__nor2_1 _15840_ (.A(_05186_),
    .B(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hd__and2_1 _15841_ (.A(_05177_),
    .B(_05196_),
    .X(_05197_));
 sky130_fd_sc_hd__o21a_1 _15842_ (.A1(_05185_),
    .A2(_05195_),
    .B1(_05194_),
    .X(_05198_));
 sky130_fd_sc_hd__inv_2 _15843_ (.A(_05168_),
    .Y(_05199_));
 sky130_fd_sc_hd__o21ai_1 _15844_ (.A1(_05199_),
    .A2(_05175_),
    .B1(_05166_),
    .Y(_05201_));
 sky130_fd_sc_hd__nand2_1 _15845_ (.A(_05196_),
    .B(_05201_),
    .Y(_05202_));
 sky130_fd_sc_hd__nand2_1 _15846_ (.A(_05198_),
    .B(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__a21oi_2 _15847_ (.A1(_05158_),
    .A2(_05197_),
    .B1(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__nand2_2 _15848_ (.A(_05152_),
    .B(_05155_),
    .Y(_05205_));
 sky130_fd_sc_hd__nand2_1 _15849_ (.A(_05145_),
    .B(_05146_),
    .Y(_05206_));
 sky130_fd_sc_hd__nand2_1 _15850_ (.A(_05206_),
    .B(_12260_),
    .Y(_05207_));
 sky130_fd_sc_hd__nand2_1 _15851_ (.A(_05207_),
    .B(_05147_),
    .Y(_05208_));
 sky130_fd_sc_hd__nor2_2 _15852_ (.A(_05205_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__and2_1 _15853_ (.A(_05139_),
    .B(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__a21oi_4 _15854_ (.A1(_04995_),
    .A2(_05004_),
    .B1(_03410_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand3_1 _15855_ (.A(_05212_),
    .B(_04954_),
    .C(_05008_),
    .Y(_05213_));
 sky130_fd_sc_hd__nand2_1 _15856_ (.A(_04948_),
    .B(_04961_),
    .Y(_05214_));
 sky130_fd_sc_hd__nand2_1 _15857_ (.A(_05214_),
    .B(_04942_),
    .Y(_05215_));
 sky130_fd_sc_hd__xor2_1 _15858_ (.A(_04957_),
    .B(_05215_),
    .X(_05216_));
 sky130_fd_sc_hd__inv_2 _15859_ (.A(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__nand2_1 _15860_ (.A(net234),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand3_2 _15861_ (.A(_05213_),
    .B(_05218_),
    .C(_07725_),
    .Y(_05219_));
 sky130_fd_sc_hd__buf_4 _15862_ (.A(_05212_),
    .X(_05220_));
 sky130_fd_sc_hd__nand2_1 _15863_ (.A(_04604_),
    .B(_04657_),
    .Y(_05221_));
 sky130_fd_sc_hd__inv_2 _15864_ (.A(_05221_),
    .Y(_05223_));
 sky130_fd_sc_hd__buf_6 _15865_ (.A(_05008_),
    .X(_05224_));
 sky130_fd_sc_hd__nand3_1 _15866_ (.A(_05220_),
    .B(_05223_),
    .C(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hd__xor2_1 _15867_ (.A(_04972_),
    .B(_04967_),
    .X(_05226_));
 sky130_fd_sc_hd__inv_2 _15868_ (.A(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__nand2_1 _15869_ (.A(_05120_),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__nand3_1 _15870_ (.A(_05225_),
    .B(_05228_),
    .C(_12051_),
    .Y(_05229_));
 sky130_fd_sc_hd__inv_2 _15871_ (.A(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hd__nand3_1 _15872_ (.A(_05220_),
    .B(_05221_),
    .C(_05224_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand2_1 _15873_ (.A(_05120_),
    .B(_05226_),
    .Y(_05232_));
 sky130_fd_sc_hd__nand3_1 _15874_ (.A(_05231_),
    .B(_05232_),
    .C(_12029_),
    .Y(_05234_));
 sky130_fd_sc_hd__o21ai_1 _15875_ (.A1(_05219_),
    .A2(_05230_),
    .B1(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__nand3_1 _15876_ (.A(_05220_),
    .B(_04976_),
    .C(_05224_),
    .Y(_05236_));
 sky130_fd_sc_hd__inv_2 _15877_ (.A(_04978_),
    .Y(_05237_));
 sky130_fd_sc_hd__o21ai_1 _15878_ (.A1(_04972_),
    .A2(_05140_),
    .B1(_04668_),
    .Y(_05238_));
 sky130_fd_sc_hd__xor2_1 _15879_ (.A(_05237_),
    .B(_05238_),
    .X(_05239_));
 sky130_fd_sc_hd__nand2_1 _15880_ (.A(net234),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__nand3_2 _15881_ (.A(_05236_),
    .B(_05240_),
    .C(_08055_),
    .Y(_05241_));
 sky130_fd_sc_hd__nand3_1 _15882_ (.A(_05220_),
    .B(_04773_),
    .C(_05224_),
    .Y(_05242_));
 sky130_fd_sc_hd__clkinvlp_2 _15883_ (.A(_05239_),
    .Y(_05243_));
 sky130_fd_sc_hd__nand2_1 _15884_ (.A(net234),
    .B(_05243_),
    .Y(_05245_));
 sky130_fd_sc_hd__nand3_1 _15885_ (.A(_05242_),
    .B(_05245_),
    .C(_08066_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand2_1 _15886_ (.A(_05241_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__nand3_1 _15887_ (.A(_05220_),
    .B(_04930_),
    .C(_05224_),
    .Y(_05248_));
 sky130_fd_sc_hd__or2b_1 _15888_ (.A(_05141_),
    .B_N(_04933_),
    .X(_05249_));
 sky130_fd_sc_hd__nand2_1 _15889_ (.A(_05249_),
    .B(_05142_),
    .Y(_05250_));
 sky130_fd_sc_hd__nand2_1 _15890_ (.A(_05120_),
    .B(_05250_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_2 _15891_ (.A(_05248_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__nand2_1 _15892_ (.A(_05252_),
    .B(_11579_),
    .Y(_05253_));
 sky130_fd_sc_hd__nand3_1 _15893_ (.A(_05248_),
    .B(_05251_),
    .C(_13588_),
    .Y(_05254_));
 sky130_fd_sc_hd__nand2_1 _15894_ (.A(_05253_),
    .B(_05254_),
    .Y(_05256_));
 sky130_fd_sc_hd__nor2_1 _15895_ (.A(_05247_),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__inv_2 _15896_ (.A(_05253_),
    .Y(_05258_));
 sky130_fd_sc_hd__o21ai_1 _15897_ (.A1(_05241_),
    .A2(_05258_),
    .B1(_05254_),
    .Y(_05259_));
 sky130_fd_sc_hd__a21oi_1 _15898_ (.A1(_05235_),
    .A2(_05257_),
    .B1(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand3_1 _15899_ (.A(_05220_),
    .B(_04958_),
    .C(_05224_),
    .Y(_05261_));
 sky130_fd_sc_hd__nand2_1 _15900_ (.A(_04958_),
    .B(_07231_),
    .Y(_05262_));
 sky130_fd_sc_hd__nand2_1 _15901_ (.A(_04960_),
    .B(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__nand2_1 _15902_ (.A(_05010_),
    .B(_05263_),
    .Y(_05264_));
 sky130_fd_sc_hd__nand3_2 _15903_ (.A(_05261_),
    .B(_05264_),
    .C(_07539_),
    .Y(_05265_));
 sky130_fd_sc_hd__nand3_1 _15904_ (.A(_05220_),
    .B(_04959_),
    .C(_05224_),
    .Y(_05267_));
 sky130_fd_sc_hd__inv_2 _15905_ (.A(_05263_),
    .Y(_05268_));
 sky130_fd_sc_hd__nand2_1 _15906_ (.A(_05120_),
    .B(_05268_),
    .Y(_05269_));
 sky130_fd_sc_hd__nand3_1 _15907_ (.A(_05267_),
    .B(_05269_),
    .C(_07560_),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2_1 _15908_ (.A(_05265_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__inv_2 _15909_ (.A(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__nand3_1 _15910_ (.A(_05120_),
    .B(_05474_),
    .C(_07308_),
    .Y(_05273_));
 sky130_fd_sc_hd__inv_2 _15911_ (.A(_05273_),
    .Y(_05274_));
 sky130_fd_sc_hd__nand2_1 _15912_ (.A(_04938_),
    .B(_04941_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand3b_1 _15913_ (.A_N(_05275_),
    .B(_05220_),
    .C(_05224_),
    .Y(_05276_));
 sky130_fd_sc_hd__nand2_1 _15914_ (.A(_04947_),
    .B(_04960_),
    .Y(_05278_));
 sky130_fd_sc_hd__nand2_1 _15915_ (.A(_05214_),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__inv_2 _15916_ (.A(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__nand2_1 _15917_ (.A(\div1i.quot[21] ),
    .B(_05280_),
    .Y(_05281_));
 sky130_fd_sc_hd__nand3_1 _15918_ (.A(_05276_),
    .B(_05281_),
    .C(_11777_),
    .Y(_05282_));
 sky130_fd_sc_hd__nand3_1 _15919_ (.A(_05220_),
    .B(_05275_),
    .C(_05224_),
    .Y(_05283_));
 sky130_fd_sc_hd__nand2_1 _15920_ (.A(\div1i.quot[21] ),
    .B(_05279_),
    .Y(_05284_));
 sky130_fd_sc_hd__nand3_1 _15921_ (.A(_05283_),
    .B(_05284_),
    .C(_11799_),
    .Y(_05285_));
 sky130_fd_sc_hd__nand2_2 _15922_ (.A(_05282_),
    .B(_05285_),
    .Y(_05286_));
 sky130_fd_sc_hd__nand3_1 _15923_ (.A(_05272_),
    .B(_05274_),
    .C(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__inv_2 _15924_ (.A(_05265_),
    .Y(_05289_));
 sky130_fd_sc_hd__nand3_2 _15925_ (.A(_05276_),
    .B(_05281_),
    .C(_11799_),
    .Y(_05290_));
 sky130_fd_sc_hd__nand3_1 _15926_ (.A(_05283_),
    .B(_05284_),
    .C(_11777_),
    .Y(_05291_));
 sky130_fd_sc_hd__a21boi_1 _15927_ (.A1(_05289_),
    .A2(_05290_),
    .B1_N(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hd__nand2_1 _15928_ (.A(_05287_),
    .B(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__clkinvlp_2 _15929_ (.A(_04954_),
    .Y(_05294_));
 sky130_fd_sc_hd__nand3_1 _15930_ (.A(_05220_),
    .B(_05294_),
    .C(_05224_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand2_1 _15931_ (.A(net234),
    .B(_05216_),
    .Y(_05296_));
 sky130_fd_sc_hd__nand3_1 _15932_ (.A(_05295_),
    .B(_05296_),
    .C(_07703_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand2_1 _15933_ (.A(_05297_),
    .B(_05219_),
    .Y(_05298_));
 sky130_fd_sc_hd__inv_2 _15934_ (.A(_05298_),
    .Y(_05300_));
 sky130_fd_sc_hd__nand2_1 _15935_ (.A(_05231_),
    .B(_05232_),
    .Y(_05301_));
 sky130_fd_sc_hd__nand2_1 _15936_ (.A(_05301_),
    .B(_12029_),
    .Y(_05302_));
 sky130_fd_sc_hd__nand3_1 _15937_ (.A(_05231_),
    .B(_05232_),
    .C(_12051_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand2_1 _15938_ (.A(_05302_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__nand2_1 _15939_ (.A(_05300_),
    .B(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__inv_2 _15940_ (.A(_05247_),
    .Y(_05306_));
 sky130_fd_sc_hd__nand2_1 _15941_ (.A(_05252_),
    .B(_13588_),
    .Y(_05307_));
 sky130_fd_sc_hd__nand3_1 _15942_ (.A(_05248_),
    .B(_05251_),
    .C(_11579_),
    .Y(_05308_));
 sky130_fd_sc_hd__nand2_1 _15943_ (.A(_05307_),
    .B(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__nand2_1 _15944_ (.A(_05306_),
    .B(_05309_),
    .Y(_05311_));
 sky130_fd_sc_hd__nor2_1 _15945_ (.A(_05305_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2_1 _15946_ (.A(_05293_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__nand2_2 _15947_ (.A(_05260_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__nand3_1 _15948_ (.A(_05197_),
    .B(_05210_),
    .C(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_2 _15949_ (.A(_05204_),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__a21o_1 _15950_ (.A1(_05076_),
    .A2(_05077_),
    .B1(_09559_),
    .X(_05317_));
 sky130_fd_sc_hd__inv_2 _15951_ (.A(_05087_),
    .Y(_05318_));
 sky130_fd_sc_hd__nand3_1 _15952_ (.A(_05317_),
    .B(_05318_),
    .C(_05078_),
    .Y(_05319_));
 sky130_fd_sc_hd__inv_2 _15953_ (.A(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__nand2_1 _15954_ (.A(_05320_),
    .B(_05105_),
    .Y(_05322_));
 sky130_fd_sc_hd__nor2_2 _15955_ (.A(_05064_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__nand2_4 _15956_ (.A(_05316_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__nand2_2 _15957_ (.A(_05115_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_1 _15958_ (.A(_05019_),
    .B(_03116_),
    .Y(_05326_));
 sky130_fd_sc_hd__xor2_1 _15959_ (.A(_03344_),
    .B(_05326_),
    .X(_05327_));
 sky130_fd_sc_hd__mux2_2 _15960_ (.A0(_05327_),
    .A1(_03247_),
    .S(_05024_),
    .X(_05328_));
 sky130_fd_sc_hd__nand2_4 _15961_ (.A(_05325_),
    .B(_05328_),
    .Y(_05329_));
 sky130_fd_sc_hd__nand3b_4 _15962_ (.A_N(_05328_),
    .B(_05115_),
    .C(_05324_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_4 _15963_ (.A(_05329_),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__buf_6 _15964_ (.A(_05331_),
    .X(_05333_));
 sky130_fd_sc_hd__buf_6 _15965_ (.A(_05333_),
    .X(\div1i.quot[20] ));
 sky130_fd_sc_hd__clkinvlp_2 _15966_ (.A(_05169_),
    .Y(_05334_));
 sky130_fd_sc_hd__nand2_1 _15967_ (.A(_05210_),
    .B(_05314_),
    .Y(_05335_));
 sky130_fd_sc_hd__nand3_2 _15968_ (.A(_05335_),
    .B(_05157_),
    .C(_05136_),
    .Y(_05336_));
 sky130_fd_sc_hd__inv_2 _15969_ (.A(_05176_),
    .Y(_05337_));
 sky130_fd_sc_hd__nand2_2 _15970_ (.A(_05336_),
    .B(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _15971_ (.A(_05338_),
    .B(_05175_),
    .Y(_05339_));
 sky130_fd_sc_hd__or2_1 _15972_ (.A(_05334_),
    .B(_05339_),
    .X(_05340_));
 sky130_fd_sc_hd__nand2_1 _15973_ (.A(_05339_),
    .B(_05334_),
    .Y(_05341_));
 sky130_fd_sc_hd__nand2_1 _15974_ (.A(_05340_),
    .B(_05341_),
    .Y(_05343_));
 sky130_fd_sc_hd__mux2_1 _15975_ (.A0(_05165_),
    .A1(_05343_),
    .S(_05333_),
    .X(_05344_));
 sky130_fd_sc_hd__or2_1 _15976_ (.A(_08527_),
    .B(_05344_),
    .X(_05345_));
 sky130_fd_sc_hd__nand2_1 _15977_ (.A(_05314_),
    .B(_05209_),
    .Y(_05346_));
 sky130_fd_sc_hd__inv_2 _15978_ (.A(_05156_),
    .Y(_05347_));
 sky130_fd_sc_hd__nand2_1 _15979_ (.A(_05346_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__inv_2 _15980_ (.A(_05138_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _15981_ (.A(_05348_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2_1 _15982_ (.A(_05350_),
    .B(_05123_),
    .Y(_05351_));
 sky130_fd_sc_hd__inv_2 _15983_ (.A(_05135_),
    .Y(_05352_));
 sky130_fd_sc_hd__nand2_1 _15984_ (.A(_05351_),
    .B(_05352_),
    .Y(_05354_));
 sky130_fd_sc_hd__nand3_1 _15985_ (.A(_05350_),
    .B(_05135_),
    .C(_05123_),
    .Y(_05355_));
 sky130_fd_sc_hd__nand2_1 _15986_ (.A(_05354_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__nand2_1 _15987_ (.A(_05356_),
    .B(_05288_),
    .Y(_05357_));
 sky130_fd_sc_hd__nand3_1 _15988_ (.A(_05346_),
    .B(_05138_),
    .C(_05347_),
    .Y(_05358_));
 sky130_fd_sc_hd__nand3_1 _15989_ (.A(_05350_),
    .B(net34),
    .C(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__clkinvlp_2 _15990_ (.A(_05359_),
    .Y(_05360_));
 sky130_fd_sc_hd__nand3_1 _15991_ (.A(_05354_),
    .B(net35),
    .C(_05355_),
    .Y(_05361_));
 sky130_fd_sc_hd__nand3_1 _15992_ (.A(_05357_),
    .B(_05360_),
    .C(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_1 _15993_ (.A(_05362_),
    .B(_05361_),
    .Y(_05363_));
 sky130_fd_sc_hd__inv_2 _15994_ (.A(_05208_),
    .Y(_05365_));
 sky130_fd_sc_hd__nand2_1 _15995_ (.A(_05314_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__nand2_1 _15996_ (.A(_05366_),
    .B(_05147_),
    .Y(_05367_));
 sky130_fd_sc_hd__clkinvlp_2 _15997_ (.A(_05205_),
    .Y(_05368_));
 sky130_fd_sc_hd__nand2_1 _15998_ (.A(_05367_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__nand3_1 _15999_ (.A(_05366_),
    .B(_05205_),
    .C(_05147_),
    .Y(_05370_));
 sky130_fd_sc_hd__nand2_1 _16000_ (.A(_05369_),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__nand2_1 _16001_ (.A(_05371_),
    .B(_05310_),
    .Y(_05372_));
 sky130_fd_sc_hd__or2_1 _16002_ (.A(_05365_),
    .B(_05314_),
    .X(_05373_));
 sky130_fd_sc_hd__nand2_1 _16003_ (.A(_05373_),
    .B(_05366_),
    .Y(_05374_));
 sky130_fd_sc_hd__nor2_1 _16004_ (.A(_05321_),
    .B(_05374_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand3_1 _16005_ (.A(_05369_),
    .B(net64),
    .C(_05370_),
    .Y(_05377_));
 sky130_fd_sc_hd__a21boi_2 _16006_ (.A1(_05372_),
    .A2(_05376_),
    .B1_N(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__nand2_1 _16007_ (.A(_05350_),
    .B(_05358_),
    .Y(_05379_));
 sky130_fd_sc_hd__nand2_1 _16008_ (.A(_05379_),
    .B(_05299_),
    .Y(_05380_));
 sky130_fd_sc_hd__nand2_1 _16009_ (.A(_05380_),
    .B(_05359_),
    .Y(_05381_));
 sky130_fd_sc_hd__inv_2 _16010_ (.A(_05381_),
    .Y(_05382_));
 sky130_fd_sc_hd__nand3_1 _16011_ (.A(_05357_),
    .B(_05382_),
    .C(_05361_),
    .Y(_05383_));
 sky130_fd_sc_hd__nor2_1 _16012_ (.A(_05378_),
    .B(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__nor2_1 _16013_ (.A(_05363_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__xor2_1 _16014_ (.A(net63),
    .B(_05374_),
    .X(_05387_));
 sky130_fd_sc_hd__inv_2 _16015_ (.A(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__and2_1 _16016_ (.A(_05372_),
    .B(_05377_),
    .X(_05389_));
 sky130_fd_sc_hd__nand2_1 _16017_ (.A(_05388_),
    .B(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__nor2_1 _16018_ (.A(_05390_),
    .B(_05383_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _16019_ (.A(_05293_),
    .B(_05300_),
    .Y(_05392_));
 sky130_fd_sc_hd__nand2_1 _16020_ (.A(_05392_),
    .B(_05219_),
    .Y(_05393_));
 sky130_fd_sc_hd__nand2_1 _16021_ (.A(_05393_),
    .B(_05304_),
    .Y(_05394_));
 sky130_fd_sc_hd__nand2_1 _16022_ (.A(_05234_),
    .B(_05229_),
    .Y(_05395_));
 sky130_fd_sc_hd__nand3_1 _16023_ (.A(_05392_),
    .B(_05219_),
    .C(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__nand2_1 _16024_ (.A(_05394_),
    .B(_05396_),
    .Y(_05398_));
 sky130_fd_sc_hd__nand2_1 _16025_ (.A(_05398_),
    .B(_05211_),
    .Y(_05399_));
 sky130_fd_sc_hd__nand3_1 _16026_ (.A(_05394_),
    .B(_05738_),
    .C(_05396_),
    .Y(_05400_));
 sky130_fd_sc_hd__nand2_1 _16027_ (.A(_05399_),
    .B(_05400_),
    .Y(_05401_));
 sky130_fd_sc_hd__nand3_1 _16028_ (.A(_05265_),
    .B(_05270_),
    .C(_05274_),
    .Y(_05402_));
 sky130_fd_sc_hd__and2_1 _16029_ (.A(_05402_),
    .B(_05265_),
    .X(_05403_));
 sky130_fd_sc_hd__xor2_2 _16030_ (.A(_05286_),
    .B(_05403_),
    .X(_05404_));
 sky130_fd_sc_hd__nand2_1 _16031_ (.A(_05404_),
    .B(_05178_),
    .Y(_05405_));
 sky130_fd_sc_hd__nand2_1 _16032_ (.A(_05271_),
    .B(_05273_),
    .Y(_05406_));
 sky130_fd_sc_hd__nand2_1 _16033_ (.A(_05406_),
    .B(_05402_),
    .Y(_05407_));
 sky130_fd_sc_hd__nand2_1 _16034_ (.A(_05407_),
    .B(_05189_),
    .Y(_05409_));
 sky130_fd_sc_hd__nand2_1 _16035_ (.A(\div1i.quot[21] ),
    .B(_07308_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand2_1 _16036_ (.A(_05410_),
    .B(_07231_),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_1 _16037_ (.A(_05411_),
    .B(_05273_),
    .Y(_05412_));
 sky130_fd_sc_hd__nand2_1 _16038_ (.A(_05412_),
    .B(_05474_),
    .Y(_05413_));
 sky130_fd_sc_hd__nor2_1 _16039_ (.A(_05189_),
    .B(_05407_),
    .Y(_05414_));
 sky130_fd_sc_hd__a21o_1 _16040_ (.A1(_05409_),
    .A2(_05413_),
    .B1(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__nand2_1 _16041_ (.A(_05405_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__o21ai_1 _16042_ (.A1(_05178_),
    .A2(_05404_),
    .B1(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_1 _16043_ (.A(_05265_),
    .B(_05291_),
    .Y(_05418_));
 sky130_fd_sc_hd__inv_2 _16044_ (.A(_05418_),
    .Y(_05420_));
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(_05402_),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21o_1 _16046_ (.A1(_05421_),
    .A2(_05290_),
    .B1(_05300_),
    .X(_05422_));
 sky130_fd_sc_hd__nand2_1 _16047_ (.A(_05422_),
    .B(_05392_),
    .Y(_05423_));
 sky130_fd_sc_hd__inv_2 _16048_ (.A(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__nand2_1 _16049_ (.A(_05424_),
    .B(net59),
    .Y(_05425_));
 sky130_fd_sc_hd__nand2_1 _16050_ (.A(_05423_),
    .B(_05705_),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_1 _16051_ (.A(_05425_),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__inv_2 _16052_ (.A(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__nand3_1 _16053_ (.A(_05401_),
    .B(_05417_),
    .C(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__nand2_1 _16054_ (.A(_05398_),
    .B(_05738_),
    .Y(_05431_));
 sky130_fd_sc_hd__inv_2 _16055_ (.A(_05425_),
    .Y(_05432_));
 sky130_fd_sc_hd__nand3_1 _16056_ (.A(_05394_),
    .B(_05211_),
    .C(_05396_),
    .Y(_05433_));
 sky130_fd_sc_hd__a21boi_1 _16057_ (.A1(_05431_),
    .A2(_05432_),
    .B1_N(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__nand2_1 _16058_ (.A(_05429_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__nor2_1 _16059_ (.A(_05298_),
    .B(_05395_),
    .Y(_05436_));
 sky130_fd_sc_hd__nand3_1 _16060_ (.A(_05421_),
    .B(_05436_),
    .C(_05290_),
    .Y(_05437_));
 sky130_fd_sc_hd__inv_2 _16061_ (.A(_05235_),
    .Y(_05438_));
 sky130_fd_sc_hd__nand2_1 _16062_ (.A(_05437_),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__nand2_1 _16063_ (.A(_05439_),
    .B(_05306_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand3_1 _16064_ (.A(_05437_),
    .B(_05247_),
    .C(_05438_),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_1 _16065_ (.A(_05440_),
    .B(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__nand2_1 _16066_ (.A(_05443_),
    .B(_05847_),
    .Y(_05444_));
 sky130_fd_sc_hd__nand3_1 _16067_ (.A(_05440_),
    .B(net61),
    .C(_05442_),
    .Y(_05445_));
 sky130_fd_sc_hd__nand2_1 _16068_ (.A(_05444_),
    .B(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__nand2_1 _16069_ (.A(_05440_),
    .B(_05241_),
    .Y(_05447_));
 sky130_fd_sc_hd__nand2_1 _16070_ (.A(_05447_),
    .B(_05309_),
    .Y(_05448_));
 sky130_fd_sc_hd__nand3_1 _16071_ (.A(_05440_),
    .B(_05241_),
    .C(_05256_),
    .Y(_05449_));
 sky130_fd_sc_hd__nand2_1 _16072_ (.A(_05448_),
    .B(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__nand2_1 _16073_ (.A(_05450_),
    .B(_05255_),
    .Y(_05451_));
 sky130_fd_sc_hd__nand3_1 _16074_ (.A(_05448_),
    .B(net62),
    .C(_05449_),
    .Y(_05453_));
 sky130_fd_sc_hd__nand3b_1 _16075_ (.A_N(_05446_),
    .B(_05451_),
    .C(_05453_),
    .Y(_05454_));
 sky130_fd_sc_hd__inv_2 _16076_ (.A(_05454_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand2_1 _16077_ (.A(_05435_),
    .B(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__inv_2 _16078_ (.A(_05445_),
    .Y(_05457_));
 sky130_fd_sc_hd__a21boi_1 _16079_ (.A1(_05451_),
    .A2(_05457_),
    .B1_N(_05453_),
    .Y(_05458_));
 sky130_fd_sc_hd__nand2_1 _16080_ (.A(_05456_),
    .B(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(_05391_),
    .B(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__nand2_1 _16082_ (.A(_05385_),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__nand2_1 _16083_ (.A(_05343_),
    .B(_06045_),
    .Y(_05462_));
 sky130_fd_sc_hd__nand3_1 _16084_ (.A(_05340_),
    .B(net37),
    .C(_05341_),
    .Y(_05464_));
 sky130_fd_sc_hd__or2_1 _16085_ (.A(_05337_),
    .B(_05336_),
    .X(_05465_));
 sky130_fd_sc_hd__nand2_1 _16086_ (.A(_05465_),
    .B(_05338_),
    .Y(_05466_));
 sky130_fd_sc_hd__nand2_1 _16087_ (.A(_05466_),
    .B(_06012_),
    .Y(_05467_));
 sky130_fd_sc_hd__nand3_1 _16088_ (.A(_05465_),
    .B(net36),
    .C(_05338_),
    .Y(_05468_));
 sky130_fd_sc_hd__nand2_1 _16089_ (.A(_05467_),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__inv_2 _16090_ (.A(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__nand3_1 _16091_ (.A(_05462_),
    .B(_05464_),
    .C(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hd__inv_2 _16092_ (.A(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__nand2_1 _16093_ (.A(_05461_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__inv_2 _16094_ (.A(_05468_),
    .Y(_05475_));
 sky130_fd_sc_hd__a21boi_2 _16095_ (.A1(_05462_),
    .A2(_05475_),
    .B1_N(_05464_),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_1 _16096_ (.A(_05473_),
    .B(_05476_),
    .Y(_05477_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(_05336_),
    .B(_05177_),
    .Y(_05478_));
 sky130_fd_sc_hd__inv_2 _16098_ (.A(_05201_),
    .Y(_05479_));
 sky130_fd_sc_hd__nand2_1 _16099_ (.A(_05478_),
    .B(_05479_),
    .Y(_05480_));
 sky130_fd_sc_hd__inv_2 _16100_ (.A(_05186_),
    .Y(_05481_));
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(_05480_),
    .B(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand3_1 _16102_ (.A(_05478_),
    .B(_05186_),
    .C(_05479_),
    .Y(_05483_));
 sky130_fd_sc_hd__nand2_1 _16103_ (.A(_05482_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__inv_2 _16104_ (.A(_05484_),
    .Y(_05486_));
 sky130_fd_sc_hd__nand2_1 _16105_ (.A(_05486_),
    .B(net38),
    .Y(_05487_));
 sky130_fd_sc_hd__nand2_1 _16106_ (.A(_05484_),
    .B(_06155_),
    .Y(_05488_));
 sky130_fd_sc_hd__nand2_1 _16107_ (.A(_05487_),
    .B(_05488_),
    .Y(_05489_));
 sky130_fd_sc_hd__inv_2 _16108_ (.A(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(_05477_),
    .B(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__inv_6 _16110_ (.A(_05333_),
    .Y(_05492_));
 sky130_fd_sc_hd__buf_6 _16111_ (.A(_05492_),
    .X(_05493_));
 sky130_fd_sc_hd__nand3_1 _16112_ (.A(_05473_),
    .B(_05489_),
    .C(_05476_),
    .Y(_05494_));
 sky130_fd_sc_hd__nand3_1 _16113_ (.A(_05491_),
    .B(_05493_),
    .C(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__nand2_1 _16114_ (.A(\div1i.quot[20] ),
    .B(_05486_),
    .Y(_05497_));
 sky130_fd_sc_hd__nand3_1 _16115_ (.A(_05495_),
    .B(net137),
    .C(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__inv_2 _16116_ (.A(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__nand2_1 _16117_ (.A(_05495_),
    .B(_05497_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_1 _16118_ (.A(_05500_),
    .B(net121),
    .Y(_05501_));
 sky130_fd_sc_hd__o21ai_1 _16119_ (.A1(_05345_),
    .A2(_05499_),
    .B1(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__nand2_1 _16120_ (.A(_05492_),
    .B(_05132_),
    .Y(_05503_));
 sky130_fd_sc_hd__nand2_1 _16121_ (.A(\div1i.quot[20] ),
    .B(_05356_),
    .Y(_05504_));
 sky130_fd_sc_hd__nand2_1 _16122_ (.A(_05503_),
    .B(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__or2_1 _16123_ (.A(_08274_),
    .B(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__nand2_1 _16124_ (.A(_05461_),
    .B(_05470_),
    .Y(_05508_));
 sky130_fd_sc_hd__nand3_1 _16125_ (.A(_05385_),
    .B(_05460_),
    .C(_05469_),
    .Y(_05509_));
 sky130_fd_sc_hd__nand3_1 _16126_ (.A(_05508_),
    .B(_05492_),
    .C(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__or2_1 _16127_ (.A(_05466_),
    .B(_05492_),
    .X(_05511_));
 sky130_fd_sc_hd__nand3_1 _16128_ (.A(_05510_),
    .B(_08406_),
    .C(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__inv_2 _16129_ (.A(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hd__nand2_1 _16130_ (.A(_05510_),
    .B(_05511_),
    .Y(_05514_));
 sky130_fd_sc_hd__nand2_1 _16131_ (.A(_05514_),
    .B(_08384_),
    .Y(_05515_));
 sky130_fd_sc_hd__o21a_1 _16132_ (.A1(_05506_),
    .A2(_05513_),
    .B1(_05515_),
    .X(_05516_));
 sky130_fd_sc_hd__nand2_1 _16133_ (.A(_05344_),
    .B(_08527_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_1 _16134_ (.A(_05345_),
    .B(_05517_),
    .Y(_05519_));
 sky130_fd_sc_hd__inv_2 _16135_ (.A(_05519_),
    .Y(_05520_));
 sky130_fd_sc_hd__nand3_1 _16136_ (.A(_05501_),
    .B(_05498_),
    .C(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__nor2_1 _16137_ (.A(_05516_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nor2_1 _16138_ (.A(_05502_),
    .B(_05522_),
    .Y(_05523_));
 sky130_fd_sc_hd__nand2_1 _16139_ (.A(_05515_),
    .B(_05512_),
    .Y(_05524_));
 sky130_fd_sc_hd__inv_4 _16140_ (.A(_05524_),
    .Y(_05525_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(_05505_),
    .B(_08274_),
    .Y(_05526_));
 sky130_fd_sc_hd__nand2_1 _16142_ (.A(_05506_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__inv_2 _16143_ (.A(_05527_),
    .Y(_05528_));
 sky130_fd_sc_hd__nand2_1 _16144_ (.A(_05525_),
    .B(_05528_),
    .Y(_05530_));
 sky130_fd_sc_hd__nor2_1 _16145_ (.A(_05530_),
    .B(_05521_),
    .Y(_05531_));
 sky130_fd_sc_hd__inv_2 _16146_ (.A(_05407_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand2_1 _16147_ (.A(_05331_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__nand2_1 _16148_ (.A(_05261_),
    .B(_05264_),
    .Y(_05534_));
 sky130_fd_sc_hd__nand3b_1 _16149_ (.A_N(_05534_),
    .B(_05329_),
    .C(_05330_),
    .Y(_05535_));
 sky130_fd_sc_hd__nand2_1 _16150_ (.A(_05533_),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__nand2_1 _16151_ (.A(_05536_),
    .B(_11777_),
    .Y(_05537_));
 sky130_fd_sc_hd__inv_2 _16152_ (.A(_05412_),
    .Y(_05538_));
 sky130_fd_sc_hd__nand2_1 _16153_ (.A(_05331_),
    .B(_05538_),
    .Y(_05539_));
 sky130_fd_sc_hd__inv_2 _16154_ (.A(_05410_),
    .Y(_05541_));
 sky130_fd_sc_hd__nand3_1 _16155_ (.A(_05329_),
    .B(_05330_),
    .C(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__nand2_1 _16156_ (.A(_05539_),
    .B(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand2_2 _16157_ (.A(_05543_),
    .B(_07539_),
    .Y(_05544_));
 sky130_fd_sc_hd__nand2_1 _16158_ (.A(_05537_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__inv_2 _16159_ (.A(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__nand3_1 _16160_ (.A(_05539_),
    .B(_05542_),
    .C(_07560_),
    .Y(_05547_));
 sky130_fd_sc_hd__nand3_2 _16161_ (.A(_05331_),
    .B(_05474_),
    .C(_07308_),
    .Y(_05548_));
 sky130_fd_sc_hd__inv_2 _16162_ (.A(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__nand3_2 _16163_ (.A(_05544_),
    .B(_05547_),
    .C(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__nand2_1 _16164_ (.A(_05546_),
    .B(_05550_),
    .Y(_05552_));
 sky130_fd_sc_hd__or2_1 _16165_ (.A(_11777_),
    .B(_05536_),
    .X(_05553_));
 sky130_fd_sc_hd__nand2_1 _16166_ (.A(_05552_),
    .B(_05553_),
    .Y(_05554_));
 sky130_fd_sc_hd__inv_2 _16167_ (.A(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__nand2_1 _16168_ (.A(_05333_),
    .B(_05398_),
    .Y(_05556_));
 sky130_fd_sc_hd__nand3_1 _16169_ (.A(_05329_),
    .B(_05330_),
    .C(_05301_),
    .Y(_05557_));
 sky130_fd_sc_hd__nand2_1 _16170_ (.A(_05556_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__nand2_1 _16171_ (.A(_05558_),
    .B(_08066_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand3_2 _16172_ (.A(_05556_),
    .B(_05557_),
    .C(_08055_),
    .Y(_05560_));
 sky130_fd_sc_hd__nand2_1 _16173_ (.A(_05559_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__inv_2 _16174_ (.A(_05561_),
    .Y(_05563_));
 sky130_fd_sc_hd__inv_2 _16175_ (.A(_05443_),
    .Y(_05564_));
 sky130_fd_sc_hd__nand2_1 _16176_ (.A(_05333_),
    .B(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hd__nand2_1 _16177_ (.A(_05242_),
    .B(_05245_),
    .Y(_05566_));
 sky130_fd_sc_hd__nand3_1 _16178_ (.A(_05329_),
    .B(_05330_),
    .C(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__nand2_1 _16179_ (.A(_05565_),
    .B(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand2_1 _16180_ (.A(_05568_),
    .B(_13588_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand3_1 _16181_ (.A(_05565_),
    .B(_05567_),
    .C(_11579_),
    .Y(_05570_));
 sky130_fd_sc_hd__nand2_1 _16182_ (.A(_05569_),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hd__inv_2 _16183_ (.A(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__nand2_1 _16184_ (.A(_05563_),
    .B(_05572_),
    .Y(_05574_));
 sky130_fd_sc_hd__clkinvlp_2 _16185_ (.A(_05404_),
    .Y(_05575_));
 sky130_fd_sc_hd__nand2_1 _16186_ (.A(_05333_),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hd__nand2_1 _16187_ (.A(_05276_),
    .B(_05281_),
    .Y(_05577_));
 sky130_fd_sc_hd__nand3_1 _16188_ (.A(_05329_),
    .B(_05330_),
    .C(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__nand2_1 _16189_ (.A(_05576_),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__nand2_1 _16190_ (.A(_05579_),
    .B(_07725_),
    .Y(_05580_));
 sky130_fd_sc_hd__nand3_1 _16191_ (.A(_05576_),
    .B(_05578_),
    .C(_07703_),
    .Y(_05581_));
 sky130_fd_sc_hd__nand2_1 _16192_ (.A(_05580_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__inv_2 _16193_ (.A(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__nand2_1 _16194_ (.A(_05333_),
    .B(_05424_),
    .Y(_05585_));
 sky130_fd_sc_hd__nand2_1 _16195_ (.A(_05295_),
    .B(_05296_),
    .Y(_05586_));
 sky130_fd_sc_hd__nand3_1 _16196_ (.A(_05329_),
    .B(_05330_),
    .C(_05586_),
    .Y(_05587_));
 sky130_fd_sc_hd__nand2_1 _16197_ (.A(_05585_),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__nand2_1 _16198_ (.A(_05588_),
    .B(_12029_),
    .Y(_05589_));
 sky130_fd_sc_hd__nand3_1 _16199_ (.A(_05585_),
    .B(_05587_),
    .C(_12051_),
    .Y(_05590_));
 sky130_fd_sc_hd__nand2_1 _16200_ (.A(_05589_),
    .B(_05590_),
    .Y(_05591_));
 sky130_fd_sc_hd__inv_2 _16201_ (.A(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand2_1 _16202_ (.A(_05583_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__nor2_1 _16203_ (.A(_05574_),
    .B(_05593_),
    .Y(_05594_));
 sky130_fd_sc_hd__nand2_1 _16204_ (.A(_05555_),
    .B(_05594_),
    .Y(_05596_));
 sky130_fd_sc_hd__inv_2 _16205_ (.A(_05590_),
    .Y(_05597_));
 sky130_fd_sc_hd__o21ai_1 _16206_ (.A1(_05580_),
    .A2(_05597_),
    .B1(_05589_),
    .Y(_05598_));
 sky130_fd_sc_hd__nor2_1 _16207_ (.A(_05561_),
    .B(_05571_),
    .Y(_05599_));
 sky130_fd_sc_hd__clkinvlp_2 _16208_ (.A(_05570_),
    .Y(_05600_));
 sky130_fd_sc_hd__o21ai_1 _16209_ (.A1(_05560_),
    .A2(_05600_),
    .B1(_05569_),
    .Y(_05601_));
 sky130_fd_sc_hd__a21oi_1 _16210_ (.A1(_05598_),
    .A2(_05599_),
    .B1(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__nand2_2 _16211_ (.A(_05596_),
    .B(_05602_),
    .Y(_05603_));
 sky130_fd_sc_hd__inv_2 _16212_ (.A(_05390_),
    .Y(_05604_));
 sky130_fd_sc_hd__nand2_1 _16213_ (.A(_05459_),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _16214_ (.A(_05605_),
    .B(_05378_),
    .Y(_05607_));
 sky130_fd_sc_hd__nand2_1 _16215_ (.A(_05607_),
    .B(_05382_),
    .Y(_05608_));
 sky130_fd_sc_hd__nand3_1 _16216_ (.A(_05605_),
    .B(_05381_),
    .C(_05378_),
    .Y(_05609_));
 sky130_fd_sc_hd__nand3_1 _16217_ (.A(_05608_),
    .B(_05492_),
    .C(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__or2_1 _16218_ (.A(_05379_),
    .B(_05492_),
    .X(_05611_));
 sky130_fd_sc_hd__nand2_1 _16219_ (.A(_05610_),
    .B(_05611_),
    .Y(_05612_));
 sky130_fd_sc_hd__nand2_1 _16220_ (.A(_05612_),
    .B(_08966_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand3_1 _16221_ (.A(_05610_),
    .B(_08944_),
    .C(_05611_),
    .Y(_05614_));
 sky130_fd_sc_hd__nand2_1 _16222_ (.A(_05333_),
    .B(_05371_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_1 _16223_ (.A1(_05154_),
    .A2(_05333_),
    .B1(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__or2_1 _16224_ (.A(_09054_),
    .B(_05616_),
    .X(_05618_));
 sky130_fd_sc_hd__nand2_1 _16225_ (.A(_05616_),
    .B(_09054_),
    .Y(_05619_));
 sky130_fd_sc_hd__nand2_1 _16226_ (.A(_05618_),
    .B(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__inv_2 _16227_ (.A(_05620_),
    .Y(_05621_));
 sky130_fd_sc_hd__nand3_1 _16228_ (.A(_05613_),
    .B(_05614_),
    .C(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__clkinvlp_2 _16229_ (.A(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hd__or2_1 _16230_ (.A(_05206_),
    .B(\div1i.quot[20] ),
    .X(_05624_));
 sky130_fd_sc_hd__or2b_1 _16231_ (.A(_05374_),
    .B_N(_05333_),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _16232_ (.A(_05624_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand2_1 _16233_ (.A(_05626_),
    .B(_11140_),
    .Y(_05627_));
 sky130_fd_sc_hd__nand3_1 _16234_ (.A(_05624_),
    .B(_05625_),
    .C(_08746_),
    .Y(_05629_));
 sky130_fd_sc_hd__nand2_2 _16235_ (.A(_05627_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_1 _16236_ (.A(_05492_),
    .B(_05252_),
    .Y(_05631_));
 sky130_fd_sc_hd__nand2_1 _16237_ (.A(\div1i.quot[20] ),
    .B(_05450_),
    .Y(_05632_));
 sky130_fd_sc_hd__nand2_1 _16238_ (.A(_05631_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__or2_1 _16239_ (.A(_12260_),
    .B(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__nand2_1 _16240_ (.A(_05633_),
    .B(_12260_),
    .Y(_05635_));
 sky130_fd_sc_hd__nand2_1 _16241_ (.A(_05634_),
    .B(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hd__nor2_1 _16242_ (.A(_05630_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__nand3_1 _16243_ (.A(_05603_),
    .B(_05623_),
    .C(_05637_),
    .Y(_05638_));
 sky130_fd_sc_hd__inv_2 _16244_ (.A(_05614_),
    .Y(_05640_));
 sky130_fd_sc_hd__o21ai_1 _16245_ (.A1(_05618_),
    .A2(_05640_),
    .B1(_05613_),
    .Y(_05641_));
 sky130_fd_sc_hd__o21a_1 _16246_ (.A1(_05634_),
    .A2(_05630_),
    .B1(_05627_),
    .X(_05642_));
 sky130_fd_sc_hd__nor2_1 _16247_ (.A(_05642_),
    .B(_05622_),
    .Y(_05643_));
 sky130_fd_sc_hd__nor2_1 _16248_ (.A(_05641_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__nand2_2 _16249_ (.A(_05644_),
    .B(_05638_),
    .Y(_05645_));
 sky130_fd_sc_hd__nand2_1 _16250_ (.A(_05531_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__nand2_2 _16251_ (.A(_05523_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_1 _16252_ (.A(_05317_),
    .B(_05078_),
    .Y(_05648_));
 sky130_fd_sc_hd__inv_2 _16253_ (.A(_05316_),
    .Y(_05649_));
 sky130_fd_sc_hd__or2_1 _16254_ (.A(_05648_),
    .B(_05649_),
    .X(_05651_));
 sky130_fd_sc_hd__nand2_1 _16255_ (.A(_05649_),
    .B(_05648_),
    .Y(_05652_));
 sky130_fd_sc_hd__nand2_1 _16256_ (.A(_05651_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__inv_2 _16257_ (.A(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_1 _16258_ (.A(_05654_),
    .B(net40),
    .Y(_05655_));
 sky130_fd_sc_hd__nand2_1 _16259_ (.A(_05653_),
    .B(_05408_),
    .Y(_05656_));
 sky130_fd_sc_hd__nand2_1 _16260_ (.A(_05655_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__inv_2 _16261_ (.A(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hd__nand2_1 _16262_ (.A(_05482_),
    .B(_05185_),
    .Y(_05659_));
 sky130_fd_sc_hd__inv_2 _16263_ (.A(_05195_),
    .Y(_05660_));
 sky130_fd_sc_hd__nand2_1 _16264_ (.A(_05659_),
    .B(_05660_),
    .Y(_05662_));
 sky130_fd_sc_hd__nand3_1 _16265_ (.A(_05482_),
    .B(_05195_),
    .C(_05185_),
    .Y(_05663_));
 sky130_fd_sc_hd__nand2_1 _16266_ (.A(_05662_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__nand2_1 _16267_ (.A(_05664_),
    .B(_05375_),
    .Y(_05665_));
 sky130_fd_sc_hd__nand3_1 _16268_ (.A(_05662_),
    .B(net39),
    .C(_05663_),
    .Y(_05666_));
 sky130_fd_sc_hd__nand3_1 _16269_ (.A(_05490_),
    .B(_05665_),
    .C(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hd__nor2_1 _16270_ (.A(_05476_),
    .B(_05667_),
    .Y(_05668_));
 sky130_fd_sc_hd__nand2_1 _16271_ (.A(_05665_),
    .B(_05666_),
    .Y(_05669_));
 sky130_fd_sc_hd__o21ai_1 _16272_ (.A1(_05487_),
    .A2(_05669_),
    .B1(_05666_),
    .Y(_05670_));
 sky130_fd_sc_hd__nor2_1 _16273_ (.A(_05668_),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__nand3b_1 _16274_ (.A_N(_05667_),
    .B(_05461_),
    .C(_05472_),
    .Y(_05673_));
 sky130_fd_sc_hd__nand2_2 _16275_ (.A(_05671_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__or2_1 _16276_ (.A(_05658_),
    .B(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__nand2_1 _16277_ (.A(_05674_),
    .B(_05658_),
    .Y(_05676_));
 sky130_fd_sc_hd__nand3_1 _16278_ (.A(_05675_),
    .B(_05493_),
    .C(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hd__nand2_1 _16279_ (.A(_05654_),
    .B(\div1i.quot[20] ),
    .Y(_05678_));
 sky130_fd_sc_hd__nand2_1 _16280_ (.A(_05677_),
    .B(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__nand2_1 _16281_ (.A(_05679_),
    .B(_09383_),
    .Y(_05680_));
 sky130_fd_sc_hd__nand3_1 _16282_ (.A(_05677_),
    .B(_09361_),
    .C(_05678_),
    .Y(_05681_));
 sky130_fd_sc_hd__mux2_1 _16283_ (.A0(_05192_),
    .A1(_05664_),
    .S(\div1i.quot[20] ),
    .X(_05682_));
 sky130_fd_sc_hd__or2_1 _16284_ (.A(_09548_),
    .B(_05682_),
    .X(_05684_));
 sky130_fd_sc_hd__nand2_1 _16285_ (.A(_05682_),
    .B(_09548_),
    .Y(_05685_));
 sky130_fd_sc_hd__nand2_1 _16286_ (.A(_05684_),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__inv_4 _16287_ (.A(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hd__nand3_1 _16288_ (.A(_05680_),
    .B(_05681_),
    .C(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hd__inv_2 _16289_ (.A(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__nand2_1 _16290_ (.A(_05647_),
    .B(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__inv_2 _16291_ (.A(_05681_),
    .Y(_05691_));
 sky130_fd_sc_hd__o21a_1 _16292_ (.A1(_05684_),
    .A2(_05691_),
    .B1(_05680_),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _16293_ (.A(_05690_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__nand2_1 _16294_ (.A(_05651_),
    .B(_05078_),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_1 _16295_ (.A(_05695_),
    .B(_05318_),
    .Y(_05696_));
 sky130_fd_sc_hd__nand3_1 _16296_ (.A(_05651_),
    .B(_05087_),
    .C(_05078_),
    .Y(_05697_));
 sky130_fd_sc_hd__nand2_1 _16297_ (.A(_05696_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__nand2_1 _16298_ (.A(_05698_),
    .B(_06814_),
    .Y(_05699_));
 sky130_fd_sc_hd__nand3_1 _16299_ (.A(_05696_),
    .B(net41),
    .C(_05697_),
    .Y(_05700_));
 sky130_fd_sc_hd__nand3_1 _16300_ (.A(_05658_),
    .B(_05699_),
    .C(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__inv_2 _16301_ (.A(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hd__nand2_1 _16302_ (.A(_05674_),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__inv_2 _16303_ (.A(_05655_),
    .Y(_05704_));
 sky130_fd_sc_hd__a21boi_2 _16304_ (.A1(_05699_),
    .A2(_05704_),
    .B1_N(_05700_),
    .Y(_05706_));
 sky130_fd_sc_hd__nand2_1 _16305_ (.A(_05703_),
    .B(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hd__inv_2 _16306_ (.A(_05097_),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_1 _16307_ (.A(_05316_),
    .B(_05320_),
    .Y(_05709_));
 sky130_fd_sc_hd__inv_2 _16308_ (.A(_05088_),
    .Y(_05710_));
 sky130_fd_sc_hd__nand2_1 _16309_ (.A(_05709_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__or2_1 _16310_ (.A(_05708_),
    .B(_05711_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_1 _16311_ (.A(_05711_),
    .B(_05708_),
    .Y(_05713_));
 sky130_fd_sc_hd__nand2_1 _16312_ (.A(_05712_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__nand2_1 _16313_ (.A(_05714_),
    .B(_06737_),
    .Y(_05715_));
 sky130_fd_sc_hd__nand3_1 _16314_ (.A(_05712_),
    .B(_06726_),
    .C(_05713_),
    .Y(_05717_));
 sky130_fd_sc_hd__nand2_1 _16315_ (.A(_05715_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__inv_2 _16316_ (.A(_05718_),
    .Y(_05719_));
 sky130_fd_sc_hd__nand2_1 _16317_ (.A(_05707_),
    .B(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__nand3_1 _16318_ (.A(_05703_),
    .B(_05718_),
    .C(_05706_),
    .Y(_05721_));
 sky130_fd_sc_hd__nand3_1 _16319_ (.A(_05720_),
    .B(_05493_),
    .C(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__or2_1 _16320_ (.A(_05493_),
    .B(_05714_),
    .X(_05723_));
 sky130_fd_sc_hd__nand2_1 _16321_ (.A(_05722_),
    .B(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__nand2_1 _16322_ (.A(_05724_),
    .B(_10009_),
    .Y(_05725_));
 sky130_fd_sc_hd__nand3_1 _16323_ (.A(_05722_),
    .B(_09987_),
    .C(_05723_),
    .Y(_05726_));
 sky130_fd_sc_hd__mux2_1 _16324_ (.A0(_05084_),
    .A1(_05698_),
    .S(\div1i.quot[20] ),
    .X(_05728_));
 sky130_fd_sc_hd__inv_2 _16325_ (.A(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__nand2_1 _16326_ (.A(_05729_),
    .B(net120),
    .Y(_05730_));
 sky130_fd_sc_hd__nand2_1 _16327_ (.A(_05728_),
    .B(_09735_),
    .Y(_05731_));
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(_05730_),
    .B(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__inv_2 _16329_ (.A(_05732_),
    .Y(_05733_));
 sky130_fd_sc_hd__nand3_1 _16330_ (.A(_05725_),
    .B(_05726_),
    .C(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__inv_2 _16331_ (.A(_05734_),
    .Y(_05735_));
 sky130_fd_sc_hd__nand2_1 _16332_ (.A(_05693_),
    .B(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand2_1 _16333_ (.A(_05725_),
    .B(_05726_),
    .Y(_05737_));
 sky130_fd_sc_hd__o21a_1 _16334_ (.A1(_05730_),
    .A2(_05737_),
    .B1(_05725_),
    .X(_05739_));
 sky130_fd_sc_hd__nand2_2 _16335_ (.A(_05736_),
    .B(_05739_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2_1 _16336_ (.A(_05713_),
    .B(_05096_),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2b_1 _16337_ (.A_N(_05741_),
    .B(_05104_),
    .Y(_05742_));
 sky130_fd_sc_hd__a21o_1 _16338_ (.A1(_05713_),
    .A2(_05096_),
    .B1(_05104_),
    .X(_05743_));
 sky130_fd_sc_hd__nand2_1 _16339_ (.A(_05742_),
    .B(_05743_),
    .Y(_05744_));
 sky130_fd_sc_hd__mux2_1 _16340_ (.A0(_05744_),
    .A1(_05101_),
    .S(_05493_),
    .X(_05745_));
 sky130_fd_sc_hd__or2_1 _16341_ (.A(_10251_),
    .B(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__nand2_1 _16342_ (.A(_05745_),
    .B(_10251_),
    .Y(_05747_));
 sky130_fd_sc_hd__nand2_1 _16343_ (.A(_05746_),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand2_1 _16344_ (.A(_05051_),
    .B(_05061_),
    .Y(_05750_));
 sky130_fd_sc_hd__inv_4 _16345_ (.A(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__a31o_1 _16346_ (.A1(_05316_),
    .A2(_05105_),
    .A3(_05320_),
    .B1(_05109_),
    .X(_05752_));
 sky130_fd_sc_hd__or2_1 _16347_ (.A(_05751_),
    .B(_05752_),
    .X(_05753_));
 sky130_fd_sc_hd__nand2_1 _16348_ (.A(_05752_),
    .B(_05751_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2_1 _16349_ (.A(_05753_),
    .B(_05754_),
    .Y(_05755_));
 sky130_fd_sc_hd__mux2_1 _16350_ (.A0(_05755_),
    .A1(_05050_),
    .S(_05493_),
    .X(_05756_));
 sky130_fd_sc_hd__or2_1 _16351_ (.A(_10481_),
    .B(_05756_),
    .X(_05757_));
 sky130_fd_sc_hd__nand2_1 _16352_ (.A(_05756_),
    .B(_10481_),
    .Y(_05758_));
 sky130_fd_sc_hd__nand2_1 _16353_ (.A(_05757_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__nor2_1 _16354_ (.A(_05748_),
    .B(_05759_),
    .Y(_05761_));
 sky130_fd_sc_hd__clkinvlp_2 _16355_ (.A(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand2_1 _16356_ (.A(_05744_),
    .B(_06704_),
    .Y(_05763_));
 sky130_fd_sc_hd__clkinvlp_2 _16357_ (.A(_05717_),
    .Y(_05764_));
 sky130_fd_sc_hd__nand3_1 _16358_ (.A(_05742_),
    .B(_05743_),
    .C(net43),
    .Y(_05765_));
 sky130_fd_sc_hd__inv_2 _16359_ (.A(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__a21o_1 _16360_ (.A1(_05763_),
    .A2(_05764_),
    .B1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__nand3_1 _16361_ (.A(_05763_),
    .B(_05719_),
    .C(_05765_),
    .Y(_05768_));
 sky130_fd_sc_hd__nor2_1 _16362_ (.A(_05706_),
    .B(_05768_),
    .Y(_05769_));
 sky130_fd_sc_hd__nor2_1 _16363_ (.A(_05767_),
    .B(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__nor2_1 _16364_ (.A(_05701_),
    .B(_05768_),
    .Y(_05772_));
 sky130_fd_sc_hd__nand2_1 _16365_ (.A(_05674_),
    .B(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__nand2_1 _16366_ (.A(_05770_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__nand2_1 _16367_ (.A(_05754_),
    .B(_05051_),
    .Y(_05775_));
 sky130_fd_sc_hd__xor2_2 _16368_ (.A(_05059_),
    .B(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__inv_2 _16369_ (.A(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__nand2_1 _16370_ (.A(_05777_),
    .B(net46),
    .Y(_05778_));
 sky130_fd_sc_hd__nand2_1 _16371_ (.A(_05776_),
    .B(_06550_),
    .Y(_05779_));
 sky130_fd_sc_hd__nand2_1 _16372_ (.A(_05755_),
    .B(_10426_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand3_1 _16373_ (.A(_05753_),
    .B(_06649_),
    .C(_05754_),
    .Y(_05781_));
 sky130_fd_sc_hd__nand2_1 _16374_ (.A(_05780_),
    .B(_05781_),
    .Y(_05783_));
 sky130_fd_sc_hd__inv_2 _16375_ (.A(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__nand3_1 _16376_ (.A(_05778_),
    .B(_05779_),
    .C(_05784_),
    .Y(_05785_));
 sky130_fd_sc_hd__inv_2 _16377_ (.A(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__nand2_1 _16378_ (.A(_05774_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__inv_2 _16379_ (.A(_05779_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21a_1 _16380_ (.A1(_05781_),
    .A2(_05788_),
    .B1(_05778_),
    .X(_05789_));
 sky130_fd_sc_hd__nand2_1 _16381_ (.A(_05787_),
    .B(_05789_),
    .Y(_05790_));
 sky130_fd_sc_hd__inv_2 _16382_ (.A(_05042_),
    .Y(_05791_));
 sky130_fd_sc_hd__a21o_1 _16383_ (.A1(_05752_),
    .A2(_05063_),
    .B1(_05110_),
    .X(_05792_));
 sky130_fd_sc_hd__or2_1 _16384_ (.A(_05791_),
    .B(_05792_),
    .X(_05794_));
 sky130_fd_sc_hd__nand2_1 _16385_ (.A(_05792_),
    .B(_05791_),
    .Y(_05795_));
 sky130_fd_sc_hd__nand2_1 _16386_ (.A(_05794_),
    .B(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hd__inv_2 _16387_ (.A(_05796_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand2_1 _16388_ (.A(_05797_),
    .B(net47),
    .Y(_05798_));
 sky130_fd_sc_hd__nand2_1 _16389_ (.A(_05796_),
    .B(_06594_),
    .Y(_05799_));
 sky130_fd_sc_hd__nand2_1 _16390_ (.A(_05798_),
    .B(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__inv_2 _16391_ (.A(_05800_),
    .Y(_05801_));
 sky130_fd_sc_hd__nand2_1 _16392_ (.A(_05790_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__nand3_1 _16393_ (.A(_05787_),
    .B(_05789_),
    .C(_05800_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand3_1 _16394_ (.A(_05802_),
    .B(_05493_),
    .C(_05803_),
    .Y(_05805_));
 sky130_fd_sc_hd__nand2_1 _16395_ (.A(_05797_),
    .B(\div1i.quot[20] ),
    .Y(_05806_));
 sky130_fd_sc_hd__nand2_1 _16396_ (.A(_05805_),
    .B(_05806_),
    .Y(_05807_));
 sky130_fd_sc_hd__nand2_1 _16397_ (.A(_05807_),
    .B(_10887_),
    .Y(_05808_));
 sky130_fd_sc_hd__nand3_2 _16398_ (.A(_05805_),
    .B(_10909_),
    .C(_05806_),
    .Y(_05809_));
 sky130_fd_sc_hd__mux2_1 _16399_ (.A0(_05776_),
    .A1(_05056_),
    .S(_05493_),
    .X(_05810_));
 sky130_fd_sc_hd__or2_1 _16400_ (.A(_10701_),
    .B(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__nand2_1 _16401_ (.A(_05810_),
    .B(_10701_),
    .Y(_05812_));
 sky130_fd_sc_hd__nand2_1 _16402_ (.A(_05811_),
    .B(_05812_),
    .Y(_05813_));
 sky130_fd_sc_hd__inv_2 _16403_ (.A(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__nand3_1 _16404_ (.A(_05808_),
    .B(_05809_),
    .C(_05814_),
    .Y(_05816_));
 sky130_fd_sc_hd__nor2_1 _16405_ (.A(_05762_),
    .B(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__nand2_4 _16406_ (.A(_05740_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__inv_2 _16407_ (.A(_05809_),
    .Y(_05819_));
 sky130_fd_sc_hd__o21ai_1 _16408_ (.A1(_05811_),
    .A2(_05819_),
    .B1(_05808_),
    .Y(_05820_));
 sky130_fd_sc_hd__o21a_1 _16409_ (.A1(_05746_),
    .A2(_05759_),
    .B1(_05757_),
    .X(_05821_));
 sky130_fd_sc_hd__nor2_1 _16410_ (.A(_05821_),
    .B(_05816_),
    .Y(_05822_));
 sky130_fd_sc_hd__nor2_2 _16411_ (.A(_05820_),
    .B(_05822_),
    .Y(_05823_));
 sky130_fd_sc_hd__nand2_4 _16412_ (.A(_05818_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__nand2_2 _16413_ (.A(_05795_),
    .B(_05041_),
    .Y(_05825_));
 sky130_fd_sc_hd__xor2_4 _16414_ (.A(_05029_),
    .B(_05825_),
    .X(_05827_));
 sky130_fd_sc_hd__nand3_2 _16415_ (.A(_05802_),
    .B(_05493_),
    .C(_05798_),
    .Y(_05828_));
 sky130_fd_sc_hd__xor2_4 _16416_ (.A(_05827_),
    .B(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__inv_2 _16417_ (.A(_05829_),
    .Y(_05830_));
 sky130_fd_sc_hd__nand2_8 _16418_ (.A(_05824_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand3_4 _16419_ (.A(_05818_),
    .B(_05823_),
    .C(_05829_),
    .Y(_05832_));
 sky130_fd_sc_hd__nand2_8 _16420_ (.A(_05832_),
    .B(_05831_),
    .Y(_05833_));
 sky130_fd_sc_hd__buf_8 _16421_ (.A(_05833_),
    .X(_05834_));
 sky130_fd_sc_hd__buf_12 _16422_ (.A(net235),
    .X(\div1i.quot[19] ));
 sky130_fd_sc_hd__inv_2 _16423_ (.A(_05636_),
    .Y(_05835_));
 sky130_fd_sc_hd__or2_1 _16424_ (.A(_05835_),
    .B(_05603_),
    .X(_05837_));
 sky130_fd_sc_hd__nand2_1 _16425_ (.A(_05603_),
    .B(_05835_),
    .Y(_05838_));
 sky130_fd_sc_hd__nand2_1 _16426_ (.A(_05837_),
    .B(_05838_),
    .Y(_05839_));
 sky130_fd_sc_hd__inv_2 _16427_ (.A(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_1 _16428_ (.A(_05840_),
    .B(net63),
    .Y(_05841_));
 sky130_fd_sc_hd__nand2_1 _16429_ (.A(_05839_),
    .B(_05321_),
    .Y(_05842_));
 sky130_fd_sc_hd__nand2_1 _16430_ (.A(_05841_),
    .B(_05842_),
    .Y(_05843_));
 sky130_fd_sc_hd__inv_2 _16431_ (.A(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__nand2_1 _16432_ (.A(_05553_),
    .B(_05537_),
    .Y(_05845_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(_05550_),
    .B(_05544_),
    .Y(_05846_));
 sky130_fd_sc_hd__xor2_1 _16434_ (.A(_05845_),
    .B(_05846_),
    .X(_05848_));
 sky130_fd_sc_hd__nand2_1 _16435_ (.A(_05848_),
    .B(_05178_),
    .Y(_05849_));
 sky130_fd_sc_hd__nand2_1 _16436_ (.A(_05544_),
    .B(_05547_),
    .Y(_05850_));
 sky130_fd_sc_hd__nand2_1 _16437_ (.A(_05850_),
    .B(_05548_),
    .Y(_05851_));
 sky130_fd_sc_hd__nand2_1 _16438_ (.A(_05851_),
    .B(_05550_),
    .Y(_05852_));
 sky130_fd_sc_hd__nand2_1 _16439_ (.A(_05852_),
    .B(_05189_),
    .Y(_05853_));
 sky130_fd_sc_hd__nand3_1 _16440_ (.A(_05851_),
    .B(net55),
    .C(_05550_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_1 _16441_ (.A1(_05496_),
    .A2(\div1i.quot[20] ),
    .B1(_05474_),
    .Y(_05855_));
 sky130_fd_sc_hd__nand3_1 _16442_ (.A(_05853_),
    .B(_05854_),
    .C(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(_05856_),
    .B(_05854_),
    .Y(_05857_));
 sky130_fd_sc_hd__nand2_1 _16444_ (.A(_05849_),
    .B(_05857_),
    .Y(_05859_));
 sky130_fd_sc_hd__inv_2 _16445_ (.A(_05848_),
    .Y(_05860_));
 sky130_fd_sc_hd__nand2_1 _16446_ (.A(_05860_),
    .B(net58),
    .Y(_05861_));
 sky130_fd_sc_hd__nand2_1 _16447_ (.A(_05859_),
    .B(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__nand2_1 _16448_ (.A(_05554_),
    .B(_05582_),
    .Y(_05863_));
 sky130_fd_sc_hd__nand3_1 _16449_ (.A(_05552_),
    .B(_05553_),
    .C(_05583_),
    .Y(_05864_));
 sky130_fd_sc_hd__nand2_1 _16450_ (.A(_05863_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__nand2_1 _16451_ (.A(_05865_),
    .B(_05705_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand3_1 _16452_ (.A(_05863_),
    .B(net59),
    .C(_05864_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand2_1 _16453_ (.A(_05866_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__inv_2 _16454_ (.A(_05868_),
    .Y(_05870_));
 sky130_fd_sc_hd__nand2_1 _16455_ (.A(_05862_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__nand2_1 _16456_ (.A(_05871_),
    .B(_05867_),
    .Y(_05872_));
 sky130_fd_sc_hd__nand2_1 _16457_ (.A(_05864_),
    .B(_05580_),
    .Y(_05873_));
 sky130_fd_sc_hd__xor2_2 _16458_ (.A(_05591_),
    .B(_05873_),
    .X(_05874_));
 sky130_fd_sc_hd__nand2_1 _16459_ (.A(_05874_),
    .B(_05738_),
    .Y(_05875_));
 sky130_fd_sc_hd__nand2_1 _16460_ (.A(_05872_),
    .B(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__inv_4 _16461_ (.A(_05874_),
    .Y(_05877_));
 sky130_fd_sc_hd__nand2_1 _16462_ (.A(_05877_),
    .B(_05211_),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_1 _16463_ (.A(_05876_),
    .B(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__or2_1 _16464_ (.A(_05593_),
    .B(_05554_),
    .X(_05881_));
 sky130_fd_sc_hd__inv_2 _16465_ (.A(_05598_),
    .Y(_05882_));
 sky130_fd_sc_hd__nand2_1 _16466_ (.A(_05881_),
    .B(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__nand2_1 _16467_ (.A(_05883_),
    .B(_05563_),
    .Y(_05884_));
 sky130_fd_sc_hd__nand3_1 _16468_ (.A(_05881_),
    .B(_05561_),
    .C(_05882_),
    .Y(_05885_));
 sky130_fd_sc_hd__nand2_1 _16469_ (.A(_05884_),
    .B(_05885_),
    .Y(_05886_));
 sky130_fd_sc_hd__inv_2 _16470_ (.A(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__nand2_1 _16471_ (.A(_05887_),
    .B(net61),
    .Y(_05888_));
 sky130_fd_sc_hd__nand2_1 _16472_ (.A(_05886_),
    .B(_05847_),
    .Y(_05889_));
 sky130_fd_sc_hd__nand2_1 _16473_ (.A(_05888_),
    .B(_05889_),
    .Y(_05890_));
 sky130_fd_sc_hd__inv_2 _16474_ (.A(_05890_),
    .Y(_05892_));
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(_05879_),
    .B(_05892_),
    .Y(_05893_));
 sky130_fd_sc_hd__nand2_1 _16476_ (.A(_05884_),
    .B(_05560_),
    .Y(_05894_));
 sky130_fd_sc_hd__nand2_1 _16477_ (.A(_05894_),
    .B(_05572_),
    .Y(_05895_));
 sky130_fd_sc_hd__buf_6 _16478_ (.A(net62),
    .X(_05896_));
 sky130_fd_sc_hd__nand3_1 _16479_ (.A(_05884_),
    .B(_05560_),
    .C(_05571_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand3_1 _16480_ (.A(_05895_),
    .B(_05896_),
    .C(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__nand2_1 _16481_ (.A(_05898_),
    .B(_05888_),
    .Y(_05899_));
 sky130_fd_sc_hd__inv_2 _16482_ (.A(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__nand2_1 _16483_ (.A(_05895_),
    .B(_05897_),
    .Y(_05901_));
 sky130_fd_sc_hd__nand2_1 _16484_ (.A(_05901_),
    .B(_05255_),
    .Y(_05903_));
 sky130_fd_sc_hd__a21boi_2 _16485_ (.A1(_05893_),
    .A2(_05900_),
    .B1_N(_05903_),
    .Y(_05904_));
 sky130_fd_sc_hd__or2_1 _16486_ (.A(_05844_),
    .B(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__nand2_1 _16487_ (.A(_05904_),
    .B(_05844_),
    .Y(_05906_));
 sky130_fd_sc_hd__nand2_1 _16488_ (.A(_05905_),
    .B(_05906_),
    .Y(_05907_));
 sky130_fd_sc_hd__nand3b_1 _16489_ (.A_N(_05907_),
    .B(_05832_),
    .C(_05831_),
    .Y(_05908_));
 sky130_fd_sc_hd__nand2_1 _16490_ (.A(_05834_),
    .B(_05840_),
    .Y(_05909_));
 sky130_fd_sc_hd__nand2_1 _16491_ (.A(_05908_),
    .B(_05909_),
    .Y(_05910_));
 sky130_fd_sc_hd__nand2_1 _16492_ (.A(_05910_),
    .B(_11140_),
    .Y(_05911_));
 sky130_fd_sc_hd__nand3_1 _16493_ (.A(_05908_),
    .B(_08746_),
    .C(_05909_),
    .Y(_05912_));
 sky130_fd_sc_hd__nand2_4 _16494_ (.A(_05911_),
    .B(_05912_),
    .Y(_05914_));
 sky130_fd_sc_hd__buf_6 _16495_ (.A(_12260_),
    .X(_05915_));
 sky130_fd_sc_hd__inv_6 _16496_ (.A(_05833_),
    .Y(_05916_));
 sky130_fd_sc_hd__nand2_1 _16497_ (.A(_05903_),
    .B(_05898_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand2_1 _16498_ (.A(_05893_),
    .B(_05888_),
    .Y(_05918_));
 sky130_fd_sc_hd__xor2_1 _16499_ (.A(_05917_),
    .B(_05918_),
    .X(_05919_));
 sky130_fd_sc_hd__nand2_1 _16500_ (.A(_05916_),
    .B(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__nand2_1 _16501_ (.A(_05834_),
    .B(_05901_),
    .Y(_05921_));
 sky130_fd_sc_hd__nand2_1 _16502_ (.A(_05920_),
    .B(_05921_),
    .Y(_05922_));
 sky130_fd_sc_hd__or2_4 _16503_ (.A(_05915_),
    .B(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__nand2_1 _16504_ (.A(_05922_),
    .B(_05915_),
    .Y(_05925_));
 sky130_fd_sc_hd__nand2_2 _16505_ (.A(_05923_),
    .B(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__nor2_2 _16506_ (.A(_05914_),
    .B(_05926_),
    .Y(_05927_));
 sky130_fd_sc_hd__inv_2 _16507_ (.A(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__nand2_1 _16508_ (.A(_05603_),
    .B(_05637_),
    .Y(_05929_));
 sky130_fd_sc_hd__nand2_1 _16509_ (.A(_05929_),
    .B(_05642_),
    .Y(_05930_));
 sky130_fd_sc_hd__nand2_1 _16510_ (.A(_05930_),
    .B(_05621_),
    .Y(_05931_));
 sky130_fd_sc_hd__nand3_1 _16511_ (.A(_05929_),
    .B(_05620_),
    .C(_05642_),
    .Y(_05932_));
 sky130_fd_sc_hd__nand2_1 _16512_ (.A(_05931_),
    .B(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__nand2_1 _16513_ (.A(_05933_),
    .B(_05299_),
    .Y(_05934_));
 sky130_fd_sc_hd__nand3_2 _16514_ (.A(_05931_),
    .B(net34),
    .C(_05932_),
    .Y(_05936_));
 sky130_fd_sc_hd__nand2_1 _16515_ (.A(_05934_),
    .B(_05936_),
    .Y(_05937_));
 sky130_fd_sc_hd__inv_4 _16516_ (.A(_05937_),
    .Y(_05938_));
 sky130_fd_sc_hd__inv_2 _16517_ (.A(_05630_),
    .Y(_05939_));
 sky130_fd_sc_hd__nand2_1 _16518_ (.A(_05838_),
    .B(_05634_),
    .Y(_05940_));
 sky130_fd_sc_hd__or2_1 _16519_ (.A(_05939_),
    .B(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__nand2_1 _16520_ (.A(_05940_),
    .B(_05939_),
    .Y(_05942_));
 sky130_fd_sc_hd__nand3_1 _16521_ (.A(_05941_),
    .B(net64),
    .C(_05942_),
    .Y(_05943_));
 sky130_fd_sc_hd__nand2_1 _16522_ (.A(_05941_),
    .B(_05942_),
    .Y(_05944_));
 sky130_fd_sc_hd__nand2_1 _16523_ (.A(_05944_),
    .B(_05310_),
    .Y(_05945_));
 sky130_fd_sc_hd__nand3_1 _16524_ (.A(_05844_),
    .B(_05943_),
    .C(_05945_),
    .Y(_05947_));
 sky130_fd_sc_hd__inv_2 _16525_ (.A(_05947_),
    .Y(_05948_));
 sky130_fd_sc_hd__nand2_1 _16526_ (.A(_05904_),
    .B(_05948_),
    .Y(_05949_));
 sky130_fd_sc_hd__inv_2 _16527_ (.A(_05841_),
    .Y(_05950_));
 sky130_fd_sc_hd__inv_2 _16528_ (.A(_05943_),
    .Y(_05951_));
 sky130_fd_sc_hd__a21oi_1 _16529_ (.A1(_05945_),
    .A2(_05950_),
    .B1(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__nand2_1 _16530_ (.A(_05949_),
    .B(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__or2_1 _16531_ (.A(_05938_),
    .B(_05953_),
    .X(_05954_));
 sky130_fd_sc_hd__inv_2 _16532_ (.A(_05954_),
    .Y(_05955_));
 sky130_fd_sc_hd__nand2_1 _16533_ (.A(_05953_),
    .B(_05938_),
    .Y(_05956_));
 sky130_fd_sc_hd__nand2_1 _16534_ (.A(_05916_),
    .B(_05956_),
    .Y(_05958_));
 sky130_fd_sc_hd__or2_4 _16535_ (.A(_05933_),
    .B(_05916_),
    .X(_05959_));
 sky130_fd_sc_hd__o211ai_1 _16536_ (.A1(_05955_),
    .A2(_05958_),
    .B1(_08944_),
    .C1(_05959_),
    .Y(_05960_));
 sky130_fd_sc_hd__o21ai_2 _16537_ (.A1(_05955_),
    .A2(_05958_),
    .B1(_05959_),
    .Y(_05961_));
 sky130_fd_sc_hd__nand2_2 _16538_ (.A(_05961_),
    .B(_08966_),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_2 _16539_ (.A(_05960_),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__inv_2 _16540_ (.A(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__nand2_1 _16541_ (.A(_05945_),
    .B(_05943_),
    .Y(_05965_));
 sky130_fd_sc_hd__nand2_1 _16542_ (.A(_05906_),
    .B(_05841_),
    .Y(_05966_));
 sky130_fd_sc_hd__xor2_1 _16543_ (.A(_05965_),
    .B(_05966_),
    .X(_05967_));
 sky130_fd_sc_hd__nand2_1 _16544_ (.A(_05967_),
    .B(_05916_),
    .Y(_05969_));
 sky130_fd_sc_hd__nand2_1 _16545_ (.A(net235),
    .B(_05944_),
    .Y(_05970_));
 sky130_fd_sc_hd__nand2_2 _16546_ (.A(_05969_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__xor2_2 _16547_ (.A(_09076_),
    .B(_05971_),
    .X(_05972_));
 sky130_fd_sc_hd__inv_2 _16548_ (.A(_05972_),
    .Y(_05973_));
 sky130_fd_sc_hd__nand2_1 _16549_ (.A(_05964_),
    .B(_05973_),
    .Y(_05974_));
 sky130_fd_sc_hd__nor2_1 _16550_ (.A(_05928_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__inv_2 _16551_ (.A(_05852_),
    .Y(_05976_));
 sky130_fd_sc_hd__nand2_1 _16552_ (.A(_05834_),
    .B(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__a21o_1 _16553_ (.A1(_05853_),
    .A2(_05854_),
    .B1(_05855_),
    .X(_05978_));
 sky130_fd_sc_hd__nand2_1 _16554_ (.A(_05978_),
    .B(_05856_),
    .Y(_05980_));
 sky130_fd_sc_hd__nand3b_1 _16555_ (.A_N(_05980_),
    .B(_05831_),
    .C(_05832_),
    .Y(_05981_));
 sky130_fd_sc_hd__nand2_2 _16556_ (.A(_05977_),
    .B(_05981_),
    .Y(_05982_));
 sky130_fd_sc_hd__buf_4 _16557_ (.A(_11777_),
    .X(_05983_));
 sky130_fd_sc_hd__nand2_2 _16558_ (.A(_05982_),
    .B(_05983_),
    .Y(_05984_));
 sky130_fd_sc_hd__nor2_1 _16559_ (.A(_05496_),
    .B(_05493_),
    .Y(_05985_));
 sky130_fd_sc_hd__or2_1 _16560_ (.A(_07242_),
    .B(_05985_),
    .X(_05986_));
 sky130_fd_sc_hd__nand2_1 _16561_ (.A(_05986_),
    .B(_05548_),
    .Y(_05987_));
 sky130_fd_sc_hd__clkinvlp_2 _16562_ (.A(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand2_2 _16563_ (.A(_05834_),
    .B(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__nand3_1 _16564_ (.A(_05831_),
    .B(_05832_),
    .C(_05985_),
    .Y(_05991_));
 sky130_fd_sc_hd__nand2_2 _16565_ (.A(_05989_),
    .B(_05991_),
    .Y(_05992_));
 sky130_fd_sc_hd__nand2_4 _16566_ (.A(_05992_),
    .B(_07539_),
    .Y(_05993_));
 sky130_fd_sc_hd__nand2_2 _16567_ (.A(_05984_),
    .B(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__inv_2 _16568_ (.A(_05994_),
    .Y(_05995_));
 sky130_fd_sc_hd__nand3_2 _16569_ (.A(_05989_),
    .B(_07560_),
    .C(_05991_),
    .Y(_05996_));
 sky130_fd_sc_hd__nand3_2 _16570_ (.A(_05834_),
    .B(_05474_),
    .C(_07308_),
    .Y(_05997_));
 sky130_fd_sc_hd__inv_2 _16571_ (.A(_05997_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand3_4 _16572_ (.A(_05993_),
    .B(_05996_),
    .C(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__or2_4 _16573_ (.A(_11777_),
    .B(_05982_),
    .X(_06000_));
 sky130_fd_sc_hd__inv_2 _16574_ (.A(_06000_),
    .Y(_06002_));
 sky130_fd_sc_hd__a21oi_1 _16575_ (.A1(_05995_),
    .A2(_05999_),
    .B1(_06002_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand2_1 _16576_ (.A(_05833_),
    .B(_05887_),
    .Y(_06004_));
 sky130_fd_sc_hd__or2_1 _16577_ (.A(_05892_),
    .B(_05879_),
    .X(_06005_));
 sky130_fd_sc_hd__nand2_1 _16578_ (.A(_06005_),
    .B(_05893_),
    .Y(_06006_));
 sky130_fd_sc_hd__inv_2 _16579_ (.A(_06006_),
    .Y(_06007_));
 sky130_fd_sc_hd__nand3_1 _16580_ (.A(_05831_),
    .B(_05832_),
    .C(_06007_),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2_1 _16581_ (.A(_06004_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__nand2_1 _16582_ (.A(_06009_),
    .B(_13588_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand3_1 _16583_ (.A(_06004_),
    .B(_11579_),
    .C(_06008_),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2_2 _16584_ (.A(_06010_),
    .B(_06011_),
    .Y(_06013_));
 sky130_fd_sc_hd__inv_2 _16585_ (.A(_06013_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_1 _16586_ (.A(_05833_),
    .B(_05877_),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2_1 _16587_ (.A(_05878_),
    .B(_05875_),
    .Y(_06016_));
 sky130_fd_sc_hd__xnor2_1 _16588_ (.A(_05872_),
    .B(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand3_1 _16589_ (.A(_05831_),
    .B(_05832_),
    .C(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__nand2_1 _16590_ (.A(_06015_),
    .B(_06018_),
    .Y(_06019_));
 sky130_fd_sc_hd__nand2_2 _16591_ (.A(_06019_),
    .B(_08055_),
    .Y(_06020_));
 sky130_fd_sc_hd__nand3_1 _16592_ (.A(_06015_),
    .B(_08066_),
    .C(_06018_),
    .Y(_06021_));
 sky130_fd_sc_hd__nand2_2 _16593_ (.A(_06020_),
    .B(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__inv_2 _16594_ (.A(_06022_),
    .Y(_06024_));
 sky130_fd_sc_hd__nand2_1 _16595_ (.A(_06014_),
    .B(_06024_),
    .Y(_06025_));
 sky130_fd_sc_hd__inv_2 _16596_ (.A(_05865_),
    .Y(_06026_));
 sky130_fd_sc_hd__nand2_1 _16597_ (.A(_05833_),
    .B(_06026_),
    .Y(_06027_));
 sky130_fd_sc_hd__or2_1 _16598_ (.A(_05870_),
    .B(_05862_),
    .X(_06028_));
 sky130_fd_sc_hd__nand2_1 _16599_ (.A(_06028_),
    .B(_05871_),
    .Y(_06029_));
 sky130_fd_sc_hd__inv_2 _16600_ (.A(_06029_),
    .Y(_06030_));
 sky130_fd_sc_hd__nand3_1 _16601_ (.A(_05831_),
    .B(_05832_),
    .C(_06030_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand2_1 _16602_ (.A(_06027_),
    .B(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__buf_6 _16603_ (.A(_12029_),
    .X(_06033_));
 sky130_fd_sc_hd__nand2_1 _16604_ (.A(_06032_),
    .B(_06033_),
    .Y(_06035_));
 sky130_fd_sc_hd__nand3_1 _16605_ (.A(_06027_),
    .B(_12051_),
    .C(_06031_),
    .Y(_06036_));
 sky130_fd_sc_hd__nand2_2 _16606_ (.A(_06035_),
    .B(_06036_),
    .Y(_06037_));
 sky130_fd_sc_hd__inv_2 _16607_ (.A(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__nand2_1 _16608_ (.A(_05833_),
    .B(_05860_),
    .Y(_06039_));
 sky130_fd_sc_hd__nand2_1 _16609_ (.A(_05861_),
    .B(_05849_),
    .Y(_06040_));
 sky130_fd_sc_hd__xnor2_1 _16610_ (.A(_05857_),
    .B(_06040_),
    .Y(_06041_));
 sky130_fd_sc_hd__nand3_2 _16611_ (.A(_05831_),
    .B(_05832_),
    .C(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__nand2_1 _16612_ (.A(_06039_),
    .B(_06042_),
    .Y(_06043_));
 sky130_fd_sc_hd__nand2_1 _16613_ (.A(_06043_),
    .B(_07725_),
    .Y(_06044_));
 sky130_fd_sc_hd__buf_6 _16614_ (.A(_07703_),
    .X(_06046_));
 sky130_fd_sc_hd__nand3_1 _16615_ (.A(_06039_),
    .B(_06046_),
    .C(_06042_),
    .Y(_06047_));
 sky130_fd_sc_hd__nand2_1 _16616_ (.A(_06044_),
    .B(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__inv_2 _16617_ (.A(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand2_1 _16618_ (.A(_06038_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__nor2_1 _16619_ (.A(_06025_),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__nand2_1 _16620_ (.A(_06003_),
    .B(_06051_),
    .Y(_06052_));
 sky130_fd_sc_hd__inv_2 _16621_ (.A(_06036_),
    .Y(_06053_));
 sky130_fd_sc_hd__o21ai_2 _16622_ (.A1(_06044_),
    .A2(_06053_),
    .B1(_06035_),
    .Y(_06054_));
 sky130_fd_sc_hd__nor2_1 _16623_ (.A(_06013_),
    .B(_06022_),
    .Y(_06055_));
 sky130_fd_sc_hd__inv_2 _16624_ (.A(_06011_),
    .Y(_06057_));
 sky130_fd_sc_hd__o21ai_1 _16625_ (.A1(_06020_),
    .A2(_06057_),
    .B1(_06010_),
    .Y(_06058_));
 sky130_fd_sc_hd__a21oi_1 _16626_ (.A1(_06054_),
    .A2(_06055_),
    .B1(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_2 _16627_ (.A(_06052_),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__nand2_1 _16628_ (.A(_05975_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__nor2_1 _16629_ (.A(_05963_),
    .B(_05972_),
    .Y(_06062_));
 sky130_fd_sc_hd__o21ai_4 _16630_ (.A1(_05914_),
    .A2(_05923_),
    .B1(_05911_),
    .Y(_06063_));
 sky130_fd_sc_hd__or2_4 _16631_ (.A(_09054_),
    .B(_05971_),
    .X(_06064_));
 sky130_fd_sc_hd__nor2_1 _16632_ (.A(_08966_),
    .B(_05961_),
    .Y(_06065_));
 sky130_fd_sc_hd__o21ai_1 _16633_ (.A1(_06064_),
    .A2(_06065_),
    .B1(_05962_),
    .Y(_06066_));
 sky130_fd_sc_hd__a21oi_1 _16634_ (.A1(_06062_),
    .A2(_06063_),
    .B1(_06066_),
    .Y(_06068_));
 sky130_fd_sc_hd__nand2_2 _16635_ (.A(_06068_),
    .B(_06061_),
    .Y(_06069_));
 sky130_fd_sc_hd__nand2_1 _16636_ (.A(_05645_),
    .B(_05528_),
    .Y(_06070_));
 sky130_fd_sc_hd__nand2_1 _16637_ (.A(_06070_),
    .B(_05506_),
    .Y(_06071_));
 sky130_fd_sc_hd__or2_1 _16638_ (.A(_05525_),
    .B(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__nand2_1 _16639_ (.A(_06071_),
    .B(_05525_),
    .Y(_06073_));
 sky130_fd_sc_hd__nand2_1 _16640_ (.A(_06072_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__nand2_2 _16641_ (.A(_06074_),
    .B(_06045_),
    .Y(_06075_));
 sky130_fd_sc_hd__nand3_1 _16642_ (.A(_06072_),
    .B(net37),
    .C(_06073_),
    .Y(_06076_));
 sky130_fd_sc_hd__nand2_1 _16643_ (.A(_06075_),
    .B(_06076_),
    .Y(_06077_));
 sky130_fd_sc_hd__nand2_1 _16644_ (.A(_05931_),
    .B(_05618_),
    .Y(_06079_));
 sky130_fd_sc_hd__nand2_1 _16645_ (.A(_05613_),
    .B(_05614_),
    .Y(_06080_));
 sky130_fd_sc_hd__inv_2 _16646_ (.A(_06080_),
    .Y(_06081_));
 sky130_fd_sc_hd__nand2_1 _16647_ (.A(_06079_),
    .B(_06081_),
    .Y(_06082_));
 sky130_fd_sc_hd__nand3_1 _16648_ (.A(_05931_),
    .B(_06080_),
    .C(_05618_),
    .Y(_06083_));
 sky130_fd_sc_hd__nand2_1 _16649_ (.A(_06082_),
    .B(_06083_),
    .Y(_06084_));
 sky130_fd_sc_hd__nand2_1 _16650_ (.A(_06084_),
    .B(_05288_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand3_2 _16651_ (.A(_06082_),
    .B(net35),
    .C(_06083_),
    .Y(_06086_));
 sky130_fd_sc_hd__nand3_1 _16652_ (.A(_06085_),
    .B(_06086_),
    .C(_05938_),
    .Y(_06087_));
 sky130_fd_sc_hd__inv_2 _16653_ (.A(_06087_),
    .Y(_06088_));
 sky130_fd_sc_hd__nand3_1 _16654_ (.A(_05904_),
    .B(_06088_),
    .C(_05948_),
    .Y(_06090_));
 sky130_fd_sc_hd__inv_2 _16655_ (.A(_05936_),
    .Y(_06091_));
 sky130_fd_sc_hd__inv_2 _16656_ (.A(_06086_),
    .Y(_06092_));
 sky130_fd_sc_hd__a21o_1 _16657_ (.A1(_06085_),
    .A2(_06091_),
    .B1(_06092_),
    .X(_06093_));
 sky130_fd_sc_hd__nor2_1 _16658_ (.A(_06087_),
    .B(_05952_),
    .Y(_06094_));
 sky130_fd_sc_hd__nor2_1 _16659_ (.A(_06093_),
    .B(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__nand2_2 _16660_ (.A(_06090_),
    .B(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__or2_1 _16661_ (.A(_05528_),
    .B(_05645_),
    .X(_06097_));
 sky130_fd_sc_hd__nand2_1 _16662_ (.A(_06097_),
    .B(_06070_),
    .Y(_06098_));
 sky130_fd_sc_hd__inv_2 _16663_ (.A(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__nand2_1 _16664_ (.A(_06099_),
    .B(net36),
    .Y(_06101_));
 sky130_fd_sc_hd__nand2_1 _16665_ (.A(_06098_),
    .B(_06012_),
    .Y(_06102_));
 sky130_fd_sc_hd__nand2_1 _16666_ (.A(_06101_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__inv_2 _16667_ (.A(_06103_),
    .Y(_06104_));
 sky130_fd_sc_hd__nand2_1 _16668_ (.A(_06096_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__nand2_1 _16669_ (.A(_06105_),
    .B(_06101_),
    .Y(_06106_));
 sky130_fd_sc_hd__xor2_1 _16670_ (.A(_06077_),
    .B(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__nand2_1 _16671_ (.A(_06107_),
    .B(_05916_),
    .Y(_06108_));
 sky130_fd_sc_hd__nand2_1 _16672_ (.A(net235),
    .B(_06074_),
    .Y(_06109_));
 sky130_fd_sc_hd__nand2_1 _16673_ (.A(_06108_),
    .B(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__nand2_1 _16674_ (.A(_06110_),
    .B(_08527_),
    .Y(_06112_));
 sky130_fd_sc_hd__nand3_2 _16675_ (.A(_06108_),
    .B(_08505_),
    .C(_06109_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand2_1 _16676_ (.A(_06112_),
    .B(_06113_),
    .Y(_06114_));
 sky130_fd_sc_hd__nand3_2 _16677_ (.A(_06104_),
    .B(_06075_),
    .C(_06076_),
    .Y(_06115_));
 sky130_fd_sc_hd__inv_2 _16678_ (.A(_06115_),
    .Y(_06116_));
 sky130_fd_sc_hd__nand2_1 _16679_ (.A(_06096_),
    .B(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__inv_2 _16680_ (.A(_05530_),
    .Y(_06118_));
 sky130_fd_sc_hd__nand2_1 _16681_ (.A(_05645_),
    .B(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__nand2_1 _16682_ (.A(_06119_),
    .B(_05516_),
    .Y(_06120_));
 sky130_fd_sc_hd__nand2_1 _16683_ (.A(_06120_),
    .B(_05520_),
    .Y(_06121_));
 sky130_fd_sc_hd__nand3_1 _16684_ (.A(_06119_),
    .B(_05519_),
    .C(_05516_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _16685_ (.A(_06121_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__nand2_1 _16686_ (.A(_06124_),
    .B(_06155_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand3_2 _16687_ (.A(_06121_),
    .B(net38),
    .C(_06123_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand2_1 _16688_ (.A(_06125_),
    .B(_06126_),
    .Y(_06127_));
 sky130_fd_sc_hd__inv_2 _16689_ (.A(_06101_),
    .Y(_06128_));
 sky130_fd_sc_hd__a21boi_2 _16690_ (.A1(_06075_),
    .A2(_06128_),
    .B1_N(_06076_),
    .Y(_06129_));
 sky130_fd_sc_hd__nand3_1 _16691_ (.A(_06117_),
    .B(_06127_),
    .C(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__clkinvlp_2 _16692_ (.A(_06130_),
    .Y(_06131_));
 sky130_fd_sc_hd__nand2_1 _16693_ (.A(_06117_),
    .B(_06129_),
    .Y(_06132_));
 sky130_fd_sc_hd__inv_2 _16694_ (.A(_06127_),
    .Y(_06134_));
 sky130_fd_sc_hd__nand2_1 _16695_ (.A(_06132_),
    .B(_06134_),
    .Y(_06135_));
 sky130_fd_sc_hd__nand2_1 _16696_ (.A(_06135_),
    .B(_05916_),
    .Y(_06136_));
 sky130_fd_sc_hd__or2_1 _16697_ (.A(_06124_),
    .B(_05916_),
    .X(_06137_));
 sky130_fd_sc_hd__o21ai_1 _16698_ (.A1(_06131_),
    .A2(_06136_),
    .B1(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__nand2b_1 _16699_ (.A_N(_06138_),
    .B(net137),
    .Y(_06139_));
 sky130_fd_sc_hd__nand2_1 _16700_ (.A(_06138_),
    .B(net121),
    .Y(_06140_));
 sky130_fd_sc_hd__nand2_1 _16701_ (.A(_06139_),
    .B(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__nor2_2 _16702_ (.A(_06114_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__nor2_1 _16703_ (.A(_06104_),
    .B(_06096_),
    .Y(_06143_));
 sky130_fd_sc_hd__nand2_1 _16704_ (.A(_05916_),
    .B(_06105_),
    .Y(_06145_));
 sky130_fd_sc_hd__nand2_1 _16705_ (.A(net235),
    .B(_06099_),
    .Y(_06146_));
 sky130_fd_sc_hd__o21ai_1 _16706_ (.A1(_06143_),
    .A2(_06145_),
    .B1(_06146_),
    .Y(_06147_));
 sky130_fd_sc_hd__or2_1 _16707_ (.A(_08384_),
    .B(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_8 _16708_ (.A(_08384_),
    .X(_06149_));
 sky130_fd_sc_hd__nand2_1 _16709_ (.A(_06147_),
    .B(_06149_),
    .Y(_06150_));
 sky130_fd_sc_hd__nand2_2 _16710_ (.A(_06148_),
    .B(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__nand2_1 _16711_ (.A(_06085_),
    .B(_06086_),
    .Y(_06152_));
 sky130_fd_sc_hd__a21o_1 _16712_ (.A1(_05956_),
    .A2(_05936_),
    .B1(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__nand3_1 _16713_ (.A(_05956_),
    .B(_06152_),
    .C(_05936_),
    .Y(_06154_));
 sky130_fd_sc_hd__a21o_1 _16714_ (.A1(_06153_),
    .A2(_06154_),
    .B1(net235),
    .X(_06156_));
 sky130_fd_sc_hd__nand2_1 _16715_ (.A(\div1i.quot[19] ),
    .B(_06084_),
    .Y(_06157_));
 sky130_fd_sc_hd__nand2_1 _16716_ (.A(_06156_),
    .B(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__buf_6 _16717_ (.A(_08274_),
    .X(_06159_));
 sky130_fd_sc_hd__nand2_1 _16718_ (.A(_06158_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__nand3_2 _16719_ (.A(_06156_),
    .B(_08296_),
    .C(_06157_),
    .Y(_06161_));
 sky130_fd_sc_hd__nand2_2 _16720_ (.A(_06160_),
    .B(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__nor2_2 _16721_ (.A(_06151_),
    .B(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__and2_1 _16722_ (.A(_06142_),
    .B(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__nand2_1 _16723_ (.A(_06069_),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__o21ai_2 _16724_ (.A1(_06161_),
    .A2(_06151_),
    .B1(_06150_),
    .Y(_06167_));
 sky130_fd_sc_hd__o21ai_1 _16725_ (.A1(_06113_),
    .A2(_06141_),
    .B1(_06140_),
    .Y(_06168_));
 sky130_fd_sc_hd__a21oi_1 _16726_ (.A1(_06167_),
    .A2(_06142_),
    .B1(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__nand2_2 _16727_ (.A(_06169_),
    .B(_06165_),
    .Y(_06170_));
 sky130_fd_sc_hd__nand2b_1 _16728_ (.A_N(_05693_),
    .B(_05732_),
    .Y(_06171_));
 sky130_fd_sc_hd__nand2_1 _16729_ (.A(_05693_),
    .B(_05733_),
    .Y(_06172_));
 sky130_fd_sc_hd__nand2_1 _16730_ (.A(_06171_),
    .B(_06172_),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_1 _16731_ (.A(_06173_),
    .B(_06737_),
    .Y(_06174_));
 sky130_fd_sc_hd__nand3_2 _16732_ (.A(_06171_),
    .B(_06726_),
    .C(_06172_),
    .Y(_06175_));
 sky130_fd_sc_hd__nand2_1 _16733_ (.A(_06174_),
    .B(_06175_),
    .Y(_06176_));
 sky130_fd_sc_hd__inv_4 _16734_ (.A(_06176_),
    .Y(_06178_));
 sky130_fd_sc_hd__nand2_1 _16735_ (.A(_06121_),
    .B(_05345_),
    .Y(_06179_));
 sky130_fd_sc_hd__nand2_1 _16736_ (.A(_05501_),
    .B(_05498_),
    .Y(_06180_));
 sky130_fd_sc_hd__inv_2 _16737_ (.A(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__nand2_1 _16738_ (.A(_06179_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__nand3_1 _16739_ (.A(_06121_),
    .B(_06180_),
    .C(_05345_),
    .Y(_06183_));
 sky130_fd_sc_hd__nand2_1 _16740_ (.A(_06182_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand2_1 _16741_ (.A(_06184_),
    .B(_05375_),
    .Y(_06185_));
 sky130_fd_sc_hd__inv_2 _16742_ (.A(_06126_),
    .Y(_06186_));
 sky130_fd_sc_hd__nand3_2 _16743_ (.A(_06182_),
    .B(net39),
    .C(_06183_),
    .Y(_06187_));
 sky130_fd_sc_hd__inv_2 _16744_ (.A(_06187_),
    .Y(_06189_));
 sky130_fd_sc_hd__a21o_1 _16745_ (.A1(_06185_),
    .A2(_06186_),
    .B1(_06189_),
    .X(_06190_));
 sky130_fd_sc_hd__nand3_1 _16746_ (.A(_06185_),
    .B(_06187_),
    .C(_06134_),
    .Y(_06191_));
 sky130_fd_sc_hd__nor2_1 _16747_ (.A(_06191_),
    .B(_06129_),
    .Y(_06192_));
 sky130_fd_sc_hd__nor2_1 _16748_ (.A(_06190_),
    .B(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__nor2_1 _16749_ (.A(_06115_),
    .B(_06191_),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_1 _16750_ (.A(_06194_),
    .B(_06096_),
    .Y(_06195_));
 sky130_fd_sc_hd__nand2_2 _16751_ (.A(_06193_),
    .B(_06195_),
    .Y(_06196_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(_05680_),
    .B(_05681_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_1 _16753_ (.A(_05647_),
    .B(_05687_),
    .Y(_06198_));
 sky130_fd_sc_hd__nand2_1 _16754_ (.A(_06198_),
    .B(_05684_),
    .Y(_06200_));
 sky130_fd_sc_hd__xor2_2 _16755_ (.A(_06197_),
    .B(_06200_),
    .X(_06201_));
 sky130_fd_sc_hd__inv_2 _16756_ (.A(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__nand2_1 _16757_ (.A(_06202_),
    .B(net41),
    .Y(_06203_));
 sky130_fd_sc_hd__or2_1 _16758_ (.A(_05687_),
    .B(_05647_),
    .X(_06204_));
 sky130_fd_sc_hd__nand2_1 _16759_ (.A(_06204_),
    .B(_06198_),
    .Y(_06205_));
 sky130_fd_sc_hd__inv_2 _16760_ (.A(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__buf_6 _16761_ (.A(net40),
    .X(_06207_));
 sky130_fd_sc_hd__nand2_1 _16762_ (.A(_06206_),
    .B(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__nand2_1 _16763_ (.A(_06205_),
    .B(_05408_),
    .Y(_06209_));
 sky130_fd_sc_hd__nand2_1 _16764_ (.A(_06208_),
    .B(_06209_),
    .Y(_06211_));
 sky130_fd_sc_hd__inv_2 _16765_ (.A(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__nand2_1 _16766_ (.A(_06201_),
    .B(_06814_),
    .Y(_06213_));
 sky130_fd_sc_hd__nand3_1 _16767_ (.A(_06203_),
    .B(_06212_),
    .C(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__inv_2 _16768_ (.A(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__nand2_1 _16769_ (.A(_06196_),
    .B(_06215_),
    .Y(_06216_));
 sky130_fd_sc_hd__inv_2 _16770_ (.A(_06208_),
    .Y(_06217_));
 sky130_fd_sc_hd__inv_2 _16771_ (.A(_06203_),
    .Y(_06218_));
 sky130_fd_sc_hd__a21oi_1 _16772_ (.A1(_06213_),
    .A2(_06217_),
    .B1(_06218_),
    .Y(_06219_));
 sky130_fd_sc_hd__nand2_1 _16773_ (.A(_06216_),
    .B(_06219_),
    .Y(_06220_));
 sky130_fd_sc_hd__or2_1 _16774_ (.A(_06178_),
    .B(_06220_),
    .X(_06222_));
 sky130_fd_sc_hd__buf_6 _16775_ (.A(_05916_),
    .X(_06223_));
 sky130_fd_sc_hd__nand2_1 _16776_ (.A(_06220_),
    .B(_06178_),
    .Y(_06224_));
 sky130_fd_sc_hd__nand3_1 _16777_ (.A(_06222_),
    .B(_06223_),
    .C(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__or2_1 _16778_ (.A(_06173_),
    .B(_05916_),
    .X(_06226_));
 sky130_fd_sc_hd__nand2_1 _16779_ (.A(_06225_),
    .B(_06226_),
    .Y(_06227_));
 sky130_fd_sc_hd__inv_2 _16780_ (.A(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__nand2_1 _16781_ (.A(_06228_),
    .B(_09987_),
    .Y(_06229_));
 sky130_fd_sc_hd__nand2_1 _16782_ (.A(_06227_),
    .B(_10009_),
    .Y(_06230_));
 sky130_fd_sc_hd__nand2_1 _16783_ (.A(_06229_),
    .B(_06230_),
    .Y(_06231_));
 sky130_fd_sc_hd__nand2_1 _16784_ (.A(_06203_),
    .B(_06213_),
    .Y(_06233_));
 sky130_fd_sc_hd__nand2_1 _16785_ (.A(_06196_),
    .B(_06212_),
    .Y(_06234_));
 sky130_fd_sc_hd__nand2_1 _16786_ (.A(_06234_),
    .B(_06208_),
    .Y(_06235_));
 sky130_fd_sc_hd__xor2_1 _16787_ (.A(_06233_),
    .B(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__nand2_1 _16788_ (.A(_06236_),
    .B(_06223_),
    .Y(_06237_));
 sky130_fd_sc_hd__nand2_1 _16789_ (.A(\div1i.quot[19] ),
    .B(_06201_),
    .Y(_06238_));
 sky130_fd_sc_hd__nand2_1 _16790_ (.A(_06237_),
    .B(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__nand2b_1 _16791_ (.A_N(_06239_),
    .B(net120),
    .Y(_06240_));
 sky130_fd_sc_hd__nand2_1 _16792_ (.A(_06239_),
    .B(_09735_),
    .Y(_06241_));
 sky130_fd_sc_hd__nand2_1 _16793_ (.A(_06240_),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__nor2_1 _16794_ (.A(_06231_),
    .B(_06242_),
    .Y(_06244_));
 sky130_fd_sc_hd__or2_1 _16795_ (.A(_06212_),
    .B(_06196_),
    .X(_06245_));
 sky130_fd_sc_hd__nand3_1 _16796_ (.A(_06245_),
    .B(_06223_),
    .C(_06234_),
    .Y(_06246_));
 sky130_fd_sc_hd__nand2_1 _16797_ (.A(\div1i.quot[19] ),
    .B(_06206_),
    .Y(_06247_));
 sky130_fd_sc_hd__nand2_1 _16798_ (.A(_06246_),
    .B(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__or2_1 _16799_ (.A(_09383_),
    .B(_06248_),
    .X(_06249_));
 sky130_fd_sc_hd__nand2_1 _16800_ (.A(_06248_),
    .B(_09383_),
    .Y(_06250_));
 sky130_fd_sc_hd__nand2_2 _16801_ (.A(_06249_),
    .B(_06250_),
    .Y(_06251_));
 sky130_fd_sc_hd__nand2_1 _16802_ (.A(_06185_),
    .B(_06187_),
    .Y(_06252_));
 sky130_fd_sc_hd__nand2_1 _16803_ (.A(_06135_),
    .B(_06126_),
    .Y(_06253_));
 sky130_fd_sc_hd__xor2_1 _16804_ (.A(_06252_),
    .B(_06253_),
    .X(_06255_));
 sky130_fd_sc_hd__nand2_1 _16805_ (.A(_06255_),
    .B(_06223_),
    .Y(_06256_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(\div1i.quot[19] ),
    .B(_06184_),
    .Y(_06257_));
 sky130_fd_sc_hd__nand2_1 _16807_ (.A(_06256_),
    .B(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__or2_1 _16808_ (.A(_09548_),
    .B(_06258_),
    .X(_06259_));
 sky130_fd_sc_hd__nand2_1 _16809_ (.A(_06258_),
    .B(_09548_),
    .Y(_06260_));
 sky130_fd_sc_hd__nand2_1 _16810_ (.A(_06259_),
    .B(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__nor2_1 _16811_ (.A(_06251_),
    .B(_06261_),
    .Y(_06262_));
 sky130_fd_sc_hd__nand3_2 _16812_ (.A(_06170_),
    .B(_06244_),
    .C(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__o21ai_2 _16813_ (.A1(_06251_),
    .A2(_06259_),
    .B1(_06250_),
    .Y(_06264_));
 sky130_fd_sc_hd__inv_2 _16814_ (.A(_06229_),
    .Y(_06266_));
 sky130_fd_sc_hd__o21ai_1 _16815_ (.A1(_06240_),
    .A2(_06266_),
    .B1(_06230_),
    .Y(_06267_));
 sky130_fd_sc_hd__a21oi_2 _16816_ (.A1(_06244_),
    .A2(_06264_),
    .B1(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_2 _16817_ (.A(_06263_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__a21o_1 _16818_ (.A1(_06172_),
    .A2(_05730_),
    .B1(_05737_),
    .X(_06270_));
 sky130_fd_sc_hd__nand3_1 _16819_ (.A(_06172_),
    .B(_05737_),
    .C(_05730_),
    .Y(_06271_));
 sky130_fd_sc_hd__nand2_1 _16820_ (.A(_06270_),
    .B(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(_06272_),
    .B(_06704_),
    .Y(_06273_));
 sky130_fd_sc_hd__inv_2 _16822_ (.A(_06175_),
    .Y(_06274_));
 sky130_fd_sc_hd__nand3_2 _16823_ (.A(_06270_),
    .B(net43),
    .C(_06271_),
    .Y(_06275_));
 sky130_fd_sc_hd__nand3_1 _16824_ (.A(_06273_),
    .B(_06274_),
    .C(_06275_),
    .Y(_06277_));
 sky130_fd_sc_hd__nand2_1 _16825_ (.A(_06277_),
    .B(_06275_),
    .Y(_06278_));
 sky130_fd_sc_hd__nand3_1 _16826_ (.A(_06273_),
    .B(_06178_),
    .C(_06275_),
    .Y(_06279_));
 sky130_fd_sc_hd__nor2_1 _16827_ (.A(_06219_),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__nor2_1 _16828_ (.A(_06278_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__inv_2 _16829_ (.A(_06279_),
    .Y(_06282_));
 sky130_fd_sc_hd__nand3_1 _16830_ (.A(_06282_),
    .B(_06196_),
    .C(_06215_),
    .Y(_06283_));
 sky130_fd_sc_hd__nand2_1 _16831_ (.A(_06281_),
    .B(_06283_),
    .Y(_06284_));
 sky130_fd_sc_hd__inv_2 _16832_ (.A(_05748_),
    .Y(_06285_));
 sky130_fd_sc_hd__or2_1 _16833_ (.A(_06285_),
    .B(_05740_),
    .X(_06286_));
 sky130_fd_sc_hd__nand2_1 _16834_ (.A(_05740_),
    .B(_06285_),
    .Y(_06288_));
 sky130_fd_sc_hd__nand2_1 _16835_ (.A(_06286_),
    .B(_06288_),
    .Y(_06289_));
 sky130_fd_sc_hd__inv_2 _16836_ (.A(_06289_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand2_1 _16837_ (.A(_06290_),
    .B(_06649_),
    .Y(_06291_));
 sky130_fd_sc_hd__nand2_1 _16838_ (.A(_06289_),
    .B(_10426_),
    .Y(_06292_));
 sky130_fd_sc_hd__nand2_1 _16839_ (.A(_06291_),
    .B(_06292_),
    .Y(_06293_));
 sky130_fd_sc_hd__inv_2 _16840_ (.A(_06293_),
    .Y(_06294_));
 sky130_fd_sc_hd__inv_2 _16841_ (.A(_05759_),
    .Y(_06295_));
 sky130_fd_sc_hd__nand2_1 _16842_ (.A(_06288_),
    .B(_05746_),
    .Y(_06296_));
 sky130_fd_sc_hd__or2_1 _16843_ (.A(_06295_),
    .B(_06296_),
    .X(_06297_));
 sky130_fd_sc_hd__nand2_1 _16844_ (.A(_06296_),
    .B(_06295_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2_1 _16845_ (.A(_06297_),
    .B(_06299_),
    .Y(_06300_));
 sky130_fd_sc_hd__nand2_1 _16846_ (.A(_06300_),
    .B(_06550_),
    .Y(_06301_));
 sky130_fd_sc_hd__nand3_1 _16847_ (.A(_06297_),
    .B(net46),
    .C(_06299_),
    .Y(_06302_));
 sky130_fd_sc_hd__nand3_1 _16848_ (.A(_06294_),
    .B(_06301_),
    .C(_06302_),
    .Y(_06303_));
 sky130_fd_sc_hd__inv_2 _16849_ (.A(_06303_),
    .Y(_06304_));
 sky130_fd_sc_hd__nand2_1 _16850_ (.A(_06284_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__inv_2 _16851_ (.A(_06301_),
    .Y(_06306_));
 sky130_fd_sc_hd__o21a_1 _16852_ (.A1(_06291_),
    .A2(_06306_),
    .B1(_06302_),
    .X(_06307_));
 sky130_fd_sc_hd__nand2_1 _16853_ (.A(_06305_),
    .B(_06307_),
    .Y(_06308_));
 sky130_fd_sc_hd__a21bo_1 _16854_ (.A1(_05740_),
    .A2(_05761_),
    .B1_N(_05821_),
    .X(_06310_));
 sky130_fd_sc_hd__or2_1 _16855_ (.A(_05814_),
    .B(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__nand2_1 _16856_ (.A(_06310_),
    .B(_05814_),
    .Y(_06312_));
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(_06311_),
    .B(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__inv_2 _16858_ (.A(_06313_),
    .Y(_06314_));
 sky130_fd_sc_hd__nand2_1 _16859_ (.A(_06314_),
    .B(net47),
    .Y(_06315_));
 sky130_fd_sc_hd__nand2_1 _16860_ (.A(_06313_),
    .B(_06594_),
    .Y(_06316_));
 sky130_fd_sc_hd__nand2_1 _16861_ (.A(_06315_),
    .B(_06316_),
    .Y(_06317_));
 sky130_fd_sc_hd__inv_2 _16862_ (.A(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__nand2_1 _16863_ (.A(_06308_),
    .B(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__nand3_1 _16864_ (.A(_06305_),
    .B(_06307_),
    .C(_06317_),
    .Y(_06321_));
 sky130_fd_sc_hd__nand3_1 _16865_ (.A(_06319_),
    .B(_06321_),
    .C(_06223_),
    .Y(_06322_));
 sky130_fd_sc_hd__nand2_1 _16866_ (.A(_06314_),
    .B(\div1i.quot[19] ),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(_06322_),
    .B(_06323_),
    .Y(_06324_));
 sky130_fd_sc_hd__nand2_2 _16868_ (.A(_06324_),
    .B(_10887_),
    .Y(_06325_));
 sky130_fd_sc_hd__nand3_2 _16869_ (.A(_06322_),
    .B(_10909_),
    .C(_06323_),
    .Y(_06326_));
 sky130_fd_sc_hd__nand2_4 _16870_ (.A(_06326_),
    .B(_06325_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand2_1 _16871_ (.A(_06224_),
    .B(_06175_),
    .Y(_06328_));
 sky130_fd_sc_hd__nand2_1 _16872_ (.A(_06273_),
    .B(_06275_),
    .Y(_06329_));
 sky130_fd_sc_hd__inv_2 _16873_ (.A(_06329_),
    .Y(_06330_));
 sky130_fd_sc_hd__nand2_1 _16874_ (.A(_06328_),
    .B(_06330_),
    .Y(_06332_));
 sky130_fd_sc_hd__nand3_1 _16875_ (.A(_06224_),
    .B(_06175_),
    .C(_06329_),
    .Y(_06333_));
 sky130_fd_sc_hd__nand2_1 _16876_ (.A(_06332_),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__nand2_1 _16877_ (.A(_06334_),
    .B(_06223_),
    .Y(_06335_));
 sky130_fd_sc_hd__nand2_1 _16878_ (.A(\div1i.quot[19] ),
    .B(_06272_),
    .Y(_06336_));
 sky130_fd_sc_hd__nand2_1 _16879_ (.A(_06335_),
    .B(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__nand2_1 _16880_ (.A(_06337_),
    .B(_10251_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand3_2 _16881_ (.A(_06335_),
    .B(_10240_),
    .C(_06336_),
    .Y(_06339_));
 sky130_fd_sc_hd__nand2_1 _16882_ (.A(_06338_),
    .B(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__inv_2 _16883_ (.A(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__nand2_1 _16884_ (.A(_06284_),
    .B(_06294_),
    .Y(_06343_));
 sky130_fd_sc_hd__nand3_1 _16885_ (.A(_06281_),
    .B(_06283_),
    .C(_06293_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand3_1 _16886_ (.A(_06343_),
    .B(_06223_),
    .C(_06344_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _16887_ (.A(\div1i.quot[19] ),
    .B(_06290_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand2_1 _16888_ (.A(_06345_),
    .B(_06346_),
    .Y(_06347_));
 sky130_fd_sc_hd__buf_6 _16889_ (.A(_10470_),
    .X(_06348_));
 sky130_fd_sc_hd__nand2_1 _16890_ (.A(_06347_),
    .B(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__nand3_1 _16891_ (.A(_06345_),
    .B(_10481_),
    .C(_06346_),
    .Y(_06350_));
 sky130_fd_sc_hd__nand2_2 _16892_ (.A(_06349_),
    .B(_06350_),
    .Y(_06351_));
 sky130_fd_sc_hd__inv_2 _16893_ (.A(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__nand2_1 _16894_ (.A(_06341_),
    .B(_06352_),
    .Y(_06354_));
 sky130_fd_sc_hd__nand2_1 _16895_ (.A(_06343_),
    .B(_06291_),
    .Y(_06355_));
 sky130_fd_sc_hd__nand2_1 _16896_ (.A(_06301_),
    .B(_06302_),
    .Y(_06356_));
 sky130_fd_sc_hd__inv_2 _16897_ (.A(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__nand2_1 _16898_ (.A(_06355_),
    .B(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand3_1 _16899_ (.A(_06343_),
    .B(_06356_),
    .C(_06291_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand2_1 _16900_ (.A(_06358_),
    .B(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand2_1 _16901_ (.A(_06360_),
    .B(_06223_),
    .Y(_06361_));
 sky130_fd_sc_hd__nand2_1 _16902_ (.A(_06300_),
    .B(\div1i.quot[19] ),
    .Y(_06362_));
 sky130_fd_sc_hd__nand2_1 _16903_ (.A(_06361_),
    .B(_06362_),
    .Y(_06363_));
 sky130_fd_sc_hd__nand2_1 _16904_ (.A(_06363_),
    .B(_10701_),
    .Y(_06365_));
 sky130_fd_sc_hd__buf_6 _16905_ (.A(_10690_),
    .X(_06366_));
 sky130_fd_sc_hd__nand3_1 _16906_ (.A(_06361_),
    .B(_06366_),
    .C(_06362_),
    .Y(_06367_));
 sky130_fd_sc_hd__nand2_1 _16907_ (.A(_06365_),
    .B(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__nor3_2 _16908_ (.A(_06327_),
    .B(_06354_),
    .C(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__nand2_2 _16909_ (.A(_06269_),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_1 _16910_ (.A(_06327_),
    .B(_06368_),
    .Y(_06371_));
 sky130_fd_sc_hd__o21ai_2 _16911_ (.A1(_06339_),
    .A2(_06351_),
    .B1(_06349_),
    .Y(_06372_));
 sky130_fd_sc_hd__inv_2 _16912_ (.A(_06326_),
    .Y(_06373_));
 sky130_fd_sc_hd__o21ai_1 _16913_ (.A1(_06367_),
    .A2(_06373_),
    .B1(_06325_),
    .Y(_06374_));
 sky130_fd_sc_hd__a21oi_2 _16914_ (.A1(_06371_),
    .A2(_06372_),
    .B1(_06374_),
    .Y(_06376_));
 sky130_fd_sc_hd__nand2_2 _16915_ (.A(_06370_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__nand2_1 _16916_ (.A(_05808_),
    .B(_05809_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_1 _16917_ (.A(_06312_),
    .B(_05811_),
    .Y(_06379_));
 sky130_fd_sc_hd__xor2_1 _16918_ (.A(_06378_),
    .B(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__nand3_1 _16919_ (.A(_06319_),
    .B(_06223_),
    .C(_06315_),
    .Y(_06381_));
 sky130_fd_sc_hd__xnor2_2 _16920_ (.A(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__nand2_4 _16921_ (.A(_06377_),
    .B(_06382_),
    .Y(_06383_));
 sky130_fd_sc_hd__clkinvlp_2 _16922_ (.A(_06382_),
    .Y(_06384_));
 sky130_fd_sc_hd__nand3_4 _16923_ (.A(_06370_),
    .B(_06376_),
    .C(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__nand2_8 _16924_ (.A(_06383_),
    .B(_06385_),
    .Y(_06387_));
 sky130_fd_sc_hd__buf_8 _16925_ (.A(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__buf_6 _16926_ (.A(_06388_),
    .X(\div1i.quot[18] ));
 sky130_fd_sc_hd__nand2_1 _16927_ (.A(_06060_),
    .B(net244),
    .Y(_06389_));
 sky130_fd_sc_hd__inv_2 _16928_ (.A(_06063_),
    .Y(_06390_));
 sky130_fd_sc_hd__nand2_1 _16929_ (.A(_06389_),
    .B(_06390_),
    .Y(_06391_));
 sky130_fd_sc_hd__nand2_2 _16930_ (.A(_06391_),
    .B(_05973_),
    .Y(_06392_));
 sky130_fd_sc_hd__nand2_1 _16931_ (.A(_06392_),
    .B(_06064_),
    .Y(_06393_));
 sky130_fd_sc_hd__nand2_1 _16932_ (.A(_06393_),
    .B(_05964_),
    .Y(_06394_));
 sky130_fd_sc_hd__nand3_1 _16933_ (.A(_06392_),
    .B(_05963_),
    .C(_06064_),
    .Y(_06395_));
 sky130_fd_sc_hd__nand2_1 _16934_ (.A(_06394_),
    .B(_06395_),
    .Y(_06397_));
 sky130_fd_sc_hd__nand2_1 _16935_ (.A(_06397_),
    .B(_05288_),
    .Y(_06398_));
 sky130_fd_sc_hd__nand3_1 _16936_ (.A(_06389_),
    .B(_05972_),
    .C(_06390_),
    .Y(_06399_));
 sky130_fd_sc_hd__nand3_2 _16937_ (.A(_06392_),
    .B(net34),
    .C(_06399_),
    .Y(_06400_));
 sky130_fd_sc_hd__inv_2 _16938_ (.A(_06400_),
    .Y(_06401_));
 sky130_fd_sc_hd__nand3_2 _16939_ (.A(_06394_),
    .B(net35),
    .C(_06395_),
    .Y(_06402_));
 sky130_fd_sc_hd__nand3_1 _16940_ (.A(_06398_),
    .B(_06401_),
    .C(_06402_),
    .Y(_06403_));
 sky130_fd_sc_hd__nand2_1 _16941_ (.A(_06403_),
    .B(_06402_),
    .Y(_06404_));
 sky130_fd_sc_hd__inv_2 _16942_ (.A(_05926_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_1 _16943_ (.A(_06060_),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand2_1 _16944_ (.A(_06406_),
    .B(_05923_),
    .Y(_06408_));
 sky130_fd_sc_hd__inv_2 _16945_ (.A(_05914_),
    .Y(_06409_));
 sky130_fd_sc_hd__nand2_1 _16946_ (.A(_06408_),
    .B(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__nand3_1 _16947_ (.A(_06406_),
    .B(_05914_),
    .C(_05923_),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_1 _16948_ (.A(_06410_),
    .B(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__nand2_1 _16949_ (.A(_06412_),
    .B(_05310_),
    .Y(_06413_));
 sky130_fd_sc_hd__or2_1 _16950_ (.A(_06405_),
    .B(_06060_),
    .X(_06414_));
 sky130_fd_sc_hd__nand2_1 _16951_ (.A(_06414_),
    .B(_06406_),
    .Y(_06415_));
 sky130_fd_sc_hd__inv_2 _16952_ (.A(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__nand2_1 _16953_ (.A(_06416_),
    .B(net63),
    .Y(_06417_));
 sky130_fd_sc_hd__inv_2 _16954_ (.A(_06417_),
    .Y(_06419_));
 sky130_fd_sc_hd__inv_2 _16955_ (.A(_06412_),
    .Y(_06420_));
 sky130_fd_sc_hd__nand2_1 _16956_ (.A(_06420_),
    .B(net64),
    .Y(_06421_));
 sky130_fd_sc_hd__inv_2 _16957_ (.A(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__a21oi_2 _16958_ (.A1(_06413_),
    .A2(_06419_),
    .B1(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__nand2_1 _16959_ (.A(_06392_),
    .B(_06399_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand2_1 _16960_ (.A(_06424_),
    .B(_05299_),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _16961_ (.A(_06425_),
    .B(_06400_),
    .Y(_06426_));
 sky130_fd_sc_hd__inv_2 _16962_ (.A(_06426_),
    .Y(_06427_));
 sky130_fd_sc_hd__nand3_1 _16963_ (.A(_06398_),
    .B(_06427_),
    .C(_06402_),
    .Y(_06428_));
 sky130_fd_sc_hd__nor2_1 _16964_ (.A(_06423_),
    .B(_06428_),
    .Y(_06430_));
 sky130_fd_sc_hd__nor2_1 _16965_ (.A(_06404_),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__inv_2 _16966_ (.A(_06428_),
    .Y(_06432_));
 sky130_fd_sc_hd__nand2_1 _16967_ (.A(_05993_),
    .B(_05996_),
    .Y(_06433_));
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(_06433_),
    .B(_05997_),
    .Y(_06434_));
 sky130_fd_sc_hd__nand2_1 _16969_ (.A(_06434_),
    .B(_05999_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(_06435_),
    .B(_05189_),
    .Y(_06436_));
 sky130_fd_sc_hd__o21ai_1 _16971_ (.A1(_05496_),
    .A2(\div1i.quot[19] ),
    .B1(_05474_),
    .Y(_06437_));
 sky130_fd_sc_hd__nand3_1 _16972_ (.A(_06434_),
    .B(net55),
    .C(_05999_),
    .Y(_06438_));
 sky130_fd_sc_hd__inv_2 _16973_ (.A(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__a21o_1 _16974_ (.A1(_06436_),
    .A2(_06437_),
    .B1(_06439_),
    .X(_06441_));
 sky130_fd_sc_hd__nand2_1 _16975_ (.A(_06000_),
    .B(_05984_),
    .Y(_06442_));
 sky130_fd_sc_hd__nand2_1 _16976_ (.A(_05999_),
    .B(_05993_),
    .Y(_06443_));
 sky130_fd_sc_hd__xor2_2 _16977_ (.A(_06442_),
    .B(_06443_),
    .X(_06444_));
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(_06444_),
    .B(_05178_),
    .Y(_06445_));
 sky130_fd_sc_hd__nand2_1 _16979_ (.A(_06441_),
    .B(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__inv_2 _16980_ (.A(_06444_),
    .Y(_06447_));
 sky130_fd_sc_hd__nand2_1 _16981_ (.A(_06447_),
    .B(net58),
    .Y(_06448_));
 sky130_fd_sc_hd__nand2_1 _16982_ (.A(_06446_),
    .B(_06448_),
    .Y(_06449_));
 sky130_fd_sc_hd__nand2_1 _16983_ (.A(_05995_),
    .B(_05999_),
    .Y(_06450_));
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(_06450_),
    .B(_06000_),
    .Y(_06452_));
 sky130_fd_sc_hd__nand2_1 _16985_ (.A(_06452_),
    .B(_06048_),
    .Y(_06453_));
 sky130_fd_sc_hd__nand3_1 _16986_ (.A(_06450_),
    .B(_06000_),
    .C(_06049_),
    .Y(_06454_));
 sky130_fd_sc_hd__nand2_1 _16987_ (.A(_06453_),
    .B(_06454_),
    .Y(_06455_));
 sky130_fd_sc_hd__nand2_1 _16988_ (.A(_06455_),
    .B(_05705_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand3_1 _16989_ (.A(_06453_),
    .B(net59),
    .C(_06454_),
    .Y(_06457_));
 sky130_fd_sc_hd__nand2_1 _16990_ (.A(_06456_),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__inv_2 _16991_ (.A(_06458_),
    .Y(_06459_));
 sky130_fd_sc_hd__nand2_1 _16992_ (.A(_06449_),
    .B(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__nand2_1 _16993_ (.A(_06460_),
    .B(_06457_),
    .Y(_06461_));
 sky130_fd_sc_hd__nand2_1 _16994_ (.A(_06454_),
    .B(_06044_),
    .Y(_06463_));
 sky130_fd_sc_hd__xor2_2 _16995_ (.A(_06037_),
    .B(_06463_),
    .X(_06464_));
 sky130_fd_sc_hd__buf_6 _16996_ (.A(_05738_),
    .X(_06465_));
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(_06464_),
    .B(_06465_),
    .Y(_06466_));
 sky130_fd_sc_hd__nand2_1 _16998_ (.A(_06461_),
    .B(_06466_),
    .Y(_06467_));
 sky130_fd_sc_hd__or2_1 _16999_ (.A(_05738_),
    .B(_06464_),
    .X(_06468_));
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(_06467_),
    .B(_06468_),
    .Y(_06469_));
 sky130_fd_sc_hd__nor2_1 _17001_ (.A(_06037_),
    .B(_06048_),
    .Y(_06470_));
 sky130_fd_sc_hd__nand3_1 _17002_ (.A(_06450_),
    .B(_06470_),
    .C(_06000_),
    .Y(_06471_));
 sky130_fd_sc_hd__inv_2 _17003_ (.A(_06054_),
    .Y(_06472_));
 sky130_fd_sc_hd__nand2_1 _17004_ (.A(_06471_),
    .B(_06472_),
    .Y(_06474_));
 sky130_fd_sc_hd__nand2_2 _17005_ (.A(_06474_),
    .B(_06024_),
    .Y(_06475_));
 sky130_fd_sc_hd__nand2_1 _17006_ (.A(_06475_),
    .B(_06020_),
    .Y(_06476_));
 sky130_fd_sc_hd__nand2_1 _17007_ (.A(_06476_),
    .B(_06014_),
    .Y(_06477_));
 sky130_fd_sc_hd__nand3_2 _17008_ (.A(_06475_),
    .B(_06013_),
    .C(_06020_),
    .Y(_06478_));
 sky130_fd_sc_hd__nand2_1 _17009_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__nand2_1 _17010_ (.A(_06479_),
    .B(_05255_),
    .Y(_06480_));
 sky130_fd_sc_hd__nand3_1 _17011_ (.A(_06471_),
    .B(_06022_),
    .C(_06472_),
    .Y(_06481_));
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(_06475_),
    .B(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__nand2_1 _17013_ (.A(_06482_),
    .B(_05847_),
    .Y(_06483_));
 sky130_fd_sc_hd__nand3_2 _17014_ (.A(_06475_),
    .B(net61),
    .C(_06481_),
    .Y(_06485_));
 sky130_fd_sc_hd__nand2_1 _17015_ (.A(_06483_),
    .B(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__inv_2 _17016_ (.A(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__nand3_1 _17017_ (.A(_06477_),
    .B(_05896_),
    .C(_06478_),
    .Y(_06488_));
 sky130_fd_sc_hd__nand3_1 _17018_ (.A(_06480_),
    .B(_06487_),
    .C(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__inv_2 _17019_ (.A(_06489_),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_1 _17020_ (.A(_06469_),
    .B(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__inv_2 _17021_ (.A(_06485_),
    .Y(_06492_));
 sky130_fd_sc_hd__a21boi_1 _17022_ (.A1(_06480_),
    .A2(_06492_),
    .B1_N(_06488_),
    .Y(_06493_));
 sky130_fd_sc_hd__nand2_1 _17023_ (.A(_06491_),
    .B(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__nand2_1 _17024_ (.A(_06421_),
    .B(_06413_),
    .Y(_06496_));
 sky130_fd_sc_hd__inv_2 _17025_ (.A(_06496_),
    .Y(_06497_));
 sky130_fd_sc_hd__nand2_1 _17026_ (.A(_06415_),
    .B(_05321_),
    .Y(_06498_));
 sky130_fd_sc_hd__nand2_1 _17027_ (.A(_06417_),
    .B(_06498_),
    .Y(_06499_));
 sky130_fd_sc_hd__inv_2 _17028_ (.A(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__nand2_1 _17029_ (.A(_06497_),
    .B(_06500_),
    .Y(_06501_));
 sky130_fd_sc_hd__inv_2 _17030_ (.A(_06501_),
    .Y(_06502_));
 sky130_fd_sc_hd__nand3_1 _17031_ (.A(_06432_),
    .B(_06494_),
    .C(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__nand2_1 _17032_ (.A(_06431_),
    .B(_06503_),
    .Y(_06504_));
 sky130_fd_sc_hd__inv_2 _17033_ (.A(_06151_),
    .Y(_06505_));
 sky130_fd_sc_hd__inv_2 _17034_ (.A(_06162_),
    .Y(_06507_));
 sky130_fd_sc_hd__nand2_1 _17035_ (.A(_06069_),
    .B(_06507_),
    .Y(_06508_));
 sky130_fd_sc_hd__nand2_1 _17036_ (.A(_06508_),
    .B(_06161_),
    .Y(_06509_));
 sky130_fd_sc_hd__or2_1 _17037_ (.A(_06505_),
    .B(_06509_),
    .X(_06510_));
 sky130_fd_sc_hd__nand2_1 _17038_ (.A(_06509_),
    .B(_06505_),
    .Y(_06511_));
 sky130_fd_sc_hd__nand2_1 _17039_ (.A(_06510_),
    .B(_06511_),
    .Y(_06512_));
 sky130_fd_sc_hd__nand2_1 _17040_ (.A(_06512_),
    .B(_06045_),
    .Y(_06513_));
 sky130_fd_sc_hd__nand3_1 _17041_ (.A(_06510_),
    .B(net37),
    .C(_06511_),
    .Y(_06514_));
 sky130_fd_sc_hd__nand2_1 _17042_ (.A(_06513_),
    .B(_06514_),
    .Y(_06515_));
 sky130_fd_sc_hd__inv_2 _17043_ (.A(_06515_),
    .Y(_06516_));
 sky130_fd_sc_hd__or2_1 _17044_ (.A(_06507_),
    .B(_06069_),
    .X(_06518_));
 sky130_fd_sc_hd__nand2_1 _17045_ (.A(_06518_),
    .B(_06508_),
    .Y(_06519_));
 sky130_fd_sc_hd__inv_2 _17046_ (.A(_06519_),
    .Y(_06520_));
 sky130_fd_sc_hd__buf_6 _17047_ (.A(net36),
    .X(_06521_));
 sky130_fd_sc_hd__nand2_1 _17048_ (.A(_06520_),
    .B(_06521_),
    .Y(_06522_));
 sky130_fd_sc_hd__nand2_1 _17049_ (.A(_06519_),
    .B(_06012_),
    .Y(_06523_));
 sky130_fd_sc_hd__nand2_1 _17050_ (.A(_06522_),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__inv_4 _17051_ (.A(_06524_),
    .Y(_06525_));
 sky130_fd_sc_hd__nand2_1 _17052_ (.A(_06516_),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__inv_4 _17053_ (.A(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__nand2_1 _17054_ (.A(_06504_),
    .B(_06527_),
    .Y(_06529_));
 sky130_fd_sc_hd__inv_2 _17055_ (.A(_06522_),
    .Y(_06530_));
 sky130_fd_sc_hd__a21boi_2 _17056_ (.A1(_06513_),
    .A2(_06530_),
    .B1_N(_06514_),
    .Y(_06531_));
 sky130_fd_sc_hd__nand2_1 _17057_ (.A(_06529_),
    .B(_06531_),
    .Y(_06532_));
 sky130_fd_sc_hd__nand2_1 _17058_ (.A(_06069_),
    .B(_06163_),
    .Y(_06533_));
 sky130_fd_sc_hd__inv_2 _17059_ (.A(_06167_),
    .Y(_06534_));
 sky130_fd_sc_hd__nand2_1 _17060_ (.A(_06533_),
    .B(_06534_),
    .Y(_06535_));
 sky130_fd_sc_hd__inv_2 _17061_ (.A(_06114_),
    .Y(_06536_));
 sky130_fd_sc_hd__nand2_1 _17062_ (.A(_06535_),
    .B(_06536_),
    .Y(_06537_));
 sky130_fd_sc_hd__nand3_1 _17063_ (.A(_06533_),
    .B(_06114_),
    .C(_06534_),
    .Y(_06538_));
 sky130_fd_sc_hd__nand2_1 _17064_ (.A(_06537_),
    .B(_06538_),
    .Y(_06540_));
 sky130_fd_sc_hd__inv_2 _17065_ (.A(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__nand2_1 _17066_ (.A(_06541_),
    .B(net38),
    .Y(_06542_));
 sky130_fd_sc_hd__nand2_1 _17067_ (.A(_06540_),
    .B(_06155_),
    .Y(_06543_));
 sky130_fd_sc_hd__nand2_1 _17068_ (.A(_06542_),
    .B(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__inv_2 _17069_ (.A(_06544_),
    .Y(_06545_));
 sky130_fd_sc_hd__nand2_1 _17070_ (.A(_06532_),
    .B(_06545_),
    .Y(_06546_));
 sky130_fd_sc_hd__inv_4 _17071_ (.A(_06387_),
    .Y(_06547_));
 sky130_fd_sc_hd__buf_6 _17072_ (.A(_06547_),
    .X(_06548_));
 sky130_fd_sc_hd__nand3_1 _17073_ (.A(_06529_),
    .B(_06544_),
    .C(_06531_),
    .Y(_06549_));
 sky130_fd_sc_hd__nand3_1 _17074_ (.A(_06546_),
    .B(_06548_),
    .C(_06549_),
    .Y(_06551_));
 sky130_fd_sc_hd__nand2_1 _17075_ (.A(_06388_),
    .B(_06541_),
    .Y(_06552_));
 sky130_fd_sc_hd__nand2_1 _17076_ (.A(_06551_),
    .B(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__buf_6 _17077_ (.A(net121),
    .X(_06554_));
 sky130_fd_sc_hd__nand2_1 _17078_ (.A(_06553_),
    .B(_06554_),
    .Y(_06555_));
 sky130_fd_sc_hd__buf_6 _17079_ (.A(net137),
    .X(_06556_));
 sky130_fd_sc_hd__nand3_1 _17080_ (.A(_06551_),
    .B(_06556_),
    .C(_06552_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_1 _17081_ (.A(_06555_),
    .B(_06557_),
    .Y(_06558_));
 sky130_fd_sc_hd__nand2_1 _17082_ (.A(_06504_),
    .B(_06525_),
    .Y(_06559_));
 sky130_fd_sc_hd__nand2_1 _17083_ (.A(_06559_),
    .B(_06522_),
    .Y(_06560_));
 sky130_fd_sc_hd__nand2_1 _17084_ (.A(_06560_),
    .B(_06516_),
    .Y(_06562_));
 sky130_fd_sc_hd__nand3_1 _17085_ (.A(_06559_),
    .B(_06515_),
    .C(_06522_),
    .Y(_06563_));
 sky130_fd_sc_hd__nand2_1 _17086_ (.A(_06562_),
    .B(_06563_),
    .Y(_06564_));
 sky130_fd_sc_hd__nand2_1 _17087_ (.A(_06564_),
    .B(_06548_),
    .Y(_06565_));
 sky130_fd_sc_hd__nand2_1 _17088_ (.A(_06388_),
    .B(_06512_),
    .Y(_06566_));
 sky130_fd_sc_hd__nand2_1 _17089_ (.A(_06565_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__buf_6 _17090_ (.A(_08527_),
    .X(_06568_));
 sky130_fd_sc_hd__nand2_1 _17091_ (.A(_06567_),
    .B(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__clkbuf_8 _17092_ (.A(_08505_),
    .X(_06570_));
 sky130_fd_sc_hd__nand3_2 _17093_ (.A(_06565_),
    .B(_06570_),
    .C(_06566_),
    .Y(_06571_));
 sky130_fd_sc_hd__nand2_1 _17094_ (.A(_06569_),
    .B(_06571_),
    .Y(_06573_));
 sky130_fd_sc_hd__nor2_1 _17095_ (.A(_06558_),
    .B(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__nand2_1 _17096_ (.A(_06502_),
    .B(_06494_),
    .Y(_06575_));
 sky130_fd_sc_hd__nand2_1 _17097_ (.A(_06575_),
    .B(_06423_),
    .Y(_06576_));
 sky130_fd_sc_hd__nand2_1 _17098_ (.A(_06576_),
    .B(_06427_),
    .Y(_06577_));
 sky130_fd_sc_hd__nand2_1 _17099_ (.A(_06577_),
    .B(_06400_),
    .Y(_06578_));
 sky130_fd_sc_hd__nand3_1 _17100_ (.A(_06578_),
    .B(_06402_),
    .C(_06398_),
    .Y(_06579_));
 sky130_fd_sc_hd__nand2_1 _17101_ (.A(_06398_),
    .B(_06402_),
    .Y(_06580_));
 sky130_fd_sc_hd__nand3_1 _17102_ (.A(_06577_),
    .B(_06400_),
    .C(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__nand2_1 _17103_ (.A(_06579_),
    .B(_06581_),
    .Y(_06582_));
 sky130_fd_sc_hd__nand2_1 _17104_ (.A(_06582_),
    .B(_06548_),
    .Y(_06584_));
 sky130_fd_sc_hd__nand2_1 _17105_ (.A(\div1i.quot[18] ),
    .B(_06397_),
    .Y(_06585_));
 sky130_fd_sc_hd__nand3_1 _17106_ (.A(_06584_),
    .B(_08296_),
    .C(_06585_),
    .Y(_06586_));
 sky130_fd_sc_hd__or2_1 _17107_ (.A(_06525_),
    .B(_06504_),
    .X(_06587_));
 sky130_fd_sc_hd__nand3_1 _17108_ (.A(_06587_),
    .B(_06548_),
    .C(_06559_),
    .Y(_06588_));
 sky130_fd_sc_hd__nand2_1 _17109_ (.A(_06388_),
    .B(_06520_),
    .Y(_06589_));
 sky130_fd_sc_hd__nand3_1 _17110_ (.A(_06588_),
    .B(_08406_),
    .C(_06589_),
    .Y(_06590_));
 sky130_fd_sc_hd__inv_2 _17111_ (.A(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__buf_6 _17112_ (.A(_08406_),
    .X(_06592_));
 sky130_fd_sc_hd__a21o_1 _17113_ (.A1(_06588_),
    .A2(_06589_),
    .B1(_06592_),
    .X(_06593_));
 sky130_fd_sc_hd__o21ai_1 _17114_ (.A1(_06586_),
    .A2(_06591_),
    .B1(_06593_),
    .Y(_06595_));
 sky130_fd_sc_hd__inv_2 _17115_ (.A(_06557_),
    .Y(_06596_));
 sky130_fd_sc_hd__o21ai_1 _17116_ (.A1(_06571_),
    .A2(_06596_),
    .B1(_06555_),
    .Y(_06597_));
 sky130_fd_sc_hd__a21oi_1 _17117_ (.A1(_06574_),
    .A2(_06595_),
    .B1(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__inv_2 _17118_ (.A(_06435_),
    .Y(_06599_));
 sky130_fd_sc_hd__nand2_1 _17119_ (.A(_06388_),
    .B(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__nand2_1 _17120_ (.A(_06436_),
    .B(_06438_),
    .Y(_06601_));
 sky130_fd_sc_hd__xor2_1 _17121_ (.A(_06437_),
    .B(_06601_),
    .X(_06602_));
 sky130_fd_sc_hd__nand3b_1 _17122_ (.A_N(_06602_),
    .B(net130),
    .C(net138),
    .Y(_06603_));
 sky130_fd_sc_hd__nand2_1 _17123_ (.A(_06600_),
    .B(_06603_),
    .Y(_06604_));
 sky130_fd_sc_hd__nand2_1 _17124_ (.A(_06604_),
    .B(_05983_),
    .Y(_06606_));
 sky130_fd_sc_hd__clkbuf_4 _17125_ (.A(_07242_),
    .X(_06607_));
 sky130_fd_sc_hd__nor2_1 _17126_ (.A(_05496_),
    .B(_06223_),
    .Y(_06608_));
 sky130_fd_sc_hd__or2_1 _17127_ (.A(_06607_),
    .B(_06608_),
    .X(_06609_));
 sky130_fd_sc_hd__nand2_1 _17128_ (.A(_06609_),
    .B(_05997_),
    .Y(_06610_));
 sky130_fd_sc_hd__inv_2 _17129_ (.A(_06610_),
    .Y(_06611_));
 sky130_fd_sc_hd__nand2_1 _17130_ (.A(_06388_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__nand3_1 _17131_ (.A(net128),
    .B(net138),
    .C(_06608_),
    .Y(_06613_));
 sky130_fd_sc_hd__nand2_1 _17132_ (.A(_06612_),
    .B(_06613_),
    .Y(_06614_));
 sky130_fd_sc_hd__buf_6 _17133_ (.A(_07539_),
    .X(_06615_));
 sky130_fd_sc_hd__nand2_2 _17134_ (.A(_06614_),
    .B(_06615_),
    .Y(_06617_));
 sky130_fd_sc_hd__nand2_1 _17135_ (.A(_06606_),
    .B(_06617_),
    .Y(_06618_));
 sky130_fd_sc_hd__inv_2 _17136_ (.A(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__buf_6 _17137_ (.A(_07560_),
    .X(_06620_));
 sky130_fd_sc_hd__nand3_1 _17138_ (.A(_06612_),
    .B(_06620_),
    .C(_06613_),
    .Y(_06621_));
 sky130_fd_sc_hd__nand3_2 _17139_ (.A(_06388_),
    .B(_05474_),
    .C(_07308_),
    .Y(_06622_));
 sky130_fd_sc_hd__inv_2 _17140_ (.A(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__nand3_2 _17141_ (.A(_06617_),
    .B(_06621_),
    .C(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__or2_4 _17142_ (.A(_05983_),
    .B(_06604_),
    .X(_06625_));
 sky130_fd_sc_hd__a21boi_2 _17143_ (.A1(_06619_),
    .A2(_06624_),
    .B1_N(_06625_),
    .Y(_06626_));
 sky130_fd_sc_hd__inv_2 _17144_ (.A(_06482_),
    .Y(_06628_));
 sky130_fd_sc_hd__nand2_1 _17145_ (.A(_06387_),
    .B(_06628_),
    .Y(_06629_));
 sky130_fd_sc_hd__nand2_1 _17146_ (.A(_06469_),
    .B(_06487_),
    .Y(_06630_));
 sky130_fd_sc_hd__nand3_1 _17147_ (.A(_06467_),
    .B(_06486_),
    .C(_06468_),
    .Y(_06631_));
 sky130_fd_sc_hd__nand2_1 _17148_ (.A(_06630_),
    .B(_06631_),
    .Y(_06632_));
 sky130_fd_sc_hd__inv_2 _17149_ (.A(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__nand3_1 _17150_ (.A(_06383_),
    .B(net138),
    .C(_06633_),
    .Y(_06634_));
 sky130_fd_sc_hd__nand2_1 _17151_ (.A(_06629_),
    .B(_06634_),
    .Y(_06635_));
 sky130_fd_sc_hd__buf_6 _17152_ (.A(_13588_),
    .X(_06636_));
 sky130_fd_sc_hd__nand2_1 _17153_ (.A(_06635_),
    .B(_06636_),
    .Y(_06637_));
 sky130_fd_sc_hd__buf_6 _17154_ (.A(_11579_),
    .X(_06639_));
 sky130_fd_sc_hd__nand3_1 _17155_ (.A(_06629_),
    .B(_06639_),
    .C(_06634_),
    .Y(_06640_));
 sky130_fd_sc_hd__nand2_1 _17156_ (.A(_06637_),
    .B(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__inv_2 _17157_ (.A(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__nand2_1 _17158_ (.A(_06388_),
    .B(_06464_),
    .Y(_06643_));
 sky130_fd_sc_hd__nand2_1 _17159_ (.A(_06468_),
    .B(_06466_),
    .Y(_06644_));
 sky130_fd_sc_hd__xor2_1 _17160_ (.A(_06461_),
    .B(_06644_),
    .X(_06645_));
 sky130_fd_sc_hd__nand3_1 _17161_ (.A(net128),
    .B(net138),
    .C(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__nand2_1 _17162_ (.A(_06643_),
    .B(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__buf_6 _17163_ (.A(_08066_),
    .X(_06648_));
 sky130_fd_sc_hd__nand2_1 _17164_ (.A(_06647_),
    .B(_06648_),
    .Y(_06650_));
 sky130_fd_sc_hd__clkbuf_8 _17165_ (.A(_08055_),
    .X(_06651_));
 sky130_fd_sc_hd__nand3_1 _17166_ (.A(_06643_),
    .B(_06651_),
    .C(_06646_),
    .Y(_06652_));
 sky130_fd_sc_hd__nand2_2 _17167_ (.A(_06650_),
    .B(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__inv_2 _17168_ (.A(_06653_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2_1 _17169_ (.A(_06642_),
    .B(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__inv_2 _17170_ (.A(_06455_),
    .Y(_06656_));
 sky130_fd_sc_hd__nand2_1 _17171_ (.A(net231),
    .B(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__or2_1 _17172_ (.A(_06459_),
    .B(_06449_),
    .X(_06658_));
 sky130_fd_sc_hd__nand2_1 _17173_ (.A(_06658_),
    .B(_06460_),
    .Y(_06659_));
 sky130_fd_sc_hd__inv_2 _17174_ (.A(_06659_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand3_1 _17175_ (.A(net128),
    .B(net138),
    .C(_06661_),
    .Y(_06662_));
 sky130_fd_sc_hd__nand2_1 _17176_ (.A(_06657_),
    .B(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__nand2_1 _17177_ (.A(_06663_),
    .B(_06033_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand3_1 _17178_ (.A(_06657_),
    .B(_12051_),
    .C(_06662_),
    .Y(_06665_));
 sky130_fd_sc_hd__nand2_1 _17179_ (.A(_06664_),
    .B(_06665_),
    .Y(_06666_));
 sky130_fd_sc_hd__inv_2 _17180_ (.A(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__nand2_1 _17181_ (.A(net231),
    .B(_06447_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_1 _17182_ (.A(_06448_),
    .B(_06445_),
    .Y(_06669_));
 sky130_fd_sc_hd__xnor2_1 _17183_ (.A(_06441_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand3_1 _17184_ (.A(net128),
    .B(net138),
    .C(_06670_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand2_1 _17185_ (.A(_06668_),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__nand2_2 _17186_ (.A(_06673_),
    .B(_07725_),
    .Y(_06674_));
 sky130_fd_sc_hd__nand3_1 _17187_ (.A(_06668_),
    .B(_06046_),
    .C(_06672_),
    .Y(_06675_));
 sky130_fd_sc_hd__nand2_2 _17188_ (.A(_06674_),
    .B(_06675_),
    .Y(_06676_));
 sky130_fd_sc_hd__clkinv_1 _17189_ (.A(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand2_1 _17190_ (.A(_06667_),
    .B(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__nor2_1 _17191_ (.A(_06655_),
    .B(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__nand2_1 _17192_ (.A(_06626_),
    .B(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__inv_2 _17193_ (.A(_06665_),
    .Y(_06681_));
 sky130_fd_sc_hd__o21ai_2 _17194_ (.A1(_06674_),
    .A2(_06681_),
    .B1(_06664_),
    .Y(_06683_));
 sky130_fd_sc_hd__nor2_1 _17195_ (.A(_06641_),
    .B(_06653_),
    .Y(_06684_));
 sky130_fd_sc_hd__inv_2 _17196_ (.A(_06640_),
    .Y(_06685_));
 sky130_fd_sc_hd__o21ai_1 _17197_ (.A1(_06652_),
    .A2(_06685_),
    .B1(_06637_),
    .Y(_06686_));
 sky130_fd_sc_hd__a21oi_1 _17198_ (.A1(_06683_),
    .A2(_06684_),
    .B1(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__nand2_2 _17199_ (.A(_06680_),
    .B(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__nand2_1 _17200_ (.A(_06494_),
    .B(_06500_),
    .Y(_06689_));
 sky130_fd_sc_hd__or2_1 _17201_ (.A(_06500_),
    .B(_06494_),
    .X(_06690_));
 sky130_fd_sc_hd__nand3_1 _17202_ (.A(_06547_),
    .B(_06689_),
    .C(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__nand2_1 _17203_ (.A(_06387_),
    .B(_06416_),
    .Y(_06692_));
 sky130_fd_sc_hd__nand2_1 _17204_ (.A(_06691_),
    .B(_06692_),
    .Y(_06694_));
 sky130_fd_sc_hd__buf_6 _17205_ (.A(_11140_),
    .X(_06695_));
 sky130_fd_sc_hd__nand2_1 _17206_ (.A(_06694_),
    .B(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__buf_6 _17207_ (.A(_08746_),
    .X(_06697_));
 sky130_fd_sc_hd__nand3_1 _17208_ (.A(_06691_),
    .B(_06697_),
    .C(_06692_),
    .Y(_06698_));
 sky130_fd_sc_hd__nand2_1 _17209_ (.A(_06696_),
    .B(_06698_),
    .Y(_06699_));
 sky130_fd_sc_hd__inv_2 _17210_ (.A(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__nand2_1 _17211_ (.A(_06480_),
    .B(_06488_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand2_1 _17212_ (.A(_06630_),
    .B(_06485_),
    .Y(_06702_));
 sky130_fd_sc_hd__xor2_1 _17213_ (.A(_06701_),
    .B(_06702_),
    .X(_06703_));
 sky130_fd_sc_hd__nand2_1 _17214_ (.A(_06703_),
    .B(_06548_),
    .Y(_06705_));
 sky130_fd_sc_hd__nand2_1 _17215_ (.A(_06388_),
    .B(_06479_),
    .Y(_06706_));
 sky130_fd_sc_hd__nand2_1 _17216_ (.A(_06705_),
    .B(_06706_),
    .Y(_06707_));
 sky130_fd_sc_hd__nand2_1 _17217_ (.A(_06707_),
    .B(_05915_),
    .Y(_06708_));
 sky130_fd_sc_hd__nand3_2 _17218_ (.A(_06705_),
    .B(_08834_),
    .C(_06706_),
    .Y(_06709_));
 sky130_fd_sc_hd__nand2_1 _17219_ (.A(_06708_),
    .B(_06709_),
    .Y(_06710_));
 sky130_fd_sc_hd__inv_4 _17220_ (.A(_06710_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_1 _17221_ (.A(_06700_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__nand2_1 _17222_ (.A(_06689_),
    .B(_06417_),
    .Y(_06713_));
 sky130_fd_sc_hd__nand2_1 _17223_ (.A(_06713_),
    .B(_06497_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand3_1 _17224_ (.A(_06689_),
    .B(_06496_),
    .C(_06417_),
    .Y(_06716_));
 sky130_fd_sc_hd__nand2_1 _17225_ (.A(_06714_),
    .B(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__nand2_1 _17226_ (.A(_06717_),
    .B(_06548_),
    .Y(_06718_));
 sky130_fd_sc_hd__nand2_1 _17227_ (.A(_06388_),
    .B(_06412_),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_1 _17228_ (.A(_06718_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__buf_6 _17229_ (.A(_09054_),
    .X(_06721_));
 sky130_fd_sc_hd__nand2_1 _17230_ (.A(_06720_),
    .B(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__clkbuf_8 _17231_ (.A(_09076_),
    .X(_06723_));
 sky130_fd_sc_hd__nand3_2 _17232_ (.A(_06718_),
    .B(_06723_),
    .C(_06719_),
    .Y(_06724_));
 sky130_fd_sc_hd__nand2_1 _17233_ (.A(_06722_),
    .B(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__or2_1 _17234_ (.A(_06424_),
    .B(_06548_),
    .X(_06727_));
 sky130_fd_sc_hd__nand3_1 _17235_ (.A(_06575_),
    .B(_06426_),
    .C(_06423_),
    .Y(_06728_));
 sky130_fd_sc_hd__nand3_1 _17236_ (.A(_06577_),
    .B(_06548_),
    .C(_06728_),
    .Y(_06729_));
 sky130_fd_sc_hd__nand2_1 _17237_ (.A(_06727_),
    .B(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__buf_6 _17238_ (.A(_08966_),
    .X(_06731_));
 sky130_fd_sc_hd__nand2_1 _17239_ (.A(_06730_),
    .B(_06731_),
    .Y(_06732_));
 sky130_fd_sc_hd__buf_4 _17240_ (.A(_08944_),
    .X(_06733_));
 sky130_fd_sc_hd__nand3_2 _17241_ (.A(_06727_),
    .B(_06729_),
    .C(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__nand2_2 _17242_ (.A(_06732_),
    .B(_06734_),
    .Y(_06735_));
 sky130_fd_sc_hd__nor2_1 _17243_ (.A(_06725_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__nor2b_1 _17244_ (.A(_06736_),
    .B_N(_06712_),
    .Y(_06738_));
 sky130_fd_sc_hd__nand2_1 _17245_ (.A(_06688_),
    .B(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__inv_2 _17246_ (.A(_06698_),
    .Y(_06740_));
 sky130_fd_sc_hd__o21ai_2 _17247_ (.A1(_06709_),
    .A2(_06740_),
    .B1(_06696_),
    .Y(_06741_));
 sky130_fd_sc_hd__inv_2 _17248_ (.A(_06734_),
    .Y(_06742_));
 sky130_fd_sc_hd__o21ai_1 _17249_ (.A1(_06724_),
    .A2(_06742_),
    .B1(_06732_),
    .Y(_06743_));
 sky130_fd_sc_hd__a21oi_1 _17250_ (.A1(_06736_),
    .A2(_06741_),
    .B1(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__nand2_2 _17251_ (.A(_06744_),
    .B(_06739_),
    .Y(_06745_));
 sky130_fd_sc_hd__nand2_1 _17252_ (.A(_06584_),
    .B(_06585_),
    .Y(_06746_));
 sky130_fd_sc_hd__nand2_1 _17253_ (.A(_06746_),
    .B(_06159_),
    .Y(_06747_));
 sky130_fd_sc_hd__nand2_1 _17254_ (.A(_06747_),
    .B(_06586_),
    .Y(_06749_));
 sky130_fd_sc_hd__nand2_1 _17255_ (.A(_06593_),
    .B(_06590_),
    .Y(_06750_));
 sky130_fd_sc_hd__nor2_1 _17256_ (.A(_06749_),
    .B(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__nand3_2 _17257_ (.A(_06745_),
    .B(_06574_),
    .C(_06751_),
    .Y(_06752_));
 sky130_fd_sc_hd__nand2_2 _17258_ (.A(_06598_),
    .B(_06752_),
    .Y(_06753_));
 sky130_fd_sc_hd__clkbuf_16 _17259_ (.A(_09361_),
    .X(_06754_));
 sky130_fd_sc_hd__inv_2 _17260_ (.A(_06261_),
    .Y(_06755_));
 sky130_fd_sc_hd__or2_1 _17261_ (.A(_06755_),
    .B(_06170_),
    .X(_06756_));
 sky130_fd_sc_hd__nand2_1 _17262_ (.A(_06170_),
    .B(_06755_),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_1 _17263_ (.A(_06756_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__inv_2 _17264_ (.A(_06758_),
    .Y(_06760_));
 sky130_fd_sc_hd__nand2_1 _17265_ (.A(_06760_),
    .B(_06207_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_1 _17266_ (.A(_06758_),
    .B(_05408_),
    .Y(_06762_));
 sky130_fd_sc_hd__nand2_1 _17267_ (.A(_06761_),
    .B(_06762_),
    .Y(_06763_));
 sky130_fd_sc_hd__inv_4 _17268_ (.A(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__nand2_1 _17269_ (.A(_06537_),
    .B(_06113_),
    .Y(_06765_));
 sky130_fd_sc_hd__inv_2 _17270_ (.A(_06141_),
    .Y(_06766_));
 sky130_fd_sc_hd__nand2_1 _17271_ (.A(_06765_),
    .B(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__nand3_1 _17272_ (.A(_06537_),
    .B(_06141_),
    .C(_06113_),
    .Y(_06768_));
 sky130_fd_sc_hd__nand2_1 _17273_ (.A(_06767_),
    .B(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__nand2_1 _17274_ (.A(_06769_),
    .B(_05375_),
    .Y(_06771_));
 sky130_fd_sc_hd__buf_6 _17275_ (.A(net39),
    .X(_06772_));
 sky130_fd_sc_hd__nand3_1 _17276_ (.A(_06767_),
    .B(_06772_),
    .C(_06768_),
    .Y(_06773_));
 sky130_fd_sc_hd__nand3_1 _17277_ (.A(_06545_),
    .B(_06771_),
    .C(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__inv_2 _17278_ (.A(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__nand3_1 _17279_ (.A(_06504_),
    .B(_06527_),
    .C(_06775_),
    .Y(_06776_));
 sky130_fd_sc_hd__inv_2 _17280_ (.A(_06771_),
    .Y(_06777_));
 sky130_fd_sc_hd__o21ai_1 _17281_ (.A1(_06542_),
    .A2(_06777_),
    .B1(_06773_),
    .Y(_06778_));
 sky130_fd_sc_hd__nor2_1 _17282_ (.A(_06531_),
    .B(_06774_),
    .Y(_06779_));
 sky130_fd_sc_hd__nor2_1 _17283_ (.A(_06778_),
    .B(_06779_),
    .Y(_06780_));
 sky130_fd_sc_hd__nand2_2 _17284_ (.A(_06776_),
    .B(_06780_),
    .Y(_06782_));
 sky130_fd_sc_hd__or2_1 _17285_ (.A(_06764_),
    .B(_06782_),
    .X(_06783_));
 sky130_fd_sc_hd__buf_6 _17286_ (.A(_06548_),
    .X(_06784_));
 sky130_fd_sc_hd__nand2_1 _17287_ (.A(_06782_),
    .B(_06764_),
    .Y(_06785_));
 sky130_fd_sc_hd__nand3_1 _17288_ (.A(_06783_),
    .B(_06784_),
    .C(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__nand2_1 _17289_ (.A(\div1i.quot[18] ),
    .B(_06760_),
    .Y(_06787_));
 sky130_fd_sc_hd__nand2_1 _17290_ (.A(_06786_),
    .B(_06787_),
    .Y(_06788_));
 sky130_fd_sc_hd__xor2_2 _17291_ (.A(_06754_),
    .B(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__nand2_1 _17292_ (.A(_06771_),
    .B(_06773_),
    .Y(_06790_));
 sky130_fd_sc_hd__nand2_1 _17293_ (.A(_06546_),
    .B(_06542_),
    .Y(_06791_));
 sky130_fd_sc_hd__xor2_1 _17294_ (.A(_06790_),
    .B(_06791_),
    .X(_06793_));
 sky130_fd_sc_hd__nand2_1 _17295_ (.A(_06793_),
    .B(_06548_),
    .Y(_06794_));
 sky130_fd_sc_hd__nand2_1 _17296_ (.A(\div1i.quot[18] ),
    .B(_06769_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand2_1 _17297_ (.A(_06794_),
    .B(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__buf_6 _17298_ (.A(_09548_),
    .X(_06797_));
 sky130_fd_sc_hd__nand2_1 _17299_ (.A(_06796_),
    .B(_06797_),
    .Y(_06798_));
 sky130_fd_sc_hd__buf_6 _17300_ (.A(_09559_),
    .X(_06799_));
 sky130_fd_sc_hd__nand3_1 _17301_ (.A(_06794_),
    .B(_06799_),
    .C(_06795_),
    .Y(_06800_));
 sky130_fd_sc_hd__nand2_1 _17302_ (.A(_06798_),
    .B(_06800_),
    .Y(_06801_));
 sky130_fd_sc_hd__nor2_1 _17303_ (.A(_06789_),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__nand2_1 _17304_ (.A(_06753_),
    .B(_06802_),
    .Y(_06804_));
 sky130_fd_sc_hd__buf_6 _17305_ (.A(_09383_),
    .X(_06805_));
 sky130_fd_sc_hd__nand2_1 _17306_ (.A(_06788_),
    .B(_06805_),
    .Y(_06806_));
 sky130_fd_sc_hd__o21a_1 _17307_ (.A1(_06800_),
    .A2(_06789_),
    .B1(_06806_),
    .X(_06807_));
 sky130_fd_sc_hd__nand2_1 _17308_ (.A(_06804_),
    .B(_06807_),
    .Y(_06808_));
 sky130_fd_sc_hd__buf_6 _17309_ (.A(_09987_),
    .X(_06809_));
 sky130_fd_sc_hd__inv_2 _17310_ (.A(_06242_),
    .Y(_06810_));
 sky130_fd_sc_hd__nand2_1 _17311_ (.A(_06170_),
    .B(_06262_),
    .Y(_06811_));
 sky130_fd_sc_hd__inv_2 _17312_ (.A(_06264_),
    .Y(_06812_));
 sky130_fd_sc_hd__nand2_1 _17313_ (.A(_06811_),
    .B(_06812_),
    .Y(_06813_));
 sky130_fd_sc_hd__or2_1 _17314_ (.A(_06810_),
    .B(_06813_),
    .X(_06815_));
 sky130_fd_sc_hd__nand2_1 _17315_ (.A(_06813_),
    .B(_06810_),
    .Y(_06816_));
 sky130_fd_sc_hd__nand2_1 _17316_ (.A(_06815_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__nand2_1 _17317_ (.A(_06817_),
    .B(_06737_),
    .Y(_06818_));
 sky130_fd_sc_hd__buf_6 _17318_ (.A(_06726_),
    .X(_06819_));
 sky130_fd_sc_hd__nand3_1 _17319_ (.A(_06815_),
    .B(_06819_),
    .C(_06816_),
    .Y(_06820_));
 sky130_fd_sc_hd__nand2_1 _17320_ (.A(_06818_),
    .B(_06820_),
    .Y(_06821_));
 sky130_fd_sc_hd__inv_2 _17321_ (.A(_06821_),
    .Y(_06822_));
 sky130_fd_sc_hd__nand2_1 _17322_ (.A(_06757_),
    .B(_06259_),
    .Y(_06823_));
 sky130_fd_sc_hd__xor2_2 _17323_ (.A(_06251_),
    .B(_06823_),
    .X(_06824_));
 sky130_fd_sc_hd__inv_2 _17324_ (.A(_06824_),
    .Y(_06826_));
 sky130_fd_sc_hd__buf_6 _17325_ (.A(net41),
    .X(_06827_));
 sky130_fd_sc_hd__nand2_1 _17326_ (.A(_06826_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__nand2_1 _17327_ (.A(_06824_),
    .B(_06814_),
    .Y(_06829_));
 sky130_fd_sc_hd__nand2_1 _17328_ (.A(_06828_),
    .B(_06829_),
    .Y(_06830_));
 sky130_fd_sc_hd__nand2b_1 _17329_ (.A_N(_06830_),
    .B(_06764_),
    .Y(_06831_));
 sky130_fd_sc_hd__inv_2 _17330_ (.A(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2_1 _17331_ (.A(_06782_),
    .B(_06832_),
    .Y(_06833_));
 sky130_fd_sc_hd__inv_2 _17332_ (.A(_06761_),
    .Y(_06834_));
 sky130_fd_sc_hd__a21boi_1 _17333_ (.A1(_06834_),
    .A2(_06829_),
    .B1_N(_06828_),
    .Y(_06835_));
 sky130_fd_sc_hd__nand2_1 _17334_ (.A(_06833_),
    .B(_06835_),
    .Y(_06837_));
 sky130_fd_sc_hd__or2_1 _17335_ (.A(_06822_),
    .B(_06837_),
    .X(_06838_));
 sky130_fd_sc_hd__nand2_1 _17336_ (.A(_06837_),
    .B(_06822_),
    .Y(_06839_));
 sky130_fd_sc_hd__nand3_1 _17337_ (.A(_06838_),
    .B(_06784_),
    .C(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__or2_1 _17338_ (.A(_06817_),
    .B(_06784_),
    .X(_06841_));
 sky130_fd_sc_hd__nand2_1 _17339_ (.A(_06840_),
    .B(_06841_),
    .Y(_06842_));
 sky130_fd_sc_hd__xor2_2 _17340_ (.A(_06809_),
    .B(_06842_),
    .X(_06843_));
 sky130_fd_sc_hd__buf_6 _17341_ (.A(_09735_),
    .X(_06844_));
 sky130_fd_sc_hd__nand2_1 _17342_ (.A(_06785_),
    .B(_06761_),
    .Y(_06845_));
 sky130_fd_sc_hd__xor2_1 _17343_ (.A(_06830_),
    .B(_06845_),
    .X(_06846_));
 sky130_fd_sc_hd__nand2_1 _17344_ (.A(_06846_),
    .B(_06784_),
    .Y(_06848_));
 sky130_fd_sc_hd__nand2_1 _17345_ (.A(\div1i.quot[18] ),
    .B(_06824_),
    .Y(_06849_));
 sky130_fd_sc_hd__nand2_1 _17346_ (.A(_06848_),
    .B(_06849_),
    .Y(_06850_));
 sky130_fd_sc_hd__or2_1 _17347_ (.A(_06844_),
    .B(_06850_),
    .X(_06851_));
 sky130_fd_sc_hd__nand2_1 _17348_ (.A(_06850_),
    .B(_06844_),
    .Y(_06852_));
 sky130_fd_sc_hd__nand2_1 _17349_ (.A(_06851_),
    .B(_06852_),
    .Y(_06853_));
 sky130_fd_sc_hd__nor2_1 _17350_ (.A(_06843_),
    .B(_06853_),
    .Y(_06854_));
 sky130_fd_sc_hd__nand2_1 _17351_ (.A(_06808_),
    .B(_06854_),
    .Y(_06855_));
 sky130_fd_sc_hd__buf_6 _17352_ (.A(net241),
    .X(_06856_));
 sky130_fd_sc_hd__nand2_1 _17353_ (.A(_06842_),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__o21a_1 _17354_ (.A1(_06851_),
    .A2(_06843_),
    .B1(_06857_),
    .X(_06859_));
 sky130_fd_sc_hd__nand2_2 _17355_ (.A(_06855_),
    .B(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__or2_1 _17356_ (.A(_06341_),
    .B(net139),
    .X(_06861_));
 sky130_fd_sc_hd__nand2_1 _17357_ (.A(net139),
    .B(_06341_),
    .Y(_06862_));
 sky130_fd_sc_hd__nand2_1 _17358_ (.A(_06861_),
    .B(_06862_),
    .Y(_06863_));
 sky130_fd_sc_hd__or2_1 _17359_ (.A(_10426_),
    .B(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__nand2_1 _17360_ (.A(_06863_),
    .B(_10426_),
    .Y(_06865_));
 sky130_fd_sc_hd__nand2_1 _17361_ (.A(_06864_),
    .B(_06865_),
    .Y(_06866_));
 sky130_fd_sc_hd__nand2_1 _17362_ (.A(_06816_),
    .B(_06240_),
    .Y(_06867_));
 sky130_fd_sc_hd__nand2b_1 _17363_ (.A_N(_06867_),
    .B(_06231_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand3_1 _17364_ (.A(_06867_),
    .B(_06230_),
    .C(_06229_),
    .Y(_06870_));
 sky130_fd_sc_hd__nand2_1 _17365_ (.A(_06868_),
    .B(_06870_),
    .Y(_06871_));
 sky130_fd_sc_hd__nand2_1 _17366_ (.A(_06871_),
    .B(_06704_),
    .Y(_06872_));
 sky130_fd_sc_hd__inv_2 _17367_ (.A(_06820_),
    .Y(_06873_));
 sky130_fd_sc_hd__buf_6 _17368_ (.A(net43),
    .X(_06874_));
 sky130_fd_sc_hd__nand3_2 _17369_ (.A(_06868_),
    .B(_06874_),
    .C(_06870_),
    .Y(_06875_));
 sky130_fd_sc_hd__inv_2 _17370_ (.A(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__a21o_1 _17371_ (.A1(_06872_),
    .A2(_06873_),
    .B1(_06876_),
    .X(_06877_));
 sky130_fd_sc_hd__nand3_1 _17372_ (.A(_06872_),
    .B(_06822_),
    .C(_06875_),
    .Y(_06878_));
 sky130_fd_sc_hd__nor2_1 _17373_ (.A(_06835_),
    .B(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__nor2_1 _17374_ (.A(_06877_),
    .B(_06879_),
    .Y(_06881_));
 sky130_fd_sc_hd__inv_2 _17375_ (.A(_06878_),
    .Y(_06882_));
 sky130_fd_sc_hd__nand3_1 _17376_ (.A(_06782_),
    .B(_06882_),
    .C(_06832_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_1 _17377_ (.A(_06881_),
    .B(_06883_),
    .Y(_06884_));
 sky130_fd_sc_hd__xor2_1 _17378_ (.A(_06866_),
    .B(_06884_),
    .X(_06885_));
 sky130_fd_sc_hd__nand2_1 _17379_ (.A(_06885_),
    .B(_06784_),
    .Y(_06886_));
 sky130_fd_sc_hd__nand2_1 _17380_ (.A(\div1i.quot[18] ),
    .B(_06863_),
    .Y(_06887_));
 sky130_fd_sc_hd__nand2_1 _17381_ (.A(_06886_),
    .B(_06887_),
    .Y(_06888_));
 sky130_fd_sc_hd__nand2_1 _17382_ (.A(_06888_),
    .B(_10481_),
    .Y(_06889_));
 sky130_fd_sc_hd__nand3_1 _17383_ (.A(_06886_),
    .B(_06348_),
    .C(_06887_),
    .Y(_06890_));
 sky130_fd_sc_hd__nand2_2 _17384_ (.A(_06889_),
    .B(_06890_),
    .Y(_06892_));
 sky130_fd_sc_hd__inv_2 _17385_ (.A(_06892_),
    .Y(_06893_));
 sky130_fd_sc_hd__nand2_1 _17386_ (.A(_06872_),
    .B(_06875_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand2_1 _17387_ (.A(_06839_),
    .B(_06820_),
    .Y(_06895_));
 sky130_fd_sc_hd__xor2_1 _17388_ (.A(_06894_),
    .B(_06895_),
    .X(_06896_));
 sky130_fd_sc_hd__nand2_1 _17389_ (.A(_06896_),
    .B(_06784_),
    .Y(_06897_));
 sky130_fd_sc_hd__clkbuf_8 _17390_ (.A(_10240_),
    .X(_06898_));
 sky130_fd_sc_hd__nand2_1 _17391_ (.A(_06871_),
    .B(\div1i.quot[18] ),
    .Y(_06899_));
 sky130_fd_sc_hd__nand3_2 _17392_ (.A(_06897_),
    .B(_06898_),
    .C(_06899_),
    .Y(_06900_));
 sky130_fd_sc_hd__nand2_1 _17393_ (.A(_06897_),
    .B(_06899_),
    .Y(_06901_));
 sky130_fd_sc_hd__buf_4 _17394_ (.A(_10251_),
    .X(_06903_));
 sky130_fd_sc_hd__nand2_1 _17395_ (.A(_06901_),
    .B(_06903_),
    .Y(_06904_));
 sky130_fd_sc_hd__nand3_1 _17396_ (.A(_06893_),
    .B(_06900_),
    .C(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__inv_2 _17397_ (.A(_06866_),
    .Y(_06906_));
 sky130_fd_sc_hd__nand2_1 _17398_ (.A(_06884_),
    .B(_06906_),
    .Y(_06907_));
 sky130_fd_sc_hd__nand2_1 _17399_ (.A(_06907_),
    .B(_06864_),
    .Y(_06908_));
 sky130_fd_sc_hd__nand2_2 _17400_ (.A(_06862_),
    .B(_06339_),
    .Y(_06909_));
 sky130_fd_sc_hd__xor2_2 _17401_ (.A(_06351_),
    .B(_06909_),
    .X(_06910_));
 sky130_fd_sc_hd__or2_4 _17402_ (.A(_06550_),
    .B(_06910_),
    .X(_06911_));
 sky130_fd_sc_hd__nand2_1 _17403_ (.A(_06910_),
    .B(_06550_),
    .Y(_06912_));
 sky130_fd_sc_hd__nand2_2 _17404_ (.A(_06911_),
    .B(_06912_),
    .Y(_06914_));
 sky130_fd_sc_hd__inv_2 _17405_ (.A(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__nand2_1 _17406_ (.A(_06908_),
    .B(_06915_),
    .Y(_06916_));
 sky130_fd_sc_hd__nand3_1 _17407_ (.A(_06907_),
    .B(_06914_),
    .C(_06864_),
    .Y(_06917_));
 sky130_fd_sc_hd__nand2_1 _17408_ (.A(_06916_),
    .B(_06917_),
    .Y(_06918_));
 sky130_fd_sc_hd__nand2_1 _17409_ (.A(_06918_),
    .B(_06784_),
    .Y(_06919_));
 sky130_fd_sc_hd__nand2_1 _17410_ (.A(_06910_),
    .B(\div1i.quot[18] ),
    .Y(_06920_));
 sky130_fd_sc_hd__nand2_1 _17411_ (.A(_06919_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__nand2_1 _17412_ (.A(_06921_),
    .B(_10701_),
    .Y(_06922_));
 sky130_fd_sc_hd__nand3_2 _17413_ (.A(_06919_),
    .B(_06366_),
    .C(_06920_),
    .Y(_06923_));
 sky130_fd_sc_hd__nand2_1 _17414_ (.A(_06922_),
    .B(_06923_),
    .Y(_06925_));
 sky130_fd_sc_hd__inv_2 _17415_ (.A(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__nand2_1 _17416_ (.A(_06915_),
    .B(_06906_),
    .Y(_06927_));
 sky130_fd_sc_hd__inv_2 _17417_ (.A(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _17418_ (.A(_06884_),
    .B(_06928_),
    .Y(_06929_));
 sky130_fd_sc_hd__o21a_1 _17419_ (.A1(_06864_),
    .A2(_06914_),
    .B1(_06911_),
    .X(_06930_));
 sky130_fd_sc_hd__nand2_1 _17420_ (.A(_06929_),
    .B(_06930_),
    .Y(_06931_));
 sky130_fd_sc_hd__a31o_1 _17421_ (.A1(net139),
    .A2(_06352_),
    .A3(_06341_),
    .B1(_06372_),
    .X(_06932_));
 sky130_fd_sc_hd__xor2_1 _17422_ (.A(_06368_),
    .B(_06932_),
    .X(_06933_));
 sky130_fd_sc_hd__inv_2 _17423_ (.A(_06933_),
    .Y(_06934_));
 sky130_fd_sc_hd__buf_6 _17424_ (.A(net47),
    .X(_06936_));
 sky130_fd_sc_hd__nand2_1 _17425_ (.A(_06934_),
    .B(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__nand2_1 _17426_ (.A(_06933_),
    .B(_06594_),
    .Y(_06938_));
 sky130_fd_sc_hd__nand2_1 _17427_ (.A(_06937_),
    .B(_06938_),
    .Y(_06939_));
 sky130_fd_sc_hd__inv_2 _17428_ (.A(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__nand2_2 _17429_ (.A(_06931_),
    .B(_06940_),
    .Y(_06941_));
 sky130_fd_sc_hd__nand3_1 _17430_ (.A(_06929_),
    .B(_06930_),
    .C(_06939_),
    .Y(_06942_));
 sky130_fd_sc_hd__nand3_2 _17431_ (.A(_06941_),
    .B(_06784_),
    .C(_06942_),
    .Y(_06943_));
 sky130_fd_sc_hd__nand2_1 _17432_ (.A(_06934_),
    .B(\div1i.quot[18] ),
    .Y(_06944_));
 sky130_fd_sc_hd__nand2_1 _17433_ (.A(_06943_),
    .B(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__buf_6 _17434_ (.A(_10887_),
    .X(_06947_));
 sky130_fd_sc_hd__nand2_2 _17435_ (.A(_06945_),
    .B(_06947_),
    .Y(_06948_));
 sky130_fd_sc_hd__buf_6 _17436_ (.A(_10909_),
    .X(_06949_));
 sky130_fd_sc_hd__nand3_2 _17437_ (.A(_06943_),
    .B(_06949_),
    .C(_06944_),
    .Y(_06950_));
 sky130_fd_sc_hd__nand2_4 _17438_ (.A(_06948_),
    .B(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__inv_2 _17439_ (.A(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__nand2_1 _17440_ (.A(_06926_),
    .B(_06952_),
    .Y(_06953_));
 sky130_fd_sc_hd__nor2_1 _17441_ (.A(_06905_),
    .B(_06953_),
    .Y(_06954_));
 sky130_fd_sc_hd__nand2_4 _17442_ (.A(_06860_),
    .B(_06954_),
    .Y(_06955_));
 sky130_fd_sc_hd__inv_2 _17443_ (.A(_06889_),
    .Y(_06956_));
 sky130_fd_sc_hd__o21ai_1 _17444_ (.A1(_06956_),
    .A2(_06900_),
    .B1(_06890_),
    .Y(_06958_));
 sky130_fd_sc_hd__nor2_1 _17445_ (.A(_06951_),
    .B(_06925_),
    .Y(_06959_));
 sky130_fd_sc_hd__o21ai_1 _17446_ (.A1(_06923_),
    .A2(_06951_),
    .B1(_06948_),
    .Y(_06960_));
 sky130_fd_sc_hd__a21oi_2 _17447_ (.A1(_06958_),
    .A2(_06959_),
    .B1(_06960_),
    .Y(_06961_));
 sky130_fd_sc_hd__nand2_4 _17448_ (.A(_06955_),
    .B(_06961_),
    .Y(_06962_));
 sky130_fd_sc_hd__a21bo_1 _17449_ (.A1(_06932_),
    .A2(_06365_),
    .B1_N(_06367_),
    .X(_06963_));
 sky130_fd_sc_hd__xor2_4 _17450_ (.A(_06327_),
    .B(_06963_),
    .X(_06964_));
 sky130_fd_sc_hd__nand3_2 _17451_ (.A(_06941_),
    .B(_06784_),
    .C(_06937_),
    .Y(_06965_));
 sky130_fd_sc_hd__xor2_4 _17452_ (.A(_06964_),
    .B(_06965_),
    .X(_06966_));
 sky130_fd_sc_hd__clkinvlp_2 _17453_ (.A(_06966_),
    .Y(_06967_));
 sky130_fd_sc_hd__nand2_8 _17454_ (.A(_06962_),
    .B(_06967_),
    .Y(_06969_));
 sky130_fd_sc_hd__nand3_4 _17455_ (.A(_06955_),
    .B(_06961_),
    .C(_06966_),
    .Y(_06970_));
 sky130_fd_sc_hd__nand2_8 _17456_ (.A(_06969_),
    .B(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__buf_8 _17457_ (.A(_06971_),
    .X(_06972_));
 sky130_fd_sc_hd__buf_12 _17458_ (.A(net157),
    .X(\div1i.quot[17] ));
 sky130_fd_sc_hd__nand2_1 _17459_ (.A(_06617_),
    .B(_06621_),
    .Y(_06973_));
 sky130_fd_sc_hd__nand2_1 _17460_ (.A(_06973_),
    .B(_06622_),
    .Y(_06974_));
 sky130_fd_sc_hd__nand2_1 _17461_ (.A(_06974_),
    .B(net237),
    .Y(_06975_));
 sky130_fd_sc_hd__inv_2 _17462_ (.A(_06975_),
    .Y(_06976_));
 sky130_fd_sc_hd__nand2_1 _17463_ (.A(_06972_),
    .B(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__buf_6 _17464_ (.A(_05496_),
    .X(_06979_));
 sky130_fd_sc_hd__buf_6 _17465_ (.A(_05474_),
    .X(_06980_));
 sky130_fd_sc_hd__o21ai_2 _17466_ (.A1(_06979_),
    .A2(\div1i.quot[18] ),
    .B1(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__buf_6 _17467_ (.A(_05189_),
    .X(_06982_));
 sky130_fd_sc_hd__nand2_1 _17468_ (.A(_06975_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__buf_6 _17469_ (.A(net55),
    .X(_06984_));
 sky130_fd_sc_hd__nand3_1 _17470_ (.A(_06974_),
    .B(_06984_),
    .C(_06624_),
    .Y(_06985_));
 sky130_fd_sc_hd__nand2_1 _17471_ (.A(_06983_),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__xor2_1 _17472_ (.A(_06981_),
    .B(_06986_),
    .X(_06987_));
 sky130_fd_sc_hd__nand3b_1 _17473_ (.A_N(_06987_),
    .B(net127),
    .C(_06970_),
    .Y(_06988_));
 sky130_fd_sc_hd__nand2_1 _17474_ (.A(_06977_),
    .B(_06988_),
    .Y(_06990_));
 sky130_fd_sc_hd__nand2_1 _17475_ (.A(_06990_),
    .B(_05983_),
    .Y(_06991_));
 sky130_fd_sc_hd__nor2_1 _17476_ (.A(_06979_),
    .B(_06784_),
    .Y(_06992_));
 sky130_fd_sc_hd__or2_1 _17477_ (.A(_06607_),
    .B(_06992_),
    .X(_06993_));
 sky130_fd_sc_hd__nand2_1 _17478_ (.A(_06993_),
    .B(_06622_),
    .Y(_06994_));
 sky130_fd_sc_hd__inv_2 _17479_ (.A(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__nand2_1 _17480_ (.A(_06972_),
    .B(_06995_),
    .Y(_06996_));
 sky130_fd_sc_hd__nand3_1 _17481_ (.A(net126),
    .B(_06970_),
    .C(_06992_),
    .Y(_06997_));
 sky130_fd_sc_hd__nand2_1 _17482_ (.A(_06996_),
    .B(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__nand2_2 _17483_ (.A(_06998_),
    .B(_06615_),
    .Y(_06999_));
 sky130_fd_sc_hd__nand2_1 _17484_ (.A(_06991_),
    .B(_06999_),
    .Y(_07001_));
 sky130_fd_sc_hd__inv_2 _17485_ (.A(_07001_),
    .Y(_07002_));
 sky130_fd_sc_hd__nand3_1 _17486_ (.A(_06996_),
    .B(_06620_),
    .C(_06997_),
    .Y(_07003_));
 sky130_fd_sc_hd__buf_6 _17487_ (.A(_07308_),
    .X(_07004_));
 sky130_fd_sc_hd__nand3_2 _17488_ (.A(_06972_),
    .B(_06980_),
    .C(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__inv_2 _17489_ (.A(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__nand3_2 _17490_ (.A(_06999_),
    .B(_07003_),
    .C(_07006_),
    .Y(_07007_));
 sky130_fd_sc_hd__or2_4 _17491_ (.A(_05983_),
    .B(_06990_),
    .X(_07008_));
 sky130_fd_sc_hd__inv_2 _17492_ (.A(_07008_),
    .Y(_07009_));
 sky130_fd_sc_hd__a21oi_2 _17493_ (.A1(_07002_),
    .A2(_07007_),
    .B1(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__nand2_1 _17494_ (.A(_06619_),
    .B(_06624_),
    .Y(_07012_));
 sky130_fd_sc_hd__nand2_1 _17495_ (.A(_07012_),
    .B(_06625_),
    .Y(_07013_));
 sky130_fd_sc_hd__clkinvlp_2 _17496_ (.A(_06683_),
    .Y(_07014_));
 sky130_fd_sc_hd__o21ai_1 _17497_ (.A1(_06678_),
    .A2(_07013_),
    .B1(_07014_),
    .Y(_07015_));
 sky130_fd_sc_hd__or2_1 _17498_ (.A(_06654_),
    .B(_07015_),
    .X(_07016_));
 sky130_fd_sc_hd__nand2_1 _17499_ (.A(_07015_),
    .B(_06654_),
    .Y(_07017_));
 sky130_fd_sc_hd__nand2_1 _17500_ (.A(_07016_),
    .B(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__inv_2 _17501_ (.A(_07018_),
    .Y(_07019_));
 sky130_fd_sc_hd__nand2_1 _17502_ (.A(net161),
    .B(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__buf_6 _17503_ (.A(net61),
    .X(_07021_));
 sky130_fd_sc_hd__nand2_1 _17504_ (.A(_07019_),
    .B(_07021_),
    .Y(_07023_));
 sky130_fd_sc_hd__buf_4 _17505_ (.A(_05847_),
    .X(_07024_));
 sky130_fd_sc_hd__nand2_1 _17506_ (.A(_07018_),
    .B(_07024_),
    .Y(_07025_));
 sky130_fd_sc_hd__nand2_1 _17507_ (.A(_07023_),
    .B(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__inv_2 _17508_ (.A(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__nand2_1 _17509_ (.A(_06626_),
    .B(_06677_),
    .Y(_07028_));
 sky130_fd_sc_hd__nand2_1 _17510_ (.A(_07013_),
    .B(_06676_),
    .Y(_07029_));
 sky130_fd_sc_hd__nand2_1 _17511_ (.A(_07028_),
    .B(_07029_),
    .Y(_07030_));
 sky130_fd_sc_hd__buf_6 _17512_ (.A(_05705_),
    .X(_07031_));
 sky130_fd_sc_hd__nand2_1 _17513_ (.A(_07030_),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__buf_6 _17514_ (.A(net59),
    .X(_07034_));
 sky130_fd_sc_hd__nand3_1 _17515_ (.A(_07028_),
    .B(_07034_),
    .C(_07029_),
    .Y(_07035_));
 sky130_fd_sc_hd__nand2_1 _17516_ (.A(_07032_),
    .B(_07035_),
    .Y(_07036_));
 sky130_fd_sc_hd__inv_2 _17517_ (.A(_07036_),
    .Y(_07037_));
 sky130_fd_sc_hd__inv_2 _17518_ (.A(_06985_),
    .Y(_07038_));
 sky130_fd_sc_hd__a21o_1 _17519_ (.A1(_06983_),
    .A2(_06981_),
    .B1(_07038_),
    .X(_07039_));
 sky130_fd_sc_hd__nand2_1 _17520_ (.A(_06625_),
    .B(_06606_),
    .Y(_07040_));
 sky130_fd_sc_hd__nand2_1 _17521_ (.A(_06624_),
    .B(_06617_),
    .Y(_07041_));
 sky130_fd_sc_hd__xor2_1 _17522_ (.A(_07040_),
    .B(_07041_),
    .X(_07042_));
 sky130_fd_sc_hd__buf_4 _17523_ (.A(_05178_),
    .X(_07043_));
 sky130_fd_sc_hd__nand2_1 _17524_ (.A(_07042_),
    .B(_07043_),
    .Y(_07045_));
 sky130_fd_sc_hd__nand2_1 _17525_ (.A(_07039_),
    .B(_07045_),
    .Y(_07046_));
 sky130_fd_sc_hd__inv_2 _17526_ (.A(_07042_),
    .Y(_07047_));
 sky130_fd_sc_hd__buf_6 _17527_ (.A(net58),
    .X(_07048_));
 sky130_fd_sc_hd__nand2_1 _17528_ (.A(_07047_),
    .B(_07048_),
    .Y(_07049_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_07046_),
    .B(_07049_),
    .Y(_07050_));
 sky130_fd_sc_hd__nand2_1 _17530_ (.A(_07037_),
    .B(_07050_),
    .Y(_07051_));
 sky130_fd_sc_hd__nand2_1 _17531_ (.A(_07051_),
    .B(_07035_),
    .Y(_07052_));
 sky130_fd_sc_hd__nand2_1 _17532_ (.A(_07028_),
    .B(_06674_),
    .Y(_07053_));
 sky130_fd_sc_hd__xor2_1 _17533_ (.A(_06666_),
    .B(_07053_),
    .X(_07054_));
 sky130_fd_sc_hd__nand2_1 _17534_ (.A(_07054_),
    .B(_06465_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand2_1 _17535_ (.A(_07052_),
    .B(_07056_),
    .Y(_07057_));
 sky130_fd_sc_hd__inv_2 _17536_ (.A(_07054_),
    .Y(_07058_));
 sky130_fd_sc_hd__nand2_1 _17537_ (.A(_07058_),
    .B(_05211_),
    .Y(_07059_));
 sky130_fd_sc_hd__nand2_1 _17538_ (.A(_07057_),
    .B(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__or2_1 _17539_ (.A(_07027_),
    .B(_07060_),
    .X(_07061_));
 sky130_fd_sc_hd__nand2_2 _17540_ (.A(_07060_),
    .B(_07027_),
    .Y(_07062_));
 sky130_fd_sc_hd__nand2_1 _17541_ (.A(_07061_),
    .B(_07062_),
    .Y(_07063_));
 sky130_fd_sc_hd__inv_2 _17542_ (.A(_07063_),
    .Y(_07064_));
 sky130_fd_sc_hd__nand3_1 _17543_ (.A(net125),
    .B(_06970_),
    .C(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__nand2_1 _17544_ (.A(_07020_),
    .B(_07065_),
    .Y(_07067_));
 sky130_fd_sc_hd__nand2_2 _17545_ (.A(_07067_),
    .B(_06636_),
    .Y(_07068_));
 sky130_fd_sc_hd__nand3_2 _17546_ (.A(_07020_),
    .B(_06639_),
    .C(_07065_),
    .Y(_07069_));
 sky130_fd_sc_hd__nand2_2 _17547_ (.A(_07068_),
    .B(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__inv_2 _17548_ (.A(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__nand2_1 _17549_ (.A(_06971_),
    .B(_07058_),
    .Y(_07072_));
 sky130_fd_sc_hd__nand2_1 _17550_ (.A(_07059_),
    .B(_07056_),
    .Y(_07073_));
 sky130_fd_sc_hd__xnor2_1 _17551_ (.A(_07052_),
    .B(_07073_),
    .Y(_07074_));
 sky130_fd_sc_hd__nand3_1 _17552_ (.A(_06969_),
    .B(_06970_),
    .C(_07074_),
    .Y(_07075_));
 sky130_fd_sc_hd__nand2_1 _17553_ (.A(_07072_),
    .B(_07075_),
    .Y(_07076_));
 sky130_fd_sc_hd__nand2_2 _17554_ (.A(_07076_),
    .B(_06651_),
    .Y(_07078_));
 sky130_fd_sc_hd__nand3_1 _17555_ (.A(_07072_),
    .B(_06648_),
    .C(_07075_),
    .Y(_07079_));
 sky130_fd_sc_hd__nand2_1 _17556_ (.A(_07078_),
    .B(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__inv_2 _17557_ (.A(_07080_),
    .Y(_07081_));
 sky130_fd_sc_hd__nand2_1 _17558_ (.A(_07071_),
    .B(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__inv_2 _17559_ (.A(_07030_),
    .Y(_07083_));
 sky130_fd_sc_hd__nand2_1 _17560_ (.A(_06971_),
    .B(_07083_),
    .Y(_07084_));
 sky130_fd_sc_hd__or2_1 _17561_ (.A(_07050_),
    .B(_07037_),
    .X(_07085_));
 sky130_fd_sc_hd__nand2_1 _17562_ (.A(_07085_),
    .B(_07051_),
    .Y(_07086_));
 sky130_fd_sc_hd__clkinvlp_2 _17563_ (.A(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__nand3_1 _17564_ (.A(net124),
    .B(_06970_),
    .C(_07087_),
    .Y(_07089_));
 sky130_fd_sc_hd__nand2_1 _17565_ (.A(_07084_),
    .B(_07089_),
    .Y(_07090_));
 sky130_fd_sc_hd__nand2_1 _17566_ (.A(_07090_),
    .B(_06033_),
    .Y(_07091_));
 sky130_fd_sc_hd__buf_6 _17567_ (.A(_12051_),
    .X(_07092_));
 sky130_fd_sc_hd__nand3_1 _17568_ (.A(_07084_),
    .B(_07092_),
    .C(_07089_),
    .Y(_07093_));
 sky130_fd_sc_hd__nand2_2 _17569_ (.A(_07091_),
    .B(_07093_),
    .Y(_07094_));
 sky130_fd_sc_hd__inv_2 _17570_ (.A(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__nand2_1 _17571_ (.A(_06971_),
    .B(_07047_),
    .Y(_07096_));
 sky130_fd_sc_hd__nand2_1 _17572_ (.A(_07049_),
    .B(_07045_),
    .Y(_07097_));
 sky130_fd_sc_hd__xnor2_1 _17573_ (.A(_07039_),
    .B(_07097_),
    .Y(_07098_));
 sky130_fd_sc_hd__nand3_1 _17574_ (.A(net123),
    .B(_06970_),
    .C(_07098_),
    .Y(_07100_));
 sky130_fd_sc_hd__nand2_1 _17575_ (.A(_07096_),
    .B(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__buf_6 _17576_ (.A(_07725_),
    .X(_07102_));
 sky130_fd_sc_hd__nand2_1 _17577_ (.A(_07101_),
    .B(_07102_),
    .Y(_07103_));
 sky130_fd_sc_hd__nand3_1 _17578_ (.A(_07096_),
    .B(_06046_),
    .C(_07100_),
    .Y(_07104_));
 sky130_fd_sc_hd__nand2_2 _17579_ (.A(_07103_),
    .B(_07104_),
    .Y(_07105_));
 sky130_fd_sc_hd__inv_2 _17580_ (.A(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__nand2_1 _17581_ (.A(_07095_),
    .B(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__nor2_1 _17582_ (.A(_07082_),
    .B(_07107_),
    .Y(_07108_));
 sky130_fd_sc_hd__nand2_1 _17583_ (.A(_07010_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__inv_2 _17584_ (.A(_07093_),
    .Y(_07111_));
 sky130_fd_sc_hd__o21ai_2 _17585_ (.A1(_07103_),
    .A2(_07111_),
    .B1(_07091_),
    .Y(_07112_));
 sky130_fd_sc_hd__nor2_1 _17586_ (.A(_07070_),
    .B(_07080_),
    .Y(_07113_));
 sky130_fd_sc_hd__inv_2 _17587_ (.A(_07069_),
    .Y(_07114_));
 sky130_fd_sc_hd__o21ai_1 _17588_ (.A1(_07078_),
    .A2(_07114_),
    .B1(_07068_),
    .Y(_07115_));
 sky130_fd_sc_hd__a21oi_1 _17589_ (.A1(_07112_),
    .A2(_07113_),
    .B1(_07115_),
    .Y(_07116_));
 sky130_fd_sc_hd__nand2_2 _17590_ (.A(_07116_),
    .B(_07109_),
    .Y(_07117_));
 sky130_fd_sc_hd__inv_2 _17591_ (.A(_06712_),
    .Y(_07118_));
 sky130_fd_sc_hd__nand2_1 _17592_ (.A(_06688_),
    .B(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__inv_2 _17593_ (.A(_06741_),
    .Y(_07120_));
 sky130_fd_sc_hd__nand2_1 _17594_ (.A(_07119_),
    .B(_07120_),
    .Y(_07122_));
 sky130_fd_sc_hd__inv_2 _17595_ (.A(_06725_),
    .Y(_07123_));
 sky130_fd_sc_hd__nand2_1 _17596_ (.A(_07122_),
    .B(_07123_),
    .Y(_07124_));
 sky130_fd_sc_hd__nand3_1 _17597_ (.A(_07119_),
    .B(_06725_),
    .C(_07120_),
    .Y(_07125_));
 sky130_fd_sc_hd__nand2_1 _17598_ (.A(_07124_),
    .B(_07125_),
    .Y(_07126_));
 sky130_fd_sc_hd__inv_2 _17599_ (.A(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__buf_6 _17600_ (.A(net34),
    .X(_07128_));
 sky130_fd_sc_hd__nand2_1 _17601_ (.A(_07127_),
    .B(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__buf_6 _17602_ (.A(_05299_),
    .X(_07130_));
 sky130_fd_sc_hd__nand2_1 _17603_ (.A(_07126_),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__nand2_1 _17604_ (.A(_07129_),
    .B(_07131_),
    .Y(_07133_));
 sky130_fd_sc_hd__inv_2 _17605_ (.A(_07133_),
    .Y(_07134_));
 sky130_fd_sc_hd__nand2_1 _17606_ (.A(_07017_),
    .B(_06652_),
    .Y(_07135_));
 sky130_fd_sc_hd__or2_1 _17607_ (.A(_06642_),
    .B(_07135_),
    .X(_07136_));
 sky130_fd_sc_hd__nand2_1 _17608_ (.A(_07135_),
    .B(_06642_),
    .Y(_07137_));
 sky130_fd_sc_hd__nand3_1 _17609_ (.A(_07136_),
    .B(_05896_),
    .C(_07137_),
    .Y(_07138_));
 sky130_fd_sc_hd__nand2_1 _17610_ (.A(_07138_),
    .B(_07023_),
    .Y(_07139_));
 sky130_fd_sc_hd__inv_2 _17611_ (.A(_07139_),
    .Y(_07140_));
 sky130_fd_sc_hd__nand2_2 _17612_ (.A(_07062_),
    .B(_07140_),
    .Y(_07141_));
 sky130_fd_sc_hd__nand2_2 _17613_ (.A(_06688_),
    .B(_06711_),
    .Y(_07142_));
 sky130_fd_sc_hd__nand2_2 _17614_ (.A(_07142_),
    .B(_06709_),
    .Y(_07144_));
 sky130_fd_sc_hd__xor2_1 _17615_ (.A(_06699_),
    .B(_07144_),
    .X(_07145_));
 sky130_fd_sc_hd__buf_6 _17616_ (.A(_05310_),
    .X(_07146_));
 sky130_fd_sc_hd__nand2_1 _17617_ (.A(_07145_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__or2_1 _17618_ (.A(_06700_),
    .B(_07144_),
    .X(_07148_));
 sky130_fd_sc_hd__buf_6 _17619_ (.A(net64),
    .X(_07149_));
 sky130_fd_sc_hd__nand2_1 _17620_ (.A(_07144_),
    .B(_06700_),
    .Y(_07150_));
 sky130_fd_sc_hd__nand3_1 _17621_ (.A(_07148_),
    .B(_07149_),
    .C(_07150_),
    .Y(_07151_));
 sky130_fd_sc_hd__or2_1 _17622_ (.A(_06711_),
    .B(_06688_),
    .X(_07152_));
 sky130_fd_sc_hd__nand2_1 _17623_ (.A(_07152_),
    .B(_07142_),
    .Y(_07153_));
 sky130_fd_sc_hd__buf_6 _17624_ (.A(_05321_),
    .X(_07155_));
 sky130_fd_sc_hd__nand2_1 _17625_ (.A(_07153_),
    .B(_07155_),
    .Y(_07156_));
 sky130_fd_sc_hd__buf_6 _17626_ (.A(net63),
    .X(_07157_));
 sky130_fd_sc_hd__nand3_2 _17627_ (.A(_07152_),
    .B(_07157_),
    .C(_07142_),
    .Y(_07158_));
 sky130_fd_sc_hd__nand2_1 _17628_ (.A(_07156_),
    .B(_07158_),
    .Y(_07159_));
 sky130_fd_sc_hd__inv_2 _17629_ (.A(_07159_),
    .Y(_07160_));
 sky130_fd_sc_hd__nand3_1 _17630_ (.A(_07147_),
    .B(_07151_),
    .C(_07160_),
    .Y(_07161_));
 sky130_fd_sc_hd__inv_2 _17631_ (.A(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__nand2_1 _17632_ (.A(_07136_),
    .B(_07137_),
    .Y(_07163_));
 sky130_fd_sc_hd__nand2_1 _17633_ (.A(_07163_),
    .B(_05255_),
    .Y(_07164_));
 sky130_fd_sc_hd__nand3_2 _17634_ (.A(_07141_),
    .B(_07162_),
    .C(_07164_),
    .Y(_07166_));
 sky130_fd_sc_hd__inv_2 _17635_ (.A(_07158_),
    .Y(_07167_));
 sky130_fd_sc_hd__a21boi_2 _17636_ (.A1(_07147_),
    .A2(_07167_),
    .B1_N(_07151_),
    .Y(_07168_));
 sky130_fd_sc_hd__nand2_1 _17637_ (.A(_07166_),
    .B(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__or2_1 _17638_ (.A(_07134_),
    .B(_07169_),
    .X(_07170_));
 sky130_fd_sc_hd__inv_6 _17639_ (.A(net161),
    .Y(_07171_));
 sky130_fd_sc_hd__nand2_1 _17640_ (.A(_07169_),
    .B(_07134_),
    .Y(_07172_));
 sky130_fd_sc_hd__nand3_1 _17641_ (.A(_07170_),
    .B(_07171_),
    .C(_07172_),
    .Y(_07173_));
 sky130_fd_sc_hd__nand2_1 _17642_ (.A(net157),
    .B(_07127_),
    .Y(_07174_));
 sky130_fd_sc_hd__nand2_1 _17643_ (.A(_07173_),
    .B(_07174_),
    .Y(_07175_));
 sky130_fd_sc_hd__nand2_1 _17644_ (.A(_07175_),
    .B(_06731_),
    .Y(_07177_));
 sky130_fd_sc_hd__nand3_1 _17645_ (.A(_07173_),
    .B(_06733_),
    .C(_07174_),
    .Y(_07178_));
 sky130_fd_sc_hd__nand2_2 _17646_ (.A(_07177_),
    .B(_07178_),
    .Y(_07179_));
 sky130_fd_sc_hd__nand3_1 _17647_ (.A(_07141_),
    .B(_07164_),
    .C(_07160_),
    .Y(_07180_));
 sky130_fd_sc_hd__nand2_1 _17648_ (.A(_07180_),
    .B(_07158_),
    .Y(_07181_));
 sky130_fd_sc_hd__nand3_1 _17649_ (.A(_07181_),
    .B(_07151_),
    .C(_07147_),
    .Y(_07182_));
 sky130_fd_sc_hd__nand2_1 _17650_ (.A(_07147_),
    .B(_07151_),
    .Y(_07183_));
 sky130_fd_sc_hd__nand3_1 _17651_ (.A(_07180_),
    .B(_07183_),
    .C(_07158_),
    .Y(_07184_));
 sky130_fd_sc_hd__a21o_1 _17652_ (.A1(_07182_),
    .A2(_07184_),
    .B1(_06972_),
    .X(_07185_));
 sky130_fd_sc_hd__nand2_1 _17653_ (.A(net157),
    .B(_07145_),
    .Y(_07186_));
 sky130_fd_sc_hd__nand2_1 _17654_ (.A(_07185_),
    .B(_07186_),
    .Y(_07188_));
 sky130_fd_sc_hd__nand2_1 _17655_ (.A(_07188_),
    .B(_06721_),
    .Y(_07189_));
 sky130_fd_sc_hd__nand3_2 _17656_ (.A(_07185_),
    .B(_06723_),
    .C(_07186_),
    .Y(_07190_));
 sky130_fd_sc_hd__nand2_2 _17657_ (.A(_07189_),
    .B(_07190_),
    .Y(_07191_));
 sky130_fd_sc_hd__nor2_2 _17658_ (.A(_07179_),
    .B(_07191_),
    .Y(_07192_));
 sky130_fd_sc_hd__a21o_1 _17659_ (.A1(_07141_),
    .A2(_07164_),
    .B1(_07160_),
    .X(_07193_));
 sky130_fd_sc_hd__nand3_1 _17660_ (.A(_07171_),
    .B(_07180_),
    .C(_07193_),
    .Y(_07194_));
 sky130_fd_sc_hd__a21o_1 _17661_ (.A1(_06969_),
    .A2(_06970_),
    .B1(_07153_),
    .X(_07195_));
 sky130_fd_sc_hd__nand2_1 _17662_ (.A(_07194_),
    .B(_07195_),
    .Y(_07196_));
 sky130_fd_sc_hd__nand2_1 _17663_ (.A(_07196_),
    .B(_06695_),
    .Y(_07197_));
 sky130_fd_sc_hd__nand3_1 _17664_ (.A(_07194_),
    .B(_06697_),
    .C(_07195_),
    .Y(_07199_));
 sky130_fd_sc_hd__nand2_2 _17665_ (.A(_07197_),
    .B(_07199_),
    .Y(_07200_));
 sky130_fd_sc_hd__nand2_1 _17666_ (.A(_07164_),
    .B(_07138_),
    .Y(_07201_));
 sky130_fd_sc_hd__nand2_1 _17667_ (.A(_07062_),
    .B(_07023_),
    .Y(_07202_));
 sky130_fd_sc_hd__xor2_1 _17668_ (.A(_07201_),
    .B(_07202_),
    .X(_07203_));
 sky130_fd_sc_hd__nand2_1 _17669_ (.A(_07171_),
    .B(_07203_),
    .Y(_07204_));
 sky130_fd_sc_hd__nand2_1 _17670_ (.A(_06972_),
    .B(_07163_),
    .Y(_07205_));
 sky130_fd_sc_hd__nand2_1 _17671_ (.A(_07204_),
    .B(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__or2_4 _17672_ (.A(_05915_),
    .B(_07206_),
    .X(_07207_));
 sky130_fd_sc_hd__nand2_1 _17673_ (.A(_07206_),
    .B(_05915_),
    .Y(_07208_));
 sky130_fd_sc_hd__nand2_2 _17674_ (.A(_07207_),
    .B(_07208_),
    .Y(_07210_));
 sky130_fd_sc_hd__nor2_2 _17675_ (.A(_07200_),
    .B(_07210_),
    .Y(_07211_));
 sky130_fd_sc_hd__nand2_1 _17676_ (.A(_07192_),
    .B(_07211_),
    .Y(_07212_));
 sky130_fd_sc_hd__inv_2 _17677_ (.A(_07212_),
    .Y(_07213_));
 sky130_fd_sc_hd__nand2_1 _17678_ (.A(_07117_),
    .B(_07213_),
    .Y(_07214_));
 sky130_fd_sc_hd__o21ai_2 _17679_ (.A1(_07207_),
    .A2(_07200_),
    .B1(_07197_),
    .Y(_07215_));
 sky130_fd_sc_hd__o21ai_1 _17680_ (.A1(_07190_),
    .A2(_07179_),
    .B1(_07177_),
    .Y(_07216_));
 sky130_fd_sc_hd__a21oi_1 _17681_ (.A1(_07215_),
    .A2(_07192_),
    .B1(_07216_),
    .Y(_07217_));
 sky130_fd_sc_hd__nand2_2 _17682_ (.A(_07217_),
    .B(_07214_),
    .Y(_07218_));
 sky130_fd_sc_hd__inv_2 _17683_ (.A(_07166_),
    .Y(_07219_));
 sky130_fd_sc_hd__nand2_1 _17684_ (.A(_07124_),
    .B(_06724_),
    .Y(_07221_));
 sky130_fd_sc_hd__clkinvlp_2 _17685_ (.A(_06735_),
    .Y(_07222_));
 sky130_fd_sc_hd__nand2_1 _17686_ (.A(_07221_),
    .B(_07222_),
    .Y(_07223_));
 sky130_fd_sc_hd__nand3_1 _17687_ (.A(_07124_),
    .B(_06735_),
    .C(_06724_),
    .Y(_07224_));
 sky130_fd_sc_hd__nand2_1 _17688_ (.A(_07223_),
    .B(_07224_),
    .Y(_07225_));
 sky130_fd_sc_hd__buf_6 _17689_ (.A(_05288_),
    .X(_07226_));
 sky130_fd_sc_hd__nand2_1 _17690_ (.A(_07225_),
    .B(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__buf_6 _17691_ (.A(net35),
    .X(_07228_));
 sky130_fd_sc_hd__nand3_1 _17692_ (.A(_07223_),
    .B(_07228_),
    .C(_07224_),
    .Y(_07229_));
 sky130_fd_sc_hd__nand3_1 _17693_ (.A(_07134_),
    .B(_07227_),
    .C(_07229_),
    .Y(_07230_));
 sky130_fd_sc_hd__inv_2 _17694_ (.A(_07230_),
    .Y(_07232_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(_07219_),
    .B(_07232_),
    .Y(_07233_));
 sky130_fd_sc_hd__nor2_1 _17696_ (.A(_07168_),
    .B(_07230_),
    .Y(_07234_));
 sky130_fd_sc_hd__nand2_1 _17697_ (.A(_07227_),
    .B(_07229_),
    .Y(_07235_));
 sky130_fd_sc_hd__o21ai_1 _17698_ (.A1(_07129_),
    .A2(_07235_),
    .B1(_07229_),
    .Y(_07236_));
 sky130_fd_sc_hd__nor2_1 _17699_ (.A(_07234_),
    .B(_07236_),
    .Y(_07237_));
 sky130_fd_sc_hd__nand2_2 _17700_ (.A(_07233_),
    .B(_07237_),
    .Y(_07238_));
 sky130_fd_sc_hd__inv_2 _17701_ (.A(_06750_),
    .Y(_07239_));
 sky130_fd_sc_hd__inv_2 _17702_ (.A(_06749_),
    .Y(_07240_));
 sky130_fd_sc_hd__nand2_1 _17703_ (.A(_06745_),
    .B(_07240_),
    .Y(_07241_));
 sky130_fd_sc_hd__nand2_1 _17704_ (.A(_07241_),
    .B(_06586_),
    .Y(_07243_));
 sky130_fd_sc_hd__or2_1 _17705_ (.A(_07239_),
    .B(_07243_),
    .X(_07244_));
 sky130_fd_sc_hd__nand2_1 _17706_ (.A(_07243_),
    .B(_07239_),
    .Y(_07245_));
 sky130_fd_sc_hd__nand2_1 _17707_ (.A(_07244_),
    .B(_07245_),
    .Y(_07246_));
 sky130_fd_sc_hd__buf_6 _17708_ (.A(_06045_),
    .X(_07247_));
 sky130_fd_sc_hd__nand2_1 _17709_ (.A(_07246_),
    .B(_07247_),
    .Y(_07248_));
 sky130_fd_sc_hd__buf_6 _17710_ (.A(net37),
    .X(_07249_));
 sky130_fd_sc_hd__nand3_1 _17711_ (.A(_07244_),
    .B(_07249_),
    .C(_07245_),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_1 _17712_ (.A(_07248_),
    .B(_07250_),
    .Y(_07251_));
 sky130_fd_sc_hd__inv_2 _17713_ (.A(_07251_),
    .Y(_07252_));
 sky130_fd_sc_hd__or2_1 _17714_ (.A(_07240_),
    .B(_06745_),
    .X(_07254_));
 sky130_fd_sc_hd__nand2_1 _17715_ (.A(_07254_),
    .B(_07241_),
    .Y(_07255_));
 sky130_fd_sc_hd__inv_2 _17716_ (.A(_07255_),
    .Y(_07256_));
 sky130_fd_sc_hd__nand2_1 _17717_ (.A(_07256_),
    .B(_06521_),
    .Y(_07257_));
 sky130_fd_sc_hd__nand2_1 _17718_ (.A(_07255_),
    .B(_06012_),
    .Y(_07258_));
 sky130_fd_sc_hd__nand2_2 _17719_ (.A(_07257_),
    .B(_07258_),
    .Y(_07259_));
 sky130_fd_sc_hd__inv_4 _17720_ (.A(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__nand2_1 _17721_ (.A(_07252_),
    .B(_07260_),
    .Y(_07261_));
 sky130_fd_sc_hd__inv_2 _17722_ (.A(_07261_),
    .Y(_07262_));
 sky130_fd_sc_hd__nand2_1 _17723_ (.A(_07238_),
    .B(_07262_),
    .Y(_07263_));
 sky130_fd_sc_hd__inv_2 _17724_ (.A(_07257_),
    .Y(_07265_));
 sky130_fd_sc_hd__a21boi_2 _17725_ (.A1(_07248_),
    .A2(_07265_),
    .B1_N(_07250_),
    .Y(_07266_));
 sky130_fd_sc_hd__nand2_1 _17726_ (.A(_07263_),
    .B(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__nand2_1 _17727_ (.A(_06745_),
    .B(_06751_),
    .Y(_07268_));
 sky130_fd_sc_hd__inv_2 _17728_ (.A(_06595_),
    .Y(_07269_));
 sky130_fd_sc_hd__nand2_1 _17729_ (.A(_07268_),
    .B(_07269_),
    .Y(_07270_));
 sky130_fd_sc_hd__inv_2 _17730_ (.A(_06573_),
    .Y(_07271_));
 sky130_fd_sc_hd__nand2_1 _17731_ (.A(_07270_),
    .B(_07271_),
    .Y(_07272_));
 sky130_fd_sc_hd__nand3_1 _17732_ (.A(_07268_),
    .B(_07269_),
    .C(_06573_),
    .Y(_07273_));
 sky130_fd_sc_hd__nand2_1 _17733_ (.A(_07272_),
    .B(_07273_),
    .Y(_07274_));
 sky130_fd_sc_hd__buf_6 _17734_ (.A(_06155_),
    .X(_07276_));
 sky130_fd_sc_hd__nand2_1 _17735_ (.A(_07274_),
    .B(_07276_),
    .Y(_07277_));
 sky130_fd_sc_hd__buf_6 _17736_ (.A(net38),
    .X(_07278_));
 sky130_fd_sc_hd__nand3_1 _17737_ (.A(_07272_),
    .B(_07273_),
    .C(_07278_),
    .Y(_07279_));
 sky130_fd_sc_hd__nand2_1 _17738_ (.A(_07277_),
    .B(_07279_),
    .Y(_07280_));
 sky130_fd_sc_hd__inv_2 _17739_ (.A(_07280_),
    .Y(_07281_));
 sky130_fd_sc_hd__nand2_1 _17740_ (.A(_07267_),
    .B(_07281_),
    .Y(_07282_));
 sky130_fd_sc_hd__nand3_1 _17741_ (.A(_07263_),
    .B(_07280_),
    .C(_07266_),
    .Y(_07283_));
 sky130_fd_sc_hd__nand3_1 _17742_ (.A(_07282_),
    .B(_07171_),
    .C(_07283_),
    .Y(_07284_));
 sky130_fd_sc_hd__or2_1 _17743_ (.A(_07274_),
    .B(_07171_),
    .X(_07285_));
 sky130_fd_sc_hd__nand2_1 _17744_ (.A(_07284_),
    .B(_07285_),
    .Y(_07287_));
 sky130_fd_sc_hd__nand2_1 _17745_ (.A(_07287_),
    .B(_06554_),
    .Y(_07288_));
 sky130_fd_sc_hd__nand3_1 _17746_ (.A(_07284_),
    .B(_06556_),
    .C(_07285_),
    .Y(_07289_));
 sky130_fd_sc_hd__nand2_2 _17747_ (.A(_07288_),
    .B(_07289_),
    .Y(_07290_));
 sky130_fd_sc_hd__nand2_1 _17748_ (.A(_07238_),
    .B(_07260_),
    .Y(_07291_));
 sky130_fd_sc_hd__nand2_1 _17749_ (.A(_07291_),
    .B(_07257_),
    .Y(_07292_));
 sky130_fd_sc_hd__nand2_1 _17750_ (.A(_07292_),
    .B(_07252_),
    .Y(_07293_));
 sky130_fd_sc_hd__nand3_1 _17751_ (.A(_07291_),
    .B(_07251_),
    .C(_07257_),
    .Y(_07294_));
 sky130_fd_sc_hd__nand2_1 _17752_ (.A(_07293_),
    .B(_07294_),
    .Y(_07295_));
 sky130_fd_sc_hd__nand2_1 _17753_ (.A(_07295_),
    .B(_07171_),
    .Y(_07296_));
 sky130_fd_sc_hd__nand2_1 _17754_ (.A(\div1i.quot[17] ),
    .B(_07246_),
    .Y(_07298_));
 sky130_fd_sc_hd__nand2_1 _17755_ (.A(_07296_),
    .B(_07298_),
    .Y(_07299_));
 sky130_fd_sc_hd__nand2_1 _17756_ (.A(_07299_),
    .B(_06568_),
    .Y(_07300_));
 sky130_fd_sc_hd__nand3_2 _17757_ (.A(_07296_),
    .B(_06570_),
    .C(_07298_),
    .Y(_07301_));
 sky130_fd_sc_hd__nand2_2 _17758_ (.A(_07300_),
    .B(_07301_),
    .Y(_07302_));
 sky130_fd_sc_hd__nor2_2 _17759_ (.A(_07290_),
    .B(_07302_),
    .Y(_07303_));
 sky130_fd_sc_hd__or2_1 _17760_ (.A(_07260_),
    .B(_07238_),
    .X(_07304_));
 sky130_fd_sc_hd__nand3_1 _17761_ (.A(_07304_),
    .B(_07171_),
    .C(_07291_),
    .Y(_07305_));
 sky130_fd_sc_hd__nand2_1 _17762_ (.A(net157),
    .B(_07256_),
    .Y(_07306_));
 sky130_fd_sc_hd__nand2_1 _17763_ (.A(_07305_),
    .B(_07306_),
    .Y(_07307_));
 sky130_fd_sc_hd__nand2_1 _17764_ (.A(_07307_),
    .B(_06149_),
    .Y(_07309_));
 sky130_fd_sc_hd__nand3_1 _17765_ (.A(_07305_),
    .B(_06592_),
    .C(_07306_),
    .Y(_07310_));
 sky130_fd_sc_hd__nand2_1 _17766_ (.A(_07309_),
    .B(_07310_),
    .Y(_07311_));
 sky130_fd_sc_hd__nand2_1 _17767_ (.A(_07172_),
    .B(_07129_),
    .Y(_07312_));
 sky130_fd_sc_hd__xor2_1 _17768_ (.A(_07235_),
    .B(_07312_),
    .X(_07313_));
 sky130_fd_sc_hd__nand2_1 _17769_ (.A(_07313_),
    .B(_07171_),
    .Y(_07314_));
 sky130_fd_sc_hd__nand2_1 _17770_ (.A(\div1i.quot[17] ),
    .B(_07225_),
    .Y(_07315_));
 sky130_fd_sc_hd__nand2_1 _17771_ (.A(_07314_),
    .B(_07315_),
    .Y(_07316_));
 sky130_fd_sc_hd__nand2_1 _17772_ (.A(_07316_),
    .B(_06159_),
    .Y(_07317_));
 sky130_fd_sc_hd__buf_6 _17773_ (.A(_08296_),
    .X(_07318_));
 sky130_fd_sc_hd__nand3_2 _17774_ (.A(_07314_),
    .B(_07318_),
    .C(_07315_),
    .Y(_07320_));
 sky130_fd_sc_hd__nand2_2 _17775_ (.A(_07317_),
    .B(_07320_),
    .Y(_07321_));
 sky130_fd_sc_hd__nor2_2 _17776_ (.A(_07311_),
    .B(_07321_),
    .Y(_07322_));
 sky130_fd_sc_hd__nand2_1 _17777_ (.A(_07303_),
    .B(_07322_),
    .Y(_07323_));
 sky130_fd_sc_hd__inv_2 _17778_ (.A(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__nand2_2 _17779_ (.A(_07218_),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__o21ai_2 _17780_ (.A1(_07320_),
    .A2(_07311_),
    .B1(_07309_),
    .Y(_07326_));
 sky130_fd_sc_hd__o21ai_1 _17781_ (.A1(_07301_),
    .A2(_07290_),
    .B1(_07288_),
    .Y(_07327_));
 sky130_fd_sc_hd__a21oi_2 _17782_ (.A1(_07303_),
    .A2(_07326_),
    .B1(_07327_),
    .Y(_07328_));
 sky130_fd_sc_hd__nand2_4 _17783_ (.A(_07325_),
    .B(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__nand2_1 _17784_ (.A(_07272_),
    .B(_06571_),
    .Y(_07331_));
 sky130_fd_sc_hd__inv_2 _17785_ (.A(_06558_),
    .Y(_07332_));
 sky130_fd_sc_hd__nand2_1 _17786_ (.A(_07331_),
    .B(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__nand3_1 _17787_ (.A(_07272_),
    .B(_06558_),
    .C(_06571_),
    .Y(_07334_));
 sky130_fd_sc_hd__nand2_1 _17788_ (.A(_07333_),
    .B(_07334_),
    .Y(_07335_));
 sky130_fd_sc_hd__nand2_1 _17789_ (.A(_07335_),
    .B(_05375_),
    .Y(_07336_));
 sky130_fd_sc_hd__nand3_1 _17790_ (.A(_07333_),
    .B(_06772_),
    .C(_07334_),
    .Y(_07337_));
 sky130_fd_sc_hd__nand3_1 _17791_ (.A(_07336_),
    .B(_07337_),
    .C(_07281_),
    .Y(_07338_));
 sky130_fd_sc_hd__nor2_1 _17792_ (.A(_07338_),
    .B(_07261_),
    .Y(_07339_));
 sky130_fd_sc_hd__nand2_2 _17793_ (.A(_07238_),
    .B(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__nor2_1 _17794_ (.A(_07338_),
    .B(_07266_),
    .Y(_07342_));
 sky130_fd_sc_hd__nand2_1 _17795_ (.A(_07336_),
    .B(_07337_),
    .Y(_07343_));
 sky130_fd_sc_hd__o21ai_1 _17796_ (.A1(_07279_),
    .A2(_07343_),
    .B1(_07337_),
    .Y(_07344_));
 sky130_fd_sc_hd__nor2_1 _17797_ (.A(_07342_),
    .B(_07344_),
    .Y(_07345_));
 sky130_fd_sc_hd__nand2_2 _17798_ (.A(_07345_),
    .B(_07340_),
    .Y(_07346_));
 sky130_fd_sc_hd__clkinvlp_2 _17799_ (.A(_06789_),
    .Y(_07347_));
 sky130_fd_sc_hd__inv_2 _17800_ (.A(_06801_),
    .Y(_07348_));
 sky130_fd_sc_hd__nand2_1 _17801_ (.A(_06753_),
    .B(_07348_),
    .Y(_07349_));
 sky130_fd_sc_hd__nand2_1 _17802_ (.A(_07349_),
    .B(_06800_),
    .Y(_07350_));
 sky130_fd_sc_hd__or2_1 _17803_ (.A(_07347_),
    .B(_07350_),
    .X(_07351_));
 sky130_fd_sc_hd__nand2_1 _17804_ (.A(_07350_),
    .B(_07347_),
    .Y(_07353_));
 sky130_fd_sc_hd__nand2_1 _17805_ (.A(_07351_),
    .B(_07353_),
    .Y(_07354_));
 sky130_fd_sc_hd__nand2_1 _17806_ (.A(_07354_),
    .B(_06814_),
    .Y(_07355_));
 sky130_fd_sc_hd__nand3_1 _17807_ (.A(_07351_),
    .B(_06827_),
    .C(_07353_),
    .Y(_07356_));
 sky130_fd_sc_hd__nand2_1 _17808_ (.A(_07355_),
    .B(_07356_),
    .Y(_07357_));
 sky130_fd_sc_hd__or2_1 _17809_ (.A(_07348_),
    .B(_06753_),
    .X(_07358_));
 sky130_fd_sc_hd__nand2_1 _17810_ (.A(_07358_),
    .B(_07349_),
    .Y(_07359_));
 sky130_fd_sc_hd__inv_2 _17811_ (.A(_07359_),
    .Y(_07360_));
 sky130_fd_sc_hd__nand2_1 _17812_ (.A(_07360_),
    .B(_06207_),
    .Y(_07361_));
 sky130_fd_sc_hd__nand2_1 _17813_ (.A(_07359_),
    .B(_05408_),
    .Y(_07362_));
 sky130_fd_sc_hd__nand2_1 _17814_ (.A(_07361_),
    .B(_07362_),
    .Y(_07364_));
 sky130_fd_sc_hd__inv_2 _17815_ (.A(_07364_),
    .Y(_07365_));
 sky130_fd_sc_hd__nand2b_1 _17816_ (.A_N(_07357_),
    .B(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__inv_2 _17817_ (.A(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__nand2_1 _17818_ (.A(_07346_),
    .B(_07367_),
    .Y(_07368_));
 sky130_fd_sc_hd__inv_2 _17819_ (.A(_07361_),
    .Y(_07369_));
 sky130_fd_sc_hd__a21boi_2 _17820_ (.A1(_07355_),
    .A2(_07369_),
    .B1_N(_07356_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand2_1 _17821_ (.A(_07368_),
    .B(_07370_),
    .Y(_07371_));
 sky130_fd_sc_hd__inv_2 _17822_ (.A(_06853_),
    .Y(_07372_));
 sky130_fd_sc_hd__nand2_1 _17823_ (.A(_06808_),
    .B(_07372_),
    .Y(_07373_));
 sky130_fd_sc_hd__nand3_1 _17824_ (.A(_06804_),
    .B(_06807_),
    .C(_06853_),
    .Y(_07375_));
 sky130_fd_sc_hd__nand2_2 _17825_ (.A(_07373_),
    .B(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__inv_2 _17826_ (.A(_07376_),
    .Y(_07377_));
 sky130_fd_sc_hd__nand2_1 _17827_ (.A(_07377_),
    .B(_06819_),
    .Y(_07378_));
 sky130_fd_sc_hd__nand2_1 _17828_ (.A(_07376_),
    .B(_06737_),
    .Y(_07379_));
 sky130_fd_sc_hd__nand2_2 _17829_ (.A(_07378_),
    .B(_07379_),
    .Y(_07380_));
 sky130_fd_sc_hd__inv_2 _17830_ (.A(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__nand2_1 _17831_ (.A(_07371_),
    .B(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__buf_6 _17832_ (.A(_07171_),
    .X(_07383_));
 sky130_fd_sc_hd__nand3_1 _17833_ (.A(_07368_),
    .B(_07380_),
    .C(_07370_),
    .Y(_07384_));
 sky130_fd_sc_hd__nand3_2 _17834_ (.A(_07382_),
    .B(_07383_),
    .C(_07384_),
    .Y(_07386_));
 sky130_fd_sc_hd__nand2_1 _17835_ (.A(\div1i.quot[17] ),
    .B(_07377_),
    .Y(_07387_));
 sky130_fd_sc_hd__nand2_1 _17836_ (.A(_07386_),
    .B(_07387_),
    .Y(_07388_));
 sky130_fd_sc_hd__nand2_1 _17837_ (.A(_07388_),
    .B(_06856_),
    .Y(_07389_));
 sky130_fd_sc_hd__nand3_1 _17838_ (.A(_07386_),
    .B(_06809_),
    .C(_07387_),
    .Y(_07390_));
 sky130_fd_sc_hd__nand2_2 _17839_ (.A(_07389_),
    .B(_07390_),
    .Y(_07391_));
 sky130_fd_sc_hd__nand2_1 _17840_ (.A(_07346_),
    .B(_07365_),
    .Y(_07392_));
 sky130_fd_sc_hd__nand2_1 _17841_ (.A(_07392_),
    .B(_07361_),
    .Y(_07393_));
 sky130_fd_sc_hd__xor2_1 _17842_ (.A(_07357_),
    .B(_07393_),
    .X(_07394_));
 sky130_fd_sc_hd__nand2_1 _17843_ (.A(_07394_),
    .B(_07383_),
    .Y(_07395_));
 sky130_fd_sc_hd__nand2_1 _17844_ (.A(\div1i.quot[17] ),
    .B(_07354_),
    .Y(_07397_));
 sky130_fd_sc_hd__nand2_1 _17845_ (.A(_07395_),
    .B(_07397_),
    .Y(_07398_));
 sky130_fd_sc_hd__nand2_1 _17846_ (.A(_07398_),
    .B(_06844_),
    .Y(_07399_));
 sky130_fd_sc_hd__buf_8 _17847_ (.A(net120),
    .X(_07400_));
 sky130_fd_sc_hd__nand3_4 _17848_ (.A(_07395_),
    .B(_07400_),
    .C(_07397_),
    .Y(_07401_));
 sky130_fd_sc_hd__nand2_2 _17849_ (.A(_07399_),
    .B(_07401_),
    .Y(_07402_));
 sky130_fd_sc_hd__nor2_2 _17850_ (.A(_07391_),
    .B(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__nand3_1 _17851_ (.A(_07340_),
    .B(_07345_),
    .C(_07364_),
    .Y(_07404_));
 sky130_fd_sc_hd__nand3_1 _17852_ (.A(_07392_),
    .B(_07171_),
    .C(_07404_),
    .Y(_07405_));
 sky130_fd_sc_hd__nand2_1 _17853_ (.A(net157),
    .B(_07360_),
    .Y(_07406_));
 sky130_fd_sc_hd__nand2_1 _17854_ (.A(_07405_),
    .B(_07406_),
    .Y(_07408_));
 sky130_fd_sc_hd__or2_1 _17855_ (.A(_06805_),
    .B(_07408_),
    .X(_07409_));
 sky130_fd_sc_hd__nand2_1 _17856_ (.A(_07408_),
    .B(_06805_),
    .Y(_07410_));
 sky130_fd_sc_hd__nand2_2 _17857_ (.A(_07409_),
    .B(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__nand2_1 _17858_ (.A(_07282_),
    .B(_07279_),
    .Y(_07412_));
 sky130_fd_sc_hd__xor2_1 _17859_ (.A(_07343_),
    .B(_07412_),
    .X(_07413_));
 sky130_fd_sc_hd__nand2_1 _17860_ (.A(_07413_),
    .B(_07383_),
    .Y(_07414_));
 sky130_fd_sc_hd__nand2_1 _17861_ (.A(\div1i.quot[17] ),
    .B(_07335_),
    .Y(_07415_));
 sky130_fd_sc_hd__nand2_1 _17862_ (.A(_07414_),
    .B(_07415_),
    .Y(_07416_));
 sky130_fd_sc_hd__nand2_1 _17863_ (.A(_07416_),
    .B(_06797_),
    .Y(_07417_));
 sky130_fd_sc_hd__nand3_2 _17864_ (.A(_07414_),
    .B(_06799_),
    .C(_07415_),
    .Y(_07419_));
 sky130_fd_sc_hd__nand3b_2 _17865_ (.A_N(_07411_),
    .B(_07417_),
    .C(_07419_),
    .Y(_07420_));
 sky130_fd_sc_hd__inv_4 _17866_ (.A(_07420_),
    .Y(_07421_));
 sky130_fd_sc_hd__nand3_4 _17867_ (.A(_07329_),
    .B(_07403_),
    .C(_07421_),
    .Y(_07422_));
 sky130_fd_sc_hd__o21ai_2 _17868_ (.A1(_07411_),
    .A2(_07419_),
    .B1(_07410_),
    .Y(_07423_));
 sky130_fd_sc_hd__o21ai_1 _17869_ (.A1(_07391_),
    .A2(_07401_),
    .B1(_07389_),
    .Y(_07424_));
 sky130_fd_sc_hd__a21oi_2 _17870_ (.A1(_07403_),
    .A2(_07423_),
    .B1(_07424_),
    .Y(_07425_));
 sky130_fd_sc_hd__nand2_4 _17871_ (.A(_07422_),
    .B(_07425_),
    .Y(_07426_));
 sky130_fd_sc_hd__nand2_1 _17872_ (.A(_07373_),
    .B(_06851_),
    .Y(_07427_));
 sky130_fd_sc_hd__inv_2 _17873_ (.A(_06843_),
    .Y(_07428_));
 sky130_fd_sc_hd__nand2_1 _17874_ (.A(_07427_),
    .B(_07428_),
    .Y(_07430_));
 sky130_fd_sc_hd__nand3_1 _17875_ (.A(_07373_),
    .B(_06843_),
    .C(_06851_),
    .Y(_07431_));
 sky130_fd_sc_hd__nand2_1 _17876_ (.A(_07430_),
    .B(_07431_),
    .Y(_07432_));
 sky130_fd_sc_hd__nand2_2 _17877_ (.A(_07432_),
    .B(_06704_),
    .Y(_07433_));
 sky130_fd_sc_hd__nand3_1 _17878_ (.A(_07430_),
    .B(_06874_),
    .C(_07431_),
    .Y(_07434_));
 sky130_fd_sc_hd__nand3_2 _17879_ (.A(_07381_),
    .B(_07433_),
    .C(_07434_),
    .Y(_07435_));
 sky130_fd_sc_hd__inv_2 _17880_ (.A(_07435_),
    .Y(_07436_));
 sky130_fd_sc_hd__nand3_2 _17881_ (.A(_07346_),
    .B(_07367_),
    .C(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__inv_2 _17882_ (.A(_07433_),
    .Y(_07438_));
 sky130_fd_sc_hd__o21ai_1 _17883_ (.A1(_07378_),
    .A2(_07438_),
    .B1(_07434_),
    .Y(_07439_));
 sky130_fd_sc_hd__nor2_1 _17884_ (.A(_07370_),
    .B(_07435_),
    .Y(_07441_));
 sky130_fd_sc_hd__nor2_1 _17885_ (.A(_07439_),
    .B(_07441_),
    .Y(_07442_));
 sky130_fd_sc_hd__nand2_2 _17886_ (.A(_07437_),
    .B(_07442_),
    .Y(_07443_));
 sky130_fd_sc_hd__inv_2 _17887_ (.A(net240),
    .Y(_07444_));
 sky130_fd_sc_hd__nand2_1 _17888_ (.A(_06904_),
    .B(_06900_),
    .Y(_07445_));
 sky130_fd_sc_hd__nand2_1 _17889_ (.A(_07444_),
    .B(_07445_),
    .Y(_07446_));
 sky130_fd_sc_hd__inv_2 _17890_ (.A(_07445_),
    .Y(_07447_));
 sky130_fd_sc_hd__nand2_2 _17891_ (.A(net240),
    .B(_07447_),
    .Y(_07448_));
 sky130_fd_sc_hd__nand2_1 _17892_ (.A(_07446_),
    .B(_07448_),
    .Y(_07449_));
 sky130_fd_sc_hd__buf_6 _17893_ (.A(_10426_),
    .X(_07450_));
 sky130_fd_sc_hd__nand2_1 _17894_ (.A(_07449_),
    .B(_07450_),
    .Y(_07452_));
 sky130_fd_sc_hd__nand3_2 _17895_ (.A(_07446_),
    .B(_06649_),
    .C(_07448_),
    .Y(_07453_));
 sky130_fd_sc_hd__nand2_1 _17896_ (.A(_07452_),
    .B(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__inv_2 _17897_ (.A(_07454_),
    .Y(_07455_));
 sky130_fd_sc_hd__nand2_2 _17898_ (.A(_07443_),
    .B(_07455_),
    .Y(_07456_));
 sky130_fd_sc_hd__nand2_1 _17899_ (.A(_07456_),
    .B(_07453_),
    .Y(_07457_));
 sky130_fd_sc_hd__nand2_1 _17900_ (.A(_07448_),
    .B(_06900_),
    .Y(_07458_));
 sky130_fd_sc_hd__xor2_2 _17901_ (.A(_06892_),
    .B(_07458_),
    .X(_07459_));
 sky130_fd_sc_hd__inv_2 _17902_ (.A(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__buf_6 _17903_ (.A(net46),
    .X(_07461_));
 sky130_fd_sc_hd__nand2_1 _17904_ (.A(_07460_),
    .B(_07461_),
    .Y(_07463_));
 sky130_fd_sc_hd__nand2_2 _17905_ (.A(_07459_),
    .B(_06550_),
    .Y(_07464_));
 sky130_fd_sc_hd__nand2_1 _17906_ (.A(_07463_),
    .B(_07464_),
    .Y(_07465_));
 sky130_fd_sc_hd__inv_2 _17907_ (.A(_07465_),
    .Y(_07466_));
 sky130_fd_sc_hd__nand2_1 _17908_ (.A(_07457_),
    .B(_07466_),
    .Y(_07467_));
 sky130_fd_sc_hd__nand3_1 _17909_ (.A(_07456_),
    .B(_07465_),
    .C(_07453_),
    .Y(_07468_));
 sky130_fd_sc_hd__nand2_1 _17910_ (.A(_07467_),
    .B(_07468_),
    .Y(_07469_));
 sky130_fd_sc_hd__nand2_1 _17911_ (.A(_07469_),
    .B(_07383_),
    .Y(_07470_));
 sky130_fd_sc_hd__nand2_1 _17912_ (.A(_07459_),
    .B(\div1i.quot[17] ),
    .Y(_07471_));
 sky130_fd_sc_hd__nand2_1 _17913_ (.A(_07470_),
    .B(_07471_),
    .Y(_07472_));
 sky130_fd_sc_hd__buf_6 _17914_ (.A(_10701_),
    .X(_07474_));
 sky130_fd_sc_hd__nand2_1 _17915_ (.A(_07472_),
    .B(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__nand3_1 _17916_ (.A(_07470_),
    .B(_06366_),
    .C(_07471_),
    .Y(_07476_));
 sky130_fd_sc_hd__nand2_1 _17917_ (.A(_07475_),
    .B(_07476_),
    .Y(_07477_));
 sky130_fd_sc_hd__inv_2 _17918_ (.A(_07477_),
    .Y(_07478_));
 sky130_fd_sc_hd__nand3_1 _17919_ (.A(_07463_),
    .B(_07464_),
    .C(_07455_),
    .Y(_07479_));
 sky130_fd_sc_hd__inv_2 _17920_ (.A(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__nand2_1 _17921_ (.A(_07480_),
    .B(_07443_),
    .Y(_07481_));
 sky130_fd_sc_hd__inv_2 _17922_ (.A(_07464_),
    .Y(_07482_));
 sky130_fd_sc_hd__o21a_1 _17923_ (.A1(_07453_),
    .A2(_07482_),
    .B1(_07463_),
    .X(_07483_));
 sky130_fd_sc_hd__nand2_1 _17924_ (.A(_07481_),
    .B(_07483_),
    .Y(_07485_));
 sky130_fd_sc_hd__o21bai_1 _17925_ (.A1(_06905_),
    .A2(_07444_),
    .B1_N(_06958_),
    .Y(_07486_));
 sky130_fd_sc_hd__or2_1 _17926_ (.A(_06926_),
    .B(_07486_),
    .X(_07487_));
 sky130_fd_sc_hd__nand2_1 _17927_ (.A(_07486_),
    .B(_06926_),
    .Y(_07488_));
 sky130_fd_sc_hd__nand2_1 _17928_ (.A(_07487_),
    .B(_07488_),
    .Y(_07489_));
 sky130_fd_sc_hd__inv_2 _17929_ (.A(_07489_),
    .Y(_07490_));
 sky130_fd_sc_hd__nand2_1 _17930_ (.A(_07490_),
    .B(_06936_),
    .Y(_07491_));
 sky130_fd_sc_hd__nand2_1 _17931_ (.A(_07489_),
    .B(_06594_),
    .Y(_07492_));
 sky130_fd_sc_hd__nand2_1 _17932_ (.A(_07491_),
    .B(_07492_),
    .Y(_07493_));
 sky130_fd_sc_hd__inv_2 _17933_ (.A(_07493_),
    .Y(_07494_));
 sky130_fd_sc_hd__nand2_1 _17934_ (.A(_07485_),
    .B(_07494_),
    .Y(_07496_));
 sky130_fd_sc_hd__nand3_1 _17935_ (.A(_07481_),
    .B(_07483_),
    .C(_07493_),
    .Y(_07497_));
 sky130_fd_sc_hd__nand3_2 _17936_ (.A(_07496_),
    .B(_07497_),
    .C(_07383_),
    .Y(_07498_));
 sky130_fd_sc_hd__nand2_1 _17937_ (.A(_07490_),
    .B(\div1i.quot[17] ),
    .Y(_07499_));
 sky130_fd_sc_hd__nand2_1 _17938_ (.A(_07498_),
    .B(_07499_),
    .Y(_07500_));
 sky130_fd_sc_hd__nand2_1 _17939_ (.A(_07500_),
    .B(_06947_),
    .Y(_07501_));
 sky130_fd_sc_hd__nand3_2 _17940_ (.A(_07498_),
    .B(_06949_),
    .C(_07499_),
    .Y(_07502_));
 sky130_fd_sc_hd__nand2_2 _17941_ (.A(_07502_),
    .B(_07501_),
    .Y(_07503_));
 sky130_fd_sc_hd__inv_2 _17942_ (.A(_07503_),
    .Y(_07504_));
 sky130_fd_sc_hd__nand2_1 _17943_ (.A(_07478_),
    .B(_07504_),
    .Y(_07505_));
 sky130_fd_sc_hd__nand3_1 _17944_ (.A(_07437_),
    .B(_07442_),
    .C(_07454_),
    .Y(_07507_));
 sky130_fd_sc_hd__nand3_1 _17945_ (.A(_07456_),
    .B(_07507_),
    .C(_07383_),
    .Y(_07508_));
 sky130_fd_sc_hd__or2_1 _17946_ (.A(_07449_),
    .B(_07383_),
    .X(_07509_));
 sky130_fd_sc_hd__nand2_1 _17947_ (.A(_07508_),
    .B(_07509_),
    .Y(_07510_));
 sky130_fd_sc_hd__or2_1 _17948_ (.A(_06348_),
    .B(_07510_),
    .X(_07511_));
 sky130_fd_sc_hd__nand2_1 _17949_ (.A(_07510_),
    .B(_06348_),
    .Y(_07512_));
 sky130_fd_sc_hd__nand2_2 _17950_ (.A(_07511_),
    .B(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__nand2_1 _17951_ (.A(_07433_),
    .B(_07434_),
    .Y(_07514_));
 sky130_fd_sc_hd__nand2_1 _17952_ (.A(_07382_),
    .B(_07378_),
    .Y(_07515_));
 sky130_fd_sc_hd__xor2_1 _17953_ (.A(_07514_),
    .B(_07515_),
    .X(_07516_));
 sky130_fd_sc_hd__nand2_1 _17954_ (.A(_07516_),
    .B(_07383_),
    .Y(_07518_));
 sky130_fd_sc_hd__nand2_1 _17955_ (.A(\div1i.quot[17] ),
    .B(_07432_),
    .Y(_07519_));
 sky130_fd_sc_hd__nand3_2 _17956_ (.A(_07518_),
    .B(_06898_),
    .C(_07519_),
    .Y(_07520_));
 sky130_fd_sc_hd__nand2_1 _17957_ (.A(_07518_),
    .B(_07519_),
    .Y(_07521_));
 sky130_fd_sc_hd__nand2_1 _17958_ (.A(_07521_),
    .B(_06903_),
    .Y(_07522_));
 sky130_fd_sc_hd__nand3b_1 _17959_ (.A_N(_07513_),
    .B(_07520_),
    .C(_07522_),
    .Y(_07523_));
 sky130_fd_sc_hd__nor2_2 _17960_ (.A(_07505_),
    .B(_07523_),
    .Y(_07524_));
 sky130_fd_sc_hd__nand2_4 _17961_ (.A(_07426_),
    .B(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__o21ai_2 _17962_ (.A1(_07513_),
    .A2(_07520_),
    .B1(_07512_),
    .Y(_07526_));
 sky130_fd_sc_hd__nor2_1 _17963_ (.A(_07503_),
    .B(_07477_),
    .Y(_07527_));
 sky130_fd_sc_hd__inv_2 _17964_ (.A(_07502_),
    .Y(_07529_));
 sky130_fd_sc_hd__o21ai_1 _17965_ (.A1(_07476_),
    .A2(_07529_),
    .B1(_07501_),
    .Y(_07530_));
 sky130_fd_sc_hd__a21oi_2 _17966_ (.A1(_07526_),
    .A2(_07527_),
    .B1(_07530_),
    .Y(_07531_));
 sky130_fd_sc_hd__nand2_2 _17967_ (.A(_07531_),
    .B(_07525_),
    .Y(_07532_));
 sky130_fd_sc_hd__nand2_2 _17968_ (.A(_07488_),
    .B(_06923_),
    .Y(_07533_));
 sky130_fd_sc_hd__xor2_4 _17969_ (.A(net140),
    .B(_07533_),
    .X(_07534_));
 sky130_fd_sc_hd__nand3_2 _17970_ (.A(_07496_),
    .B(_07383_),
    .C(_07491_),
    .Y(_07535_));
 sky130_fd_sc_hd__xor2_4 _17971_ (.A(_07534_),
    .B(_07535_),
    .X(_07536_));
 sky130_fd_sc_hd__clkinvlp_2 _17972_ (.A(_07536_),
    .Y(_07537_));
 sky130_fd_sc_hd__nand2_4 _17973_ (.A(_07532_),
    .B(_07537_),
    .Y(_07538_));
 sky130_fd_sc_hd__nand3_4 _17974_ (.A(_07525_),
    .B(_07531_),
    .C(_07536_),
    .Y(_07540_));
 sky130_fd_sc_hd__nand2_8 _17975_ (.A(_07540_),
    .B(_07538_),
    .Y(_07541_));
 sky130_fd_sc_hd__buf_8 _17976_ (.A(_07541_),
    .X(_07542_));
 sky130_fd_sc_hd__buf_6 _17977_ (.A(_07542_),
    .X(\div1i.quot[16] ));
 sky130_fd_sc_hd__nand2_1 _17978_ (.A(_07117_),
    .B(_07211_),
    .Y(_07543_));
 sky130_fd_sc_hd__inv_2 _17979_ (.A(_07215_),
    .Y(_07544_));
 sky130_fd_sc_hd__nand2_1 _17980_ (.A(_07543_),
    .B(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__inv_2 _17981_ (.A(_07191_),
    .Y(_07546_));
 sky130_fd_sc_hd__nand2_2 _17982_ (.A(_07545_),
    .B(_07546_),
    .Y(_07547_));
 sky130_fd_sc_hd__nand2_1 _17983_ (.A(_07547_),
    .B(_07190_),
    .Y(_07548_));
 sky130_fd_sc_hd__inv_2 _17984_ (.A(_07179_),
    .Y(_07550_));
 sky130_fd_sc_hd__nand2_1 _17985_ (.A(_07548_),
    .B(_07550_),
    .Y(_07551_));
 sky130_fd_sc_hd__nand3_2 _17986_ (.A(_07547_),
    .B(_07190_),
    .C(_07179_),
    .Y(_07552_));
 sky130_fd_sc_hd__nand2_1 _17987_ (.A(_07551_),
    .B(_07552_),
    .Y(_07553_));
 sky130_fd_sc_hd__nand2_1 _17988_ (.A(_07553_),
    .B(_07226_),
    .Y(_07554_));
 sky130_fd_sc_hd__nand3_1 _17989_ (.A(_07543_),
    .B(_07191_),
    .C(_07544_),
    .Y(_07555_));
 sky130_fd_sc_hd__nand3_2 _17990_ (.A(_07547_),
    .B(_07128_),
    .C(_07555_),
    .Y(_07556_));
 sky130_fd_sc_hd__inv_2 _17991_ (.A(_07556_),
    .Y(_07557_));
 sky130_fd_sc_hd__nand3_2 _17992_ (.A(_07551_),
    .B(_07228_),
    .C(_07552_),
    .Y(_07558_));
 sky130_fd_sc_hd__nand3_1 _17993_ (.A(_07554_),
    .B(_07557_),
    .C(_07558_),
    .Y(_07559_));
 sky130_fd_sc_hd__nand2_1 _17994_ (.A(_07559_),
    .B(_07558_),
    .Y(_07561_));
 sky130_fd_sc_hd__inv_2 _17995_ (.A(_07210_),
    .Y(_07562_));
 sky130_fd_sc_hd__nand2_1 _17996_ (.A(_07117_),
    .B(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__nand2_1 _17997_ (.A(_07563_),
    .B(_07207_),
    .Y(_07564_));
 sky130_fd_sc_hd__inv_2 _17998_ (.A(_07200_),
    .Y(_07565_));
 sky130_fd_sc_hd__nand2_1 _17999_ (.A(_07564_),
    .B(_07565_),
    .Y(_07566_));
 sky130_fd_sc_hd__nand3_1 _18000_ (.A(_07563_),
    .B(_07200_),
    .C(_07207_),
    .Y(_07567_));
 sky130_fd_sc_hd__nand2_1 _18001_ (.A(_07566_),
    .B(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__nand2_1 _18002_ (.A(_07568_),
    .B(_07146_),
    .Y(_07569_));
 sky130_fd_sc_hd__or2_1 _18003_ (.A(_07562_),
    .B(_07117_),
    .X(_07570_));
 sky130_fd_sc_hd__nand2_1 _18004_ (.A(_07570_),
    .B(_07563_),
    .Y(_07572_));
 sky130_fd_sc_hd__inv_2 _18005_ (.A(_07572_),
    .Y(_07573_));
 sky130_fd_sc_hd__nand2_1 _18006_ (.A(_07573_),
    .B(_07157_),
    .Y(_07574_));
 sky130_fd_sc_hd__inv_2 _18007_ (.A(_07574_),
    .Y(_07575_));
 sky130_fd_sc_hd__inv_2 _18008_ (.A(_07568_),
    .Y(_07576_));
 sky130_fd_sc_hd__nand2_1 _18009_ (.A(_07576_),
    .B(_07149_),
    .Y(_07577_));
 sky130_fd_sc_hd__inv_2 _18010_ (.A(_07577_),
    .Y(_07578_));
 sky130_fd_sc_hd__a21oi_1 _18011_ (.A1(_07569_),
    .A2(_07575_),
    .B1(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__nand2_1 _18012_ (.A(_07547_),
    .B(_07555_),
    .Y(_07580_));
 sky130_fd_sc_hd__nand2_1 _18013_ (.A(_07580_),
    .B(_07130_),
    .Y(_07581_));
 sky130_fd_sc_hd__nand2_1 _18014_ (.A(_07581_),
    .B(_07556_),
    .Y(_07583_));
 sky130_fd_sc_hd__inv_2 _18015_ (.A(_07583_),
    .Y(_07584_));
 sky130_fd_sc_hd__nand3_1 _18016_ (.A(_07554_),
    .B(_07584_),
    .C(_07558_),
    .Y(_07585_));
 sky130_fd_sc_hd__nor2_1 _18017_ (.A(_07579_),
    .B(_07585_),
    .Y(_07586_));
 sky130_fd_sc_hd__nor2_1 _18018_ (.A(_07561_),
    .B(_07586_),
    .Y(_07587_));
 sky130_fd_sc_hd__inv_2 _18019_ (.A(_07585_),
    .Y(_07588_));
 sky130_fd_sc_hd__nand2_1 _18020_ (.A(_06999_),
    .B(_07003_),
    .Y(_07589_));
 sky130_fd_sc_hd__nand2_1 _18021_ (.A(_07589_),
    .B(_07005_),
    .Y(_07590_));
 sky130_fd_sc_hd__nand2_1 _18022_ (.A(_07590_),
    .B(net136),
    .Y(_07591_));
 sky130_fd_sc_hd__nand2_1 _18023_ (.A(_07591_),
    .B(_06982_),
    .Y(_07592_));
 sky130_fd_sc_hd__o21ai_2 _18024_ (.A1(_06979_),
    .A2(\div1i.quot[17] ),
    .B1(_06980_),
    .Y(_07594_));
 sky130_fd_sc_hd__nand3_1 _18025_ (.A(_07590_),
    .B(_06984_),
    .C(net136),
    .Y(_07595_));
 sky130_fd_sc_hd__inv_2 _18026_ (.A(_07595_),
    .Y(_07596_));
 sky130_fd_sc_hd__a21o_1 _18027_ (.A1(_07592_),
    .A2(_07594_),
    .B1(_07596_),
    .X(_07597_));
 sky130_fd_sc_hd__nand2_1 _18028_ (.A(_07008_),
    .B(_06991_),
    .Y(_07598_));
 sky130_fd_sc_hd__nand2_1 _18029_ (.A(net136),
    .B(_06999_),
    .Y(_07599_));
 sky130_fd_sc_hd__xor2_2 _18030_ (.A(_07598_),
    .B(_07599_),
    .X(_07600_));
 sky130_fd_sc_hd__nand2_1 _18031_ (.A(_07600_),
    .B(_07043_),
    .Y(_07601_));
 sky130_fd_sc_hd__nand2_1 _18032_ (.A(_07597_),
    .B(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__inv_2 _18033_ (.A(_07600_),
    .Y(_07603_));
 sky130_fd_sc_hd__nand2_1 _18034_ (.A(_07603_),
    .B(_07048_),
    .Y(_07605_));
 sky130_fd_sc_hd__nand2_1 _18035_ (.A(_07602_),
    .B(_07605_),
    .Y(_07606_));
 sky130_fd_sc_hd__nand2_1 _18036_ (.A(_07002_),
    .B(_07007_),
    .Y(_07607_));
 sky130_fd_sc_hd__nand2_1 _18037_ (.A(_07607_),
    .B(_07008_),
    .Y(_07608_));
 sky130_fd_sc_hd__nand2_1 _18038_ (.A(_07608_),
    .B(_07105_),
    .Y(_07609_));
 sky130_fd_sc_hd__nand3_1 _18039_ (.A(_07607_),
    .B(_07008_),
    .C(_07106_),
    .Y(_07610_));
 sky130_fd_sc_hd__nand2_1 _18040_ (.A(_07609_),
    .B(_07610_),
    .Y(_07611_));
 sky130_fd_sc_hd__nand2_1 _18041_ (.A(_07611_),
    .B(_07031_),
    .Y(_07612_));
 sky130_fd_sc_hd__nand3_1 _18042_ (.A(_07609_),
    .B(_07034_),
    .C(_07610_),
    .Y(_07613_));
 sky130_fd_sc_hd__nand2_1 _18043_ (.A(_07612_),
    .B(_07613_),
    .Y(_07614_));
 sky130_fd_sc_hd__inv_2 _18044_ (.A(_07614_),
    .Y(_07616_));
 sky130_fd_sc_hd__nand2_1 _18045_ (.A(_07606_),
    .B(_07616_),
    .Y(_07617_));
 sky130_fd_sc_hd__nand2_2 _18046_ (.A(_07617_),
    .B(_07613_),
    .Y(_07618_));
 sky130_fd_sc_hd__nand2_1 _18047_ (.A(_07610_),
    .B(_07103_),
    .Y(_07619_));
 sky130_fd_sc_hd__xor2_2 _18048_ (.A(_07094_),
    .B(_07619_),
    .X(_07620_));
 sky130_fd_sc_hd__nand2_1 _18049_ (.A(_07620_),
    .B(_06465_),
    .Y(_07621_));
 sky130_fd_sc_hd__nand2_2 _18050_ (.A(_07618_),
    .B(_07621_),
    .Y(_07622_));
 sky130_fd_sc_hd__or2_1 _18051_ (.A(_06465_),
    .B(_07620_),
    .X(_07623_));
 sky130_fd_sc_hd__nand2_1 _18052_ (.A(_07622_),
    .B(_07623_),
    .Y(_07624_));
 sky130_fd_sc_hd__nor2_1 _18053_ (.A(_07094_),
    .B(_07105_),
    .Y(_07625_));
 sky130_fd_sc_hd__nand3_1 _18054_ (.A(_07607_),
    .B(_07625_),
    .C(_07008_),
    .Y(_07627_));
 sky130_fd_sc_hd__inv_2 _18055_ (.A(_07112_),
    .Y(_07628_));
 sky130_fd_sc_hd__nand2_1 _18056_ (.A(_07627_),
    .B(_07628_),
    .Y(_07629_));
 sky130_fd_sc_hd__nand2_1 _18057_ (.A(_07629_),
    .B(_07081_),
    .Y(_07630_));
 sky130_fd_sc_hd__nand2_1 _18058_ (.A(_07630_),
    .B(_07078_),
    .Y(_07631_));
 sky130_fd_sc_hd__nand2_1 _18059_ (.A(_07631_),
    .B(_07071_),
    .Y(_07632_));
 sky130_fd_sc_hd__nand3_1 _18060_ (.A(_07630_),
    .B(_07070_),
    .C(_07078_),
    .Y(_07633_));
 sky130_fd_sc_hd__nand2_1 _18061_ (.A(_07632_),
    .B(_07633_),
    .Y(_07634_));
 sky130_fd_sc_hd__nand2_1 _18062_ (.A(_07634_),
    .B(_05255_),
    .Y(_07635_));
 sky130_fd_sc_hd__nand3_1 _18063_ (.A(_07627_),
    .B(_07080_),
    .C(_07628_),
    .Y(_07636_));
 sky130_fd_sc_hd__nand2_1 _18064_ (.A(_07630_),
    .B(_07636_),
    .Y(_07638_));
 sky130_fd_sc_hd__nand2_1 _18065_ (.A(_07638_),
    .B(_07024_),
    .Y(_07639_));
 sky130_fd_sc_hd__nand3_2 _18066_ (.A(_07630_),
    .B(_07021_),
    .C(_07636_),
    .Y(_07640_));
 sky130_fd_sc_hd__nand2_1 _18067_ (.A(_07639_),
    .B(_07640_),
    .Y(_07641_));
 sky130_fd_sc_hd__inv_2 _18068_ (.A(_07641_),
    .Y(_07642_));
 sky130_fd_sc_hd__nand3_1 _18069_ (.A(_07632_),
    .B(_05896_),
    .C(_07633_),
    .Y(_07643_));
 sky130_fd_sc_hd__nand3_1 _18070_ (.A(_07635_),
    .B(_07642_),
    .C(_07643_),
    .Y(_07644_));
 sky130_fd_sc_hd__inv_2 _18071_ (.A(_07644_),
    .Y(_07645_));
 sky130_fd_sc_hd__nand2_1 _18072_ (.A(_07624_),
    .B(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__inv_2 _18073_ (.A(_07640_),
    .Y(_07647_));
 sky130_fd_sc_hd__a21boi_1 _18074_ (.A1(_07635_),
    .A2(_07647_),
    .B1_N(_07643_),
    .Y(_07649_));
 sky130_fd_sc_hd__nand2_2 _18075_ (.A(_07646_),
    .B(_07649_),
    .Y(_07650_));
 sky130_fd_sc_hd__nand2_1 _18076_ (.A(_07577_),
    .B(_07569_),
    .Y(_07651_));
 sky130_fd_sc_hd__inv_2 _18077_ (.A(_07651_),
    .Y(_07652_));
 sky130_fd_sc_hd__nand2_1 _18078_ (.A(_07572_),
    .B(_07155_),
    .Y(_07653_));
 sky130_fd_sc_hd__nand2_1 _18079_ (.A(_07574_),
    .B(_07653_),
    .Y(_07654_));
 sky130_fd_sc_hd__inv_4 _18080_ (.A(_07654_),
    .Y(_07655_));
 sky130_fd_sc_hd__nand2_1 _18081_ (.A(_07652_),
    .B(_07655_),
    .Y(_07656_));
 sky130_fd_sc_hd__inv_2 _18082_ (.A(_07656_),
    .Y(_07657_));
 sky130_fd_sc_hd__nand3_1 _18083_ (.A(_07588_),
    .B(_07650_),
    .C(_07657_),
    .Y(_07658_));
 sky130_fd_sc_hd__nand2_2 _18084_ (.A(_07587_),
    .B(_07658_),
    .Y(_07660_));
 sky130_fd_sc_hd__inv_2 _18085_ (.A(_07311_),
    .Y(_07661_));
 sky130_fd_sc_hd__inv_2 _18086_ (.A(_07321_),
    .Y(_07662_));
 sky130_fd_sc_hd__nand2_1 _18087_ (.A(_07218_),
    .B(_07662_),
    .Y(_07663_));
 sky130_fd_sc_hd__nand2_1 _18088_ (.A(_07663_),
    .B(_07320_),
    .Y(_07664_));
 sky130_fd_sc_hd__or2_1 _18089_ (.A(_07661_),
    .B(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__nand2_1 _18090_ (.A(_07664_),
    .B(_07661_),
    .Y(_07666_));
 sky130_fd_sc_hd__nand2_1 _18091_ (.A(_07665_),
    .B(_07666_),
    .Y(_07667_));
 sky130_fd_sc_hd__nand2_1 _18092_ (.A(_07667_),
    .B(_07247_),
    .Y(_07668_));
 sky130_fd_sc_hd__nand3_1 _18093_ (.A(_07665_),
    .B(_07249_),
    .C(_07666_),
    .Y(_07669_));
 sky130_fd_sc_hd__nand2_1 _18094_ (.A(_07668_),
    .B(_07669_),
    .Y(_07671_));
 sky130_fd_sc_hd__inv_2 _18095_ (.A(_07671_),
    .Y(_07672_));
 sky130_fd_sc_hd__or2_1 _18096_ (.A(_07662_),
    .B(_07218_),
    .X(_07673_));
 sky130_fd_sc_hd__nand2_1 _18097_ (.A(_07673_),
    .B(_07663_),
    .Y(_07674_));
 sky130_fd_sc_hd__inv_2 _18098_ (.A(_07674_),
    .Y(_07675_));
 sky130_fd_sc_hd__nand2_1 _18099_ (.A(_07675_),
    .B(_06521_),
    .Y(_07676_));
 sky130_fd_sc_hd__buf_6 _18100_ (.A(_06012_),
    .X(_07677_));
 sky130_fd_sc_hd__nand2_1 _18101_ (.A(_07674_),
    .B(_07677_),
    .Y(_07678_));
 sky130_fd_sc_hd__nand2_1 _18102_ (.A(_07676_),
    .B(_07678_),
    .Y(_07679_));
 sky130_fd_sc_hd__inv_4 _18103_ (.A(_07679_),
    .Y(_07680_));
 sky130_fd_sc_hd__nand2_1 _18104_ (.A(_07672_),
    .B(_07680_),
    .Y(_07682_));
 sky130_fd_sc_hd__inv_4 _18105_ (.A(_07682_),
    .Y(_07683_));
 sky130_fd_sc_hd__nand2_1 _18106_ (.A(_07660_),
    .B(_07683_),
    .Y(_07684_));
 sky130_fd_sc_hd__inv_2 _18107_ (.A(_07676_),
    .Y(_07685_));
 sky130_fd_sc_hd__a21boi_2 _18108_ (.A1(_07668_),
    .A2(_07685_),
    .B1_N(_07669_),
    .Y(_07686_));
 sky130_fd_sc_hd__nand2_1 _18109_ (.A(_07684_),
    .B(_07686_),
    .Y(_07687_));
 sky130_fd_sc_hd__nand2_1 _18110_ (.A(_07218_),
    .B(_07322_),
    .Y(_07688_));
 sky130_fd_sc_hd__inv_2 _18111_ (.A(_07326_),
    .Y(_07689_));
 sky130_fd_sc_hd__nand2_1 _18112_ (.A(_07688_),
    .B(_07689_),
    .Y(_07690_));
 sky130_fd_sc_hd__inv_2 _18113_ (.A(_07302_),
    .Y(_07691_));
 sky130_fd_sc_hd__nand2_1 _18114_ (.A(_07690_),
    .B(_07691_),
    .Y(_07693_));
 sky130_fd_sc_hd__nand3_1 _18115_ (.A(_07688_),
    .B(_07302_),
    .C(_07689_),
    .Y(_07694_));
 sky130_fd_sc_hd__nand2_1 _18116_ (.A(_07693_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__inv_2 _18117_ (.A(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__nand2_1 _18118_ (.A(_07696_),
    .B(_07278_),
    .Y(_07697_));
 sky130_fd_sc_hd__nand2_1 _18119_ (.A(_07695_),
    .B(_07276_),
    .Y(_07698_));
 sky130_fd_sc_hd__nand2_1 _18120_ (.A(_07697_),
    .B(_07698_),
    .Y(_07699_));
 sky130_fd_sc_hd__inv_2 _18121_ (.A(_07699_),
    .Y(_07700_));
 sky130_fd_sc_hd__nand2_1 _18122_ (.A(_07687_),
    .B(_07700_),
    .Y(_07701_));
 sky130_fd_sc_hd__inv_6 _18123_ (.A(_07541_),
    .Y(_07702_));
 sky130_fd_sc_hd__nand3_1 _18124_ (.A(_07684_),
    .B(_07699_),
    .C(_07686_),
    .Y(_07704_));
 sky130_fd_sc_hd__nand3_1 _18125_ (.A(_07701_),
    .B(_07702_),
    .C(_07704_),
    .Y(_07705_));
 sky130_fd_sc_hd__nand2_1 _18126_ (.A(_07542_),
    .B(_07696_),
    .Y(_07706_));
 sky130_fd_sc_hd__nand2_1 _18127_ (.A(_07705_),
    .B(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__nand2_1 _18128_ (.A(_07707_),
    .B(_06554_),
    .Y(_07708_));
 sky130_fd_sc_hd__nand3_1 _18129_ (.A(_07705_),
    .B(_06556_),
    .C(_07706_),
    .Y(_07709_));
 sky130_fd_sc_hd__nand2_1 _18130_ (.A(_07708_),
    .B(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__nand2_1 _18131_ (.A(_07660_),
    .B(_07680_),
    .Y(_07711_));
 sky130_fd_sc_hd__nand2_1 _18132_ (.A(_07711_),
    .B(_07676_),
    .Y(_07712_));
 sky130_fd_sc_hd__nand2_1 _18133_ (.A(_07712_),
    .B(_07672_),
    .Y(_07713_));
 sky130_fd_sc_hd__nand3_1 _18134_ (.A(_07711_),
    .B(_07671_),
    .C(_07676_),
    .Y(_07715_));
 sky130_fd_sc_hd__nand2_1 _18135_ (.A(_07713_),
    .B(_07715_),
    .Y(_07716_));
 sky130_fd_sc_hd__nand2_1 _18136_ (.A(_07716_),
    .B(_07702_),
    .Y(_07717_));
 sky130_fd_sc_hd__nand2_1 _18137_ (.A(_07542_),
    .B(_07667_),
    .Y(_07718_));
 sky130_fd_sc_hd__nand2_1 _18138_ (.A(_07717_),
    .B(_07718_),
    .Y(_07719_));
 sky130_fd_sc_hd__nand2_1 _18139_ (.A(_07719_),
    .B(_06568_),
    .Y(_07720_));
 sky130_fd_sc_hd__nand3_2 _18140_ (.A(_07717_),
    .B(_06570_),
    .C(_07718_),
    .Y(_07721_));
 sky130_fd_sc_hd__nand2_1 _18141_ (.A(_07720_),
    .B(_07721_),
    .Y(_07722_));
 sky130_fd_sc_hd__nor2_1 _18142_ (.A(_07710_),
    .B(_07722_),
    .Y(_07723_));
 sky130_fd_sc_hd__nand2_1 _18143_ (.A(_07657_),
    .B(_07650_),
    .Y(_07724_));
 sky130_fd_sc_hd__nand2_1 _18144_ (.A(_07724_),
    .B(_07579_),
    .Y(_07726_));
 sky130_fd_sc_hd__nand2_1 _18145_ (.A(_07726_),
    .B(_07584_),
    .Y(_07727_));
 sky130_fd_sc_hd__nand2_1 _18146_ (.A(_07727_),
    .B(_07556_),
    .Y(_07728_));
 sky130_fd_sc_hd__nand3_1 _18147_ (.A(_07728_),
    .B(_07558_),
    .C(_07554_),
    .Y(_07729_));
 sky130_fd_sc_hd__nand2_1 _18148_ (.A(_07554_),
    .B(_07558_),
    .Y(_07730_));
 sky130_fd_sc_hd__nand3_1 _18149_ (.A(_07727_),
    .B(_07556_),
    .C(_07730_),
    .Y(_07731_));
 sky130_fd_sc_hd__nand2_1 _18150_ (.A(_07729_),
    .B(_07731_),
    .Y(_07732_));
 sky130_fd_sc_hd__nand2_1 _18151_ (.A(_07732_),
    .B(_07702_),
    .Y(_07733_));
 sky130_fd_sc_hd__nand2_1 _18152_ (.A(_07542_),
    .B(_07553_),
    .Y(_07734_));
 sky130_fd_sc_hd__nand3_1 _18153_ (.A(_07733_),
    .B(_07318_),
    .C(_07734_),
    .Y(_07735_));
 sky130_fd_sc_hd__or2_1 _18154_ (.A(_07680_),
    .B(_07660_),
    .X(_07737_));
 sky130_fd_sc_hd__nand3_1 _18155_ (.A(_07737_),
    .B(_07702_),
    .C(_07711_),
    .Y(_07738_));
 sky130_fd_sc_hd__nand2_1 _18156_ (.A(_07542_),
    .B(_07675_),
    .Y(_07739_));
 sky130_fd_sc_hd__nand3_1 _18157_ (.A(_07738_),
    .B(_06592_),
    .C(_07739_),
    .Y(_07740_));
 sky130_fd_sc_hd__inv_2 _18158_ (.A(_07740_),
    .Y(_07741_));
 sky130_fd_sc_hd__a21o_1 _18159_ (.A1(_07738_),
    .A2(_07739_),
    .B1(_06592_),
    .X(_07742_));
 sky130_fd_sc_hd__o21ai_1 _18160_ (.A1(_07735_),
    .A2(_07741_),
    .B1(_07742_),
    .Y(_07743_));
 sky130_fd_sc_hd__inv_2 _18161_ (.A(_07709_),
    .Y(_07744_));
 sky130_fd_sc_hd__o21ai_1 _18162_ (.A1(_07721_),
    .A2(_07744_),
    .B1(_07708_),
    .Y(_07745_));
 sky130_fd_sc_hd__a21oi_1 _18163_ (.A1(_07723_),
    .A2(_07743_),
    .B1(_07745_),
    .Y(_07746_));
 sky130_fd_sc_hd__inv_2 _18164_ (.A(_07591_),
    .Y(_07748_));
 sky130_fd_sc_hd__nand2_1 _18165_ (.A(_07542_),
    .B(_07748_),
    .Y(_07749_));
 sky130_fd_sc_hd__nand2_1 _18166_ (.A(_07592_),
    .B(_07595_),
    .Y(_07750_));
 sky130_fd_sc_hd__xor2_1 _18167_ (.A(_07594_),
    .B(_07750_),
    .X(_07751_));
 sky130_fd_sc_hd__nand3b_1 _18168_ (.A_N(_07751_),
    .B(_07538_),
    .C(_07540_),
    .Y(_07752_));
 sky130_fd_sc_hd__nand2_1 _18169_ (.A(_07749_),
    .B(_07752_),
    .Y(_07753_));
 sky130_fd_sc_hd__nand2_1 _18170_ (.A(_07753_),
    .B(_05983_),
    .Y(_07754_));
 sky130_fd_sc_hd__nor2_1 _18171_ (.A(_06979_),
    .B(_07383_),
    .Y(_07755_));
 sky130_fd_sc_hd__or2_1 _18172_ (.A(_06607_),
    .B(_07755_),
    .X(_07756_));
 sky130_fd_sc_hd__nand2_1 _18173_ (.A(_07756_),
    .B(_07005_),
    .Y(_07757_));
 sky130_fd_sc_hd__inv_2 _18174_ (.A(_07757_),
    .Y(_07759_));
 sky130_fd_sc_hd__nand2_1 _18175_ (.A(_07541_),
    .B(_07759_),
    .Y(_07760_));
 sky130_fd_sc_hd__nand3_1 _18176_ (.A(_07538_),
    .B(_07540_),
    .C(_07755_),
    .Y(_07761_));
 sky130_fd_sc_hd__nand2_1 _18177_ (.A(_07760_),
    .B(_07761_),
    .Y(_07762_));
 sky130_fd_sc_hd__nand2_1 _18178_ (.A(_07762_),
    .B(_06615_),
    .Y(_07763_));
 sky130_fd_sc_hd__nand2_1 _18179_ (.A(_07754_),
    .B(_07763_),
    .Y(_07764_));
 sky130_fd_sc_hd__inv_2 _18180_ (.A(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__nand3_1 _18181_ (.A(_07760_),
    .B(_06620_),
    .C(_07761_),
    .Y(_07766_));
 sky130_fd_sc_hd__nand3_2 _18182_ (.A(_07542_),
    .B(_06980_),
    .C(_07004_),
    .Y(_07767_));
 sky130_fd_sc_hd__inv_2 _18183_ (.A(_07767_),
    .Y(_07768_));
 sky130_fd_sc_hd__nand3_4 _18184_ (.A(_07763_),
    .B(_07766_),
    .C(_07768_),
    .Y(_07770_));
 sky130_fd_sc_hd__or2_4 _18185_ (.A(_05983_),
    .B(_07753_),
    .X(_07771_));
 sky130_fd_sc_hd__a21boi_2 _18186_ (.A1(_07765_),
    .A2(_07770_),
    .B1_N(_07771_),
    .Y(_07772_));
 sky130_fd_sc_hd__clkinvlp_2 _18187_ (.A(_07638_),
    .Y(_07773_));
 sky130_fd_sc_hd__nand2_1 _18188_ (.A(_07541_),
    .B(_07773_),
    .Y(_07774_));
 sky130_fd_sc_hd__nand2_1 _18189_ (.A(_07624_),
    .B(_07642_),
    .Y(_07775_));
 sky130_fd_sc_hd__nand3_1 _18190_ (.A(_07622_),
    .B(_07641_),
    .C(_07623_),
    .Y(_07776_));
 sky130_fd_sc_hd__nand2_1 _18191_ (.A(_07775_),
    .B(_07776_),
    .Y(_07777_));
 sky130_fd_sc_hd__inv_2 _18192_ (.A(_07777_),
    .Y(_07778_));
 sky130_fd_sc_hd__nand3_1 _18193_ (.A(_07538_),
    .B(_07540_),
    .C(_07778_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand2_1 _18194_ (.A(_07774_),
    .B(_07779_),
    .Y(_07781_));
 sky130_fd_sc_hd__nand2_1 _18195_ (.A(_07781_),
    .B(_06636_),
    .Y(_07782_));
 sky130_fd_sc_hd__nand3_1 _18196_ (.A(_07774_),
    .B(_06639_),
    .C(_07779_),
    .Y(_07783_));
 sky130_fd_sc_hd__nand2_1 _18197_ (.A(_07782_),
    .B(_07783_),
    .Y(_07784_));
 sky130_fd_sc_hd__clkinvlp_2 _18198_ (.A(_07784_),
    .Y(_07785_));
 sky130_fd_sc_hd__nand2_1 _18199_ (.A(_07542_),
    .B(_07620_),
    .Y(_07786_));
 sky130_fd_sc_hd__nand2_1 _18200_ (.A(_07623_),
    .B(_07621_),
    .Y(_07787_));
 sky130_fd_sc_hd__xor2_1 _18201_ (.A(_07618_),
    .B(_07787_),
    .X(_07788_));
 sky130_fd_sc_hd__nand3_1 _18202_ (.A(_07538_),
    .B(_07540_),
    .C(_07788_),
    .Y(_07789_));
 sky130_fd_sc_hd__nand2_1 _18203_ (.A(_07786_),
    .B(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__nand2_1 _18204_ (.A(_07790_),
    .B(_06648_),
    .Y(_07792_));
 sky130_fd_sc_hd__nand3_2 _18205_ (.A(_07786_),
    .B(_06651_),
    .C(_07789_),
    .Y(_07793_));
 sky130_fd_sc_hd__nand2_2 _18206_ (.A(_07792_),
    .B(_07793_),
    .Y(_07794_));
 sky130_fd_sc_hd__inv_2 _18207_ (.A(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__nand2_1 _18208_ (.A(_07785_),
    .B(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__inv_2 _18209_ (.A(_07611_),
    .Y(_07797_));
 sky130_fd_sc_hd__nand2_1 _18210_ (.A(_07541_),
    .B(_07797_),
    .Y(_07798_));
 sky130_fd_sc_hd__or2_1 _18211_ (.A(_07616_),
    .B(_07606_),
    .X(_07799_));
 sky130_fd_sc_hd__nand2_1 _18212_ (.A(_07799_),
    .B(_07617_),
    .Y(_07800_));
 sky130_fd_sc_hd__clkinvlp_2 _18213_ (.A(_07800_),
    .Y(_07801_));
 sky130_fd_sc_hd__nand3_1 _18214_ (.A(_07538_),
    .B(_07540_),
    .C(_07801_),
    .Y(_07803_));
 sky130_fd_sc_hd__nand2_1 _18215_ (.A(_07798_),
    .B(_07803_),
    .Y(_07804_));
 sky130_fd_sc_hd__nand2_1 _18216_ (.A(_07804_),
    .B(_06033_),
    .Y(_07805_));
 sky130_fd_sc_hd__nand3_1 _18217_ (.A(_07798_),
    .B(_07092_),
    .C(_07803_),
    .Y(_07806_));
 sky130_fd_sc_hd__nand2_1 _18218_ (.A(_07805_),
    .B(_07806_),
    .Y(_07807_));
 sky130_fd_sc_hd__inv_2 _18219_ (.A(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__nand2_1 _18220_ (.A(_07541_),
    .B(_07603_),
    .Y(_07809_));
 sky130_fd_sc_hd__nand2_1 _18221_ (.A(_07605_),
    .B(_07601_),
    .Y(_07810_));
 sky130_fd_sc_hd__xnor2_1 _18222_ (.A(_07597_),
    .B(_07810_),
    .Y(_07811_));
 sky130_fd_sc_hd__nand3_1 _18223_ (.A(net135),
    .B(_07540_),
    .C(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__nand2_1 _18224_ (.A(_07809_),
    .B(_07812_),
    .Y(_07814_));
 sky130_fd_sc_hd__nand2_2 _18225_ (.A(_07814_),
    .B(_07102_),
    .Y(_07815_));
 sky130_fd_sc_hd__nand3_1 _18226_ (.A(_07809_),
    .B(_06046_),
    .C(_07812_),
    .Y(_07816_));
 sky130_fd_sc_hd__nand2_2 _18227_ (.A(_07815_),
    .B(_07816_),
    .Y(_07817_));
 sky130_fd_sc_hd__clkinv_1 _18228_ (.A(_07817_),
    .Y(_07818_));
 sky130_fd_sc_hd__nand2_1 _18229_ (.A(_07808_),
    .B(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__nor2_1 _18230_ (.A(_07796_),
    .B(_07819_),
    .Y(_07820_));
 sky130_fd_sc_hd__nand2_1 _18231_ (.A(_07772_),
    .B(_07820_),
    .Y(_07821_));
 sky130_fd_sc_hd__inv_2 _18232_ (.A(_07806_),
    .Y(_07822_));
 sky130_fd_sc_hd__o21ai_2 _18233_ (.A1(_07815_),
    .A2(_07822_),
    .B1(_07805_),
    .Y(_07823_));
 sky130_fd_sc_hd__nor2_1 _18234_ (.A(_07784_),
    .B(_07794_),
    .Y(_07825_));
 sky130_fd_sc_hd__clkinvlp_2 _18235_ (.A(_07783_),
    .Y(_07826_));
 sky130_fd_sc_hd__o21ai_1 _18236_ (.A1(_07793_),
    .A2(_07826_),
    .B1(_07782_),
    .Y(_07827_));
 sky130_fd_sc_hd__a21oi_1 _18237_ (.A1(_07823_),
    .A2(_07825_),
    .B1(_07827_),
    .Y(_07828_));
 sky130_fd_sc_hd__nand2_2 _18238_ (.A(_07821_),
    .B(_07828_),
    .Y(_07829_));
 sky130_fd_sc_hd__nand2_2 _18239_ (.A(_07650_),
    .B(_07655_),
    .Y(_07830_));
 sky130_fd_sc_hd__or2_1 _18240_ (.A(_07655_),
    .B(_07650_),
    .X(_07831_));
 sky130_fd_sc_hd__nand3_1 _18241_ (.A(_07702_),
    .B(_07830_),
    .C(_07831_),
    .Y(_07832_));
 sky130_fd_sc_hd__nand2_1 _18242_ (.A(_07541_),
    .B(_07573_),
    .Y(_07833_));
 sky130_fd_sc_hd__nand2_1 _18243_ (.A(_07832_),
    .B(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__nand2_1 _18244_ (.A(_07834_),
    .B(_06695_),
    .Y(_07836_));
 sky130_fd_sc_hd__nand3_2 _18245_ (.A(_07832_),
    .B(_06697_),
    .C(_07833_),
    .Y(_07837_));
 sky130_fd_sc_hd__nand2_2 _18246_ (.A(_07836_),
    .B(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__inv_2 _18247_ (.A(_07838_),
    .Y(_07839_));
 sky130_fd_sc_hd__nand2_1 _18248_ (.A(_07635_),
    .B(_07643_),
    .Y(_07840_));
 sky130_fd_sc_hd__nand2_1 _18249_ (.A(_07775_),
    .B(_07640_),
    .Y(_07841_));
 sky130_fd_sc_hd__xor2_1 _18250_ (.A(_07840_),
    .B(_07841_),
    .X(_07842_));
 sky130_fd_sc_hd__nand2_1 _18251_ (.A(_07842_),
    .B(_07702_),
    .Y(_07843_));
 sky130_fd_sc_hd__nand2_1 _18252_ (.A(_07542_),
    .B(_07634_),
    .Y(_07844_));
 sky130_fd_sc_hd__nand2_1 _18253_ (.A(_07843_),
    .B(_07844_),
    .Y(_07845_));
 sky130_fd_sc_hd__nand2_1 _18254_ (.A(_07845_),
    .B(_05915_),
    .Y(_07847_));
 sky130_fd_sc_hd__nand3_1 _18255_ (.A(_07843_),
    .B(_08834_),
    .C(_07844_),
    .Y(_07848_));
 sky130_fd_sc_hd__nand2_1 _18256_ (.A(_07847_),
    .B(_07848_),
    .Y(_07849_));
 sky130_fd_sc_hd__inv_2 _18257_ (.A(_07849_),
    .Y(_07850_));
 sky130_fd_sc_hd__nand2_1 _18258_ (.A(_07839_),
    .B(_07850_),
    .Y(_07851_));
 sky130_fd_sc_hd__nand2_1 _18259_ (.A(_07830_),
    .B(_07574_),
    .Y(_07852_));
 sky130_fd_sc_hd__nand2_1 _18260_ (.A(_07852_),
    .B(_07652_),
    .Y(_07853_));
 sky130_fd_sc_hd__nand3_1 _18261_ (.A(_07830_),
    .B(_07651_),
    .C(_07574_),
    .Y(_07854_));
 sky130_fd_sc_hd__nand2_1 _18262_ (.A(_07853_),
    .B(_07854_),
    .Y(_07855_));
 sky130_fd_sc_hd__nand2_1 _18263_ (.A(_07855_),
    .B(_07702_),
    .Y(_07856_));
 sky130_fd_sc_hd__nand2_1 _18264_ (.A(_07542_),
    .B(_07568_),
    .Y(_07858_));
 sky130_fd_sc_hd__nand2_1 _18265_ (.A(_07856_),
    .B(_07858_),
    .Y(_07859_));
 sky130_fd_sc_hd__nand2_1 _18266_ (.A(_07859_),
    .B(_06721_),
    .Y(_07860_));
 sky130_fd_sc_hd__nand3_2 _18267_ (.A(_07856_),
    .B(_06723_),
    .C(_07858_),
    .Y(_07861_));
 sky130_fd_sc_hd__nand2_1 _18268_ (.A(_07860_),
    .B(_07861_),
    .Y(_07862_));
 sky130_fd_sc_hd__or2_1 _18269_ (.A(_07580_),
    .B(_07702_),
    .X(_07863_));
 sky130_fd_sc_hd__nand3_1 _18270_ (.A(_07724_),
    .B(_07583_),
    .C(_07579_),
    .Y(_07864_));
 sky130_fd_sc_hd__nand3_2 _18271_ (.A(_07727_),
    .B(_07702_),
    .C(_07864_),
    .Y(_07865_));
 sky130_fd_sc_hd__nand2_1 _18272_ (.A(_07863_),
    .B(_07865_),
    .Y(_07866_));
 sky130_fd_sc_hd__nand2_1 _18273_ (.A(_07866_),
    .B(_06731_),
    .Y(_07867_));
 sky130_fd_sc_hd__nand3_2 _18274_ (.A(_07863_),
    .B(_07865_),
    .C(_06733_),
    .Y(_07869_));
 sky130_fd_sc_hd__nand2_2 _18275_ (.A(_07867_),
    .B(_07869_),
    .Y(_07870_));
 sky130_fd_sc_hd__nor2_1 _18276_ (.A(_07862_),
    .B(_07870_),
    .Y(_07871_));
 sky130_fd_sc_hd__nor2b_1 _18277_ (.A(_07851_),
    .B_N(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__nand2_1 _18278_ (.A(_07829_),
    .B(_07872_),
    .Y(_07873_));
 sky130_fd_sc_hd__clkinvlp_2 _18279_ (.A(_07837_),
    .Y(_07874_));
 sky130_fd_sc_hd__o21ai_1 _18280_ (.A1(_07848_),
    .A2(_07874_),
    .B1(_07836_),
    .Y(_07875_));
 sky130_fd_sc_hd__inv_2 _18281_ (.A(_07869_),
    .Y(_07876_));
 sky130_fd_sc_hd__o21ai_1 _18282_ (.A1(_07861_),
    .A2(_07876_),
    .B1(_07867_),
    .Y(_07877_));
 sky130_fd_sc_hd__a21oi_1 _18283_ (.A1(_07871_),
    .A2(_07875_),
    .B1(_07877_),
    .Y(_07878_));
 sky130_fd_sc_hd__nand2_2 _18284_ (.A(_07873_),
    .B(_07878_),
    .Y(_07880_));
 sky130_fd_sc_hd__nand2_1 _18285_ (.A(_07733_),
    .B(_07734_),
    .Y(_07881_));
 sky130_fd_sc_hd__nand2_1 _18286_ (.A(_07881_),
    .B(_06159_),
    .Y(_07882_));
 sky130_fd_sc_hd__nand2_1 _18287_ (.A(_07882_),
    .B(_07735_),
    .Y(_07883_));
 sky130_fd_sc_hd__nand2_1 _18288_ (.A(_07742_),
    .B(_07740_),
    .Y(_07884_));
 sky130_fd_sc_hd__nor2_1 _18289_ (.A(_07883_),
    .B(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__nand3_2 _18290_ (.A(_07880_),
    .B(_07723_),
    .C(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__nand2_2 _18291_ (.A(_07746_),
    .B(_07886_),
    .Y(_07887_));
 sky130_fd_sc_hd__nand2_1 _18292_ (.A(_07417_),
    .B(_07419_),
    .Y(_07888_));
 sky130_fd_sc_hd__inv_4 _18293_ (.A(_07888_),
    .Y(_07889_));
 sky130_fd_sc_hd__or2_1 _18294_ (.A(_07889_),
    .B(_07329_),
    .X(_07891_));
 sky130_fd_sc_hd__nand2_1 _18295_ (.A(_07329_),
    .B(_07889_),
    .Y(_07892_));
 sky130_fd_sc_hd__nand2_1 _18296_ (.A(_07891_),
    .B(_07892_),
    .Y(_07893_));
 sky130_fd_sc_hd__inv_2 _18297_ (.A(_07893_),
    .Y(_07894_));
 sky130_fd_sc_hd__nand2_1 _18298_ (.A(_07894_),
    .B(_06207_),
    .Y(_07895_));
 sky130_fd_sc_hd__nand2_1 _18299_ (.A(_07893_),
    .B(_05408_),
    .Y(_07896_));
 sky130_fd_sc_hd__nand2_1 _18300_ (.A(_07895_),
    .B(_07896_),
    .Y(_07897_));
 sky130_fd_sc_hd__inv_2 _18301_ (.A(_07897_),
    .Y(_07898_));
 sky130_fd_sc_hd__nand2_1 _18302_ (.A(_07693_),
    .B(_07301_),
    .Y(_07899_));
 sky130_fd_sc_hd__inv_2 _18303_ (.A(_07290_),
    .Y(_07900_));
 sky130_fd_sc_hd__nand2_1 _18304_ (.A(_07899_),
    .B(_07900_),
    .Y(_07902_));
 sky130_fd_sc_hd__nand3_1 _18305_ (.A(_07693_),
    .B(_07290_),
    .C(_07301_),
    .Y(_07903_));
 sky130_fd_sc_hd__nand2_1 _18306_ (.A(_07902_),
    .B(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__buf_6 _18307_ (.A(_05375_),
    .X(_07905_));
 sky130_fd_sc_hd__nand2_1 _18308_ (.A(_07904_),
    .B(_07905_),
    .Y(_07906_));
 sky130_fd_sc_hd__nand3_1 _18309_ (.A(_07902_),
    .B(_06772_),
    .C(_07903_),
    .Y(_07907_));
 sky130_fd_sc_hd__nand3_1 _18310_ (.A(_07700_),
    .B(_07906_),
    .C(_07907_),
    .Y(_07908_));
 sky130_fd_sc_hd__inv_2 _18311_ (.A(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__nand3_1 _18312_ (.A(_07660_),
    .B(_07683_),
    .C(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__inv_2 _18313_ (.A(_07906_),
    .Y(_07911_));
 sky130_fd_sc_hd__o21ai_1 _18314_ (.A1(_07697_),
    .A2(_07911_),
    .B1(_07907_),
    .Y(_07913_));
 sky130_fd_sc_hd__nor2_1 _18315_ (.A(_07686_),
    .B(_07908_),
    .Y(_07914_));
 sky130_fd_sc_hd__nor2_1 _18316_ (.A(_07913_),
    .B(_07914_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_2 _18317_ (.A(_07910_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__or2_1 _18318_ (.A(_07898_),
    .B(_07916_),
    .X(_07917_));
 sky130_fd_sc_hd__buf_6 _18319_ (.A(_07702_),
    .X(_07918_));
 sky130_fd_sc_hd__nand2_1 _18320_ (.A(_07916_),
    .B(_07898_),
    .Y(_07919_));
 sky130_fd_sc_hd__nand3_1 _18321_ (.A(_07917_),
    .B(_07918_),
    .C(_07919_),
    .Y(_07920_));
 sky130_fd_sc_hd__nand2_1 _18322_ (.A(\div1i.quot[16] ),
    .B(_07894_),
    .Y(_07921_));
 sky130_fd_sc_hd__nand2_1 _18323_ (.A(_07920_),
    .B(_07921_),
    .Y(_07922_));
 sky130_fd_sc_hd__xor2_2 _18324_ (.A(_06754_),
    .B(_07922_),
    .X(_07924_));
 sky130_fd_sc_hd__nand2_1 _18325_ (.A(_07906_),
    .B(_07907_),
    .Y(_07925_));
 sky130_fd_sc_hd__nand2_1 _18326_ (.A(_07701_),
    .B(_07697_),
    .Y(_07926_));
 sky130_fd_sc_hd__xor2_1 _18327_ (.A(_07925_),
    .B(_07926_),
    .X(_07927_));
 sky130_fd_sc_hd__nand2_1 _18328_ (.A(_07927_),
    .B(_07918_),
    .Y(_07928_));
 sky130_fd_sc_hd__nand2_1 _18329_ (.A(\div1i.quot[16] ),
    .B(_07904_),
    .Y(_07929_));
 sky130_fd_sc_hd__nand2_1 _18330_ (.A(_07928_),
    .B(_07929_),
    .Y(_07930_));
 sky130_fd_sc_hd__nand2_1 _18331_ (.A(_07930_),
    .B(_06797_),
    .Y(_07931_));
 sky130_fd_sc_hd__nand3_1 _18332_ (.A(_07928_),
    .B(_06799_),
    .C(_07929_),
    .Y(_07932_));
 sky130_fd_sc_hd__nand2_1 _18333_ (.A(_07931_),
    .B(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__nor2_1 _18334_ (.A(_07924_),
    .B(_07933_),
    .Y(_07935_));
 sky130_fd_sc_hd__nand2_1 _18335_ (.A(_07887_),
    .B(_07935_),
    .Y(_07936_));
 sky130_fd_sc_hd__nand2_1 _18336_ (.A(_07922_),
    .B(_06805_),
    .Y(_07937_));
 sky130_fd_sc_hd__o21a_1 _18337_ (.A1(_07932_),
    .A2(_07924_),
    .B1(_07937_),
    .X(_07938_));
 sky130_fd_sc_hd__nand2_1 _18338_ (.A(_07936_),
    .B(_07938_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_1 _18339_ (.A(_07329_),
    .B(_07421_),
    .Y(_07940_));
 sky130_fd_sc_hd__inv_2 _18340_ (.A(_07423_),
    .Y(_07941_));
 sky130_fd_sc_hd__a21o_1 _18341_ (.A1(_07940_),
    .A2(_07941_),
    .B1(_07402_),
    .X(_07942_));
 sky130_fd_sc_hd__nand3_1 _18342_ (.A(_07940_),
    .B(_07402_),
    .C(_07941_),
    .Y(_07943_));
 sky130_fd_sc_hd__nand2_1 _18343_ (.A(_07942_),
    .B(_07943_),
    .Y(_07944_));
 sky130_fd_sc_hd__inv_2 _18344_ (.A(_07944_),
    .Y(_07946_));
 sky130_fd_sc_hd__nand2_1 _18345_ (.A(_07946_),
    .B(_06819_),
    .Y(_07947_));
 sky130_fd_sc_hd__buf_6 _18346_ (.A(_06737_),
    .X(_07948_));
 sky130_fd_sc_hd__nand2_1 _18347_ (.A(_07944_),
    .B(_07948_),
    .Y(_07949_));
 sky130_fd_sc_hd__nand2_1 _18348_ (.A(_07947_),
    .B(_07949_),
    .Y(_07950_));
 sky130_fd_sc_hd__inv_4 _18349_ (.A(_07950_),
    .Y(_07951_));
 sky130_fd_sc_hd__nand2_1 _18350_ (.A(_07892_),
    .B(_07419_),
    .Y(_07952_));
 sky130_fd_sc_hd__xor2_2 _18351_ (.A(_07411_),
    .B(_07952_),
    .X(_07953_));
 sky130_fd_sc_hd__inv_2 _18352_ (.A(_07953_),
    .Y(_07954_));
 sky130_fd_sc_hd__nand2_1 _18353_ (.A(_07954_),
    .B(_06827_),
    .Y(_07955_));
 sky130_fd_sc_hd__buf_6 _18354_ (.A(_06814_),
    .X(_07957_));
 sky130_fd_sc_hd__nand2_1 _18355_ (.A(_07953_),
    .B(_07957_),
    .Y(_07958_));
 sky130_fd_sc_hd__nand2_1 _18356_ (.A(_07955_),
    .B(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__or2_1 _18357_ (.A(_07897_),
    .B(_07959_),
    .X(_07960_));
 sky130_fd_sc_hd__inv_4 _18358_ (.A(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand2_1 _18359_ (.A(_07916_),
    .B(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__inv_2 _18360_ (.A(_07895_),
    .Y(_07963_));
 sky130_fd_sc_hd__a21boi_1 _18361_ (.A1(_07963_),
    .A2(_07958_),
    .B1_N(_07955_),
    .Y(_07964_));
 sky130_fd_sc_hd__nand2_1 _18362_ (.A(_07962_),
    .B(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__or2_1 _18363_ (.A(_07951_),
    .B(_07965_),
    .X(_07966_));
 sky130_fd_sc_hd__nand2_1 _18364_ (.A(_07965_),
    .B(_07951_),
    .Y(_07968_));
 sky130_fd_sc_hd__nand3_1 _18365_ (.A(_07966_),
    .B(_07918_),
    .C(_07968_),
    .Y(_07969_));
 sky130_fd_sc_hd__nand2_1 _18366_ (.A(\div1i.quot[16] ),
    .B(_07946_),
    .Y(_07970_));
 sky130_fd_sc_hd__nand2_1 _18367_ (.A(_07969_),
    .B(_07970_),
    .Y(_07971_));
 sky130_fd_sc_hd__xor2_2 _18368_ (.A(_06809_),
    .B(_07971_),
    .X(_07972_));
 sky130_fd_sc_hd__nand2_1 _18369_ (.A(_07919_),
    .B(_07895_),
    .Y(_07973_));
 sky130_fd_sc_hd__xor2_1 _18370_ (.A(_07959_),
    .B(_07973_),
    .X(_07974_));
 sky130_fd_sc_hd__nand2_1 _18371_ (.A(_07974_),
    .B(_07918_),
    .Y(_07975_));
 sky130_fd_sc_hd__nand2_1 _18372_ (.A(\div1i.quot[16] ),
    .B(_07953_),
    .Y(_07976_));
 sky130_fd_sc_hd__nand2_1 _18373_ (.A(_07975_),
    .B(_07976_),
    .Y(_07977_));
 sky130_fd_sc_hd__or2_1 _18374_ (.A(_06844_),
    .B(_07977_),
    .X(_07979_));
 sky130_fd_sc_hd__nand2_1 _18375_ (.A(_07977_),
    .B(_06844_),
    .Y(_07980_));
 sky130_fd_sc_hd__nand2_1 _18376_ (.A(_07979_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__nor2_1 _18377_ (.A(_07972_),
    .B(_07981_),
    .Y(_07982_));
 sky130_fd_sc_hd__nand2_1 _18378_ (.A(_07939_),
    .B(_07982_),
    .Y(_07983_));
 sky130_fd_sc_hd__nand2_1 _18379_ (.A(_07971_),
    .B(_06856_),
    .Y(_07984_));
 sky130_fd_sc_hd__o21a_1 _18380_ (.A1(_07979_),
    .A2(_07972_),
    .B1(_07984_),
    .X(_07985_));
 sky130_fd_sc_hd__nand2_2 _18381_ (.A(_07983_),
    .B(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__a21o_1 _18382_ (.A1(_07520_),
    .A2(_07522_),
    .B1(_07426_),
    .X(_07987_));
 sky130_fd_sc_hd__nand3_1 _18383_ (.A(_07426_),
    .B(_07520_),
    .C(_07522_),
    .Y(_07988_));
 sky130_fd_sc_hd__nand2_1 _18384_ (.A(_07987_),
    .B(_07988_),
    .Y(_07990_));
 sky130_fd_sc_hd__or2_1 _18385_ (.A(_07450_),
    .B(_07990_),
    .X(_07991_));
 sky130_fd_sc_hd__nand2_1 _18386_ (.A(_07990_),
    .B(_07450_),
    .Y(_07992_));
 sky130_fd_sc_hd__nand2_1 _18387_ (.A(_07991_),
    .B(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__inv_4 _18388_ (.A(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__nand2_1 _18389_ (.A(_07942_),
    .B(_07401_),
    .Y(_07995_));
 sky130_fd_sc_hd__clkinvlp_2 _18390_ (.A(_07391_),
    .Y(_07996_));
 sky130_fd_sc_hd__nand2_1 _18391_ (.A(_07995_),
    .B(_07996_),
    .Y(_07997_));
 sky130_fd_sc_hd__nand3_1 _18392_ (.A(_07942_),
    .B(_07391_),
    .C(_07401_),
    .Y(_07998_));
 sky130_fd_sc_hd__nand2_1 _18393_ (.A(_07997_),
    .B(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__buf_6 _18394_ (.A(_06704_),
    .X(_08001_));
 sky130_fd_sc_hd__nand2_1 _18395_ (.A(_07999_),
    .B(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__nand3_2 _18396_ (.A(_07997_),
    .B(_06874_),
    .C(_07998_),
    .Y(_08003_));
 sky130_fd_sc_hd__nand3_1 _18397_ (.A(_07951_),
    .B(_08002_),
    .C(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__inv_2 _18398_ (.A(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__nand3_1 _18399_ (.A(_07916_),
    .B(_07961_),
    .C(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__inv_2 _18400_ (.A(_07947_),
    .Y(_08007_));
 sky130_fd_sc_hd__inv_2 _18401_ (.A(_08003_),
    .Y(_08008_));
 sky130_fd_sc_hd__a21o_1 _18402_ (.A1(_08002_),
    .A2(_08007_),
    .B1(_08008_),
    .X(_08009_));
 sky130_fd_sc_hd__nor2_1 _18403_ (.A(_07964_),
    .B(_08004_),
    .Y(_08010_));
 sky130_fd_sc_hd__nor2_1 _18404_ (.A(_08009_),
    .B(_08010_),
    .Y(_08012_));
 sky130_fd_sc_hd__nand2_2 _18405_ (.A(_08006_),
    .B(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__or2_1 _18406_ (.A(_07994_),
    .B(_08013_),
    .X(_08014_));
 sky130_fd_sc_hd__nand2_1 _18407_ (.A(_08013_),
    .B(_07994_),
    .Y(_08015_));
 sky130_fd_sc_hd__nand2_1 _18408_ (.A(_08014_),
    .B(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand2_1 _18409_ (.A(_08016_),
    .B(_07918_),
    .Y(_08017_));
 sky130_fd_sc_hd__nand2_1 _18410_ (.A(\div1i.quot[16] ),
    .B(_07990_),
    .Y(_08018_));
 sky130_fd_sc_hd__nand2_1 _18411_ (.A(_08017_),
    .B(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__buf_6 _18412_ (.A(_10481_),
    .X(_08020_));
 sky130_fd_sc_hd__nand2_1 _18413_ (.A(_08019_),
    .B(_08020_),
    .Y(_08021_));
 sky130_fd_sc_hd__nand3_1 _18414_ (.A(_08017_),
    .B(_06348_),
    .C(_08018_),
    .Y(_08023_));
 sky130_fd_sc_hd__nand2_2 _18415_ (.A(_08021_),
    .B(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__inv_2 _18416_ (.A(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__nand2_1 _18417_ (.A(_08002_),
    .B(_08003_),
    .Y(_08026_));
 sky130_fd_sc_hd__nand2_1 _18418_ (.A(_07968_),
    .B(_07947_),
    .Y(_08027_));
 sky130_fd_sc_hd__xor2_1 _18419_ (.A(_08026_),
    .B(_08027_),
    .X(_08028_));
 sky130_fd_sc_hd__nand2_1 _18420_ (.A(_08028_),
    .B(_07918_),
    .Y(_08029_));
 sky130_fd_sc_hd__nand2_1 _18421_ (.A(_07999_),
    .B(\div1i.quot[16] ),
    .Y(_08030_));
 sky130_fd_sc_hd__nand2_1 _18422_ (.A(_08029_),
    .B(_08030_),
    .Y(_08031_));
 sky130_fd_sc_hd__nand2_1 _18423_ (.A(_08031_),
    .B(_06903_),
    .Y(_08032_));
 sky130_fd_sc_hd__nand3_2 _18424_ (.A(_08029_),
    .B(_06898_),
    .C(_08030_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand3_1 _18425_ (.A(_08025_),
    .B(_08032_),
    .C(_08034_),
    .Y(_08035_));
 sky130_fd_sc_hd__nand2_1 _18426_ (.A(_08015_),
    .B(_07991_),
    .Y(_08036_));
 sky130_fd_sc_hd__nand2_1 _18427_ (.A(_07988_),
    .B(_07520_),
    .Y(_08037_));
 sky130_fd_sc_hd__xor2_2 _18428_ (.A(_07513_),
    .B(_08037_),
    .X(_08038_));
 sky130_fd_sc_hd__inv_2 _18429_ (.A(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__nand2_1 _18430_ (.A(_08039_),
    .B(_07461_),
    .Y(_08040_));
 sky130_fd_sc_hd__buf_6 _18431_ (.A(_06550_),
    .X(_08041_));
 sky130_fd_sc_hd__nand2_1 _18432_ (.A(_08038_),
    .B(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__nand2_1 _18433_ (.A(_08040_),
    .B(_08042_),
    .Y(_08043_));
 sky130_fd_sc_hd__inv_2 _18434_ (.A(_08043_),
    .Y(_08045_));
 sky130_fd_sc_hd__nand2_1 _18435_ (.A(_08036_),
    .B(_08045_),
    .Y(_08046_));
 sky130_fd_sc_hd__nand3_1 _18436_ (.A(_08015_),
    .B(_08043_),
    .C(_07991_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand2_1 _18437_ (.A(_08046_),
    .B(_08047_),
    .Y(_08048_));
 sky130_fd_sc_hd__nand2_1 _18438_ (.A(_08048_),
    .B(_07918_),
    .Y(_08049_));
 sky130_fd_sc_hd__nand2_1 _18439_ (.A(_08038_),
    .B(\div1i.quot[16] ),
    .Y(_08050_));
 sky130_fd_sc_hd__nand2_1 _18440_ (.A(_08049_),
    .B(_08050_),
    .Y(_08051_));
 sky130_fd_sc_hd__nand2_1 _18441_ (.A(_08051_),
    .B(_07474_),
    .Y(_08052_));
 sky130_fd_sc_hd__nand3_2 _18442_ (.A(_08049_),
    .B(_06366_),
    .C(_08050_),
    .Y(_08053_));
 sky130_fd_sc_hd__nand2_1 _18443_ (.A(_08052_),
    .B(_08053_),
    .Y(_08054_));
 sky130_fd_sc_hd__inv_2 _18444_ (.A(_08054_),
    .Y(_08056_));
 sky130_fd_sc_hd__nand2_1 _18445_ (.A(_08045_),
    .B(_07994_),
    .Y(_08057_));
 sky130_fd_sc_hd__inv_2 _18446_ (.A(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__nand2_1 _18447_ (.A(_08013_),
    .B(_08058_),
    .Y(_08059_));
 sky130_fd_sc_hd__o21a_1 _18448_ (.A1(_07991_),
    .A2(_08043_),
    .B1(_08040_),
    .X(_08060_));
 sky130_fd_sc_hd__nand2_1 _18449_ (.A(_08059_),
    .B(_08060_),
    .Y(_08061_));
 sky130_fd_sc_hd__a21oi_1 _18450_ (.A1(_07422_),
    .A2(_07425_),
    .B1(_07523_),
    .Y(_08062_));
 sky130_fd_sc_hd__or2_1 _18451_ (.A(_07526_),
    .B(_08062_),
    .X(_08063_));
 sky130_fd_sc_hd__or2_1 _18452_ (.A(_07478_),
    .B(_08063_),
    .X(_08064_));
 sky130_fd_sc_hd__nand2_1 _18453_ (.A(_08063_),
    .B(_07478_),
    .Y(_08065_));
 sky130_fd_sc_hd__nand2_1 _18454_ (.A(_08064_),
    .B(_08065_),
    .Y(_08067_));
 sky130_fd_sc_hd__inv_2 _18455_ (.A(_08067_),
    .Y(_08068_));
 sky130_fd_sc_hd__nand2_1 _18456_ (.A(_08068_),
    .B(_06936_),
    .Y(_08069_));
 sky130_fd_sc_hd__nand2_1 _18457_ (.A(_08067_),
    .B(_06594_),
    .Y(_08070_));
 sky130_fd_sc_hd__nand2_1 _18458_ (.A(_08069_),
    .B(_08070_),
    .Y(_08071_));
 sky130_fd_sc_hd__clkinvlp_2 _18459_ (.A(_08071_),
    .Y(_08072_));
 sky130_fd_sc_hd__nand2_1 _18460_ (.A(_08061_),
    .B(_08072_),
    .Y(_08073_));
 sky130_fd_sc_hd__nand3_1 _18461_ (.A(_08059_),
    .B(_08060_),
    .C(_08071_),
    .Y(_08074_));
 sky130_fd_sc_hd__nand3_2 _18462_ (.A(_08073_),
    .B(_07918_),
    .C(_08074_),
    .Y(_08075_));
 sky130_fd_sc_hd__nand2_1 _18463_ (.A(_08068_),
    .B(\div1i.quot[16] ),
    .Y(_08076_));
 sky130_fd_sc_hd__nand2_1 _18464_ (.A(_08075_),
    .B(_08076_),
    .Y(_08078_));
 sky130_fd_sc_hd__nand2_2 _18465_ (.A(_08078_),
    .B(_06947_),
    .Y(_08079_));
 sky130_fd_sc_hd__nand3_2 _18466_ (.A(_08075_),
    .B(_06949_),
    .C(_08076_),
    .Y(_08080_));
 sky130_fd_sc_hd__nand2_4 _18467_ (.A(_08080_),
    .B(_08079_),
    .Y(_08081_));
 sky130_fd_sc_hd__inv_2 _18468_ (.A(_08081_),
    .Y(_08082_));
 sky130_fd_sc_hd__nand2_1 _18469_ (.A(_08056_),
    .B(_08082_),
    .Y(_08083_));
 sky130_fd_sc_hd__nor2_1 _18470_ (.A(_08035_),
    .B(_08083_),
    .Y(_08084_));
 sky130_fd_sc_hd__nand2_4 _18471_ (.A(_07986_),
    .B(_08084_),
    .Y(_08085_));
 sky130_fd_sc_hd__o21ai_2 _18472_ (.A1(_08034_),
    .A2(_08024_),
    .B1(_08023_),
    .Y(_08086_));
 sky130_fd_sc_hd__nor2_1 _18473_ (.A(_08081_),
    .B(_08054_),
    .Y(_08087_));
 sky130_fd_sc_hd__o21ai_1 _18474_ (.A1(_08053_),
    .A2(_08081_),
    .B1(_08079_),
    .Y(_08089_));
 sky130_fd_sc_hd__a21oi_2 _18475_ (.A1(_08086_),
    .A2(_08087_),
    .B1(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__nand2_4 _18476_ (.A(_08085_),
    .B(_08090_),
    .Y(_08091_));
 sky130_fd_sc_hd__nand2_1 _18477_ (.A(_08065_),
    .B(_07476_),
    .Y(_08092_));
 sky130_fd_sc_hd__xor2_1 _18478_ (.A(_07503_),
    .B(_08092_),
    .X(_08093_));
 sky130_fd_sc_hd__nand3_1 _18479_ (.A(_08073_),
    .B(_07918_),
    .C(_08069_),
    .Y(_08094_));
 sky130_fd_sc_hd__xnor2_2 _18480_ (.A(_08093_),
    .B(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__nand2_8 _18481_ (.A(_08091_),
    .B(_08095_),
    .Y(_08096_));
 sky130_fd_sc_hd__clkinvlp_2 _18482_ (.A(_08095_),
    .Y(_08097_));
 sky130_fd_sc_hd__nand3_4 _18483_ (.A(_08085_),
    .B(_08090_),
    .C(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__nand2_8 _18484_ (.A(_08096_),
    .B(_08098_),
    .Y(_08100_));
 sky130_fd_sc_hd__buf_8 _18485_ (.A(_08100_),
    .X(_08101_));
 sky130_fd_sc_hd__buf_8 _18486_ (.A(net221),
    .X(\div1i.quot[15] ));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_07763_),
    .B(_07766_),
    .Y(_08102_));
 sky130_fd_sc_hd__nand2_1 _18488_ (.A(_08102_),
    .B(_07767_),
    .Y(_08103_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(_08103_),
    .B(_07770_),
    .Y(_08104_));
 sky130_fd_sc_hd__inv_2 _18490_ (.A(_08104_),
    .Y(_08105_));
 sky130_fd_sc_hd__nand2_1 _18491_ (.A(_08101_),
    .B(_08105_),
    .Y(_08106_));
 sky130_fd_sc_hd__o21ai_1 _18492_ (.A1(_06979_),
    .A2(\div1i.quot[16] ),
    .B1(_06980_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand2_1 _18493_ (.A(_08104_),
    .B(_06982_),
    .Y(_08108_));
 sky130_fd_sc_hd__nand3_1 _18494_ (.A(_08103_),
    .B(_06984_),
    .C(_07770_),
    .Y(_08110_));
 sky130_fd_sc_hd__nand2_1 _18495_ (.A(_08108_),
    .B(_08110_),
    .Y(_08111_));
 sky130_fd_sc_hd__xor2_1 _18496_ (.A(_08107_),
    .B(_08111_),
    .X(_08112_));
 sky130_fd_sc_hd__nand3b_1 _18497_ (.A_N(_08112_),
    .B(_08096_),
    .C(_08098_),
    .Y(_08113_));
 sky130_fd_sc_hd__nand2_1 _18498_ (.A(_08106_),
    .B(_08113_),
    .Y(_08114_));
 sky130_fd_sc_hd__nand2_1 _18499_ (.A(_08114_),
    .B(_05983_),
    .Y(_08115_));
 sky130_fd_sc_hd__nor2_1 _18500_ (.A(_06979_),
    .B(_07918_),
    .Y(_08116_));
 sky130_fd_sc_hd__or2_1 _18501_ (.A(_06607_),
    .B(_08116_),
    .X(_08117_));
 sky130_fd_sc_hd__nand2_1 _18502_ (.A(_08117_),
    .B(_07767_),
    .Y(_08118_));
 sky130_fd_sc_hd__inv_2 _18503_ (.A(_08118_),
    .Y(_08119_));
 sky130_fd_sc_hd__nand2_1 _18504_ (.A(_08101_),
    .B(_08119_),
    .Y(_08121_));
 sky130_fd_sc_hd__nand3_1 _18505_ (.A(_08096_),
    .B(_08098_),
    .C(_08116_),
    .Y(_08122_));
 sky130_fd_sc_hd__nand2_1 _18506_ (.A(_08121_),
    .B(_08122_),
    .Y(_08123_));
 sky130_fd_sc_hd__nand2_2 _18507_ (.A(_08123_),
    .B(_06615_),
    .Y(_08124_));
 sky130_fd_sc_hd__nand2_1 _18508_ (.A(_08115_),
    .B(_08124_),
    .Y(_08125_));
 sky130_fd_sc_hd__inv_2 _18509_ (.A(_08125_),
    .Y(_08126_));
 sky130_fd_sc_hd__nand3_2 _18510_ (.A(_08121_),
    .B(_06620_),
    .C(_08122_),
    .Y(_08127_));
 sky130_fd_sc_hd__nand3_2 _18511_ (.A(_08101_),
    .B(_06980_),
    .C(_07004_),
    .Y(_08128_));
 sky130_fd_sc_hd__inv_2 _18512_ (.A(_08128_),
    .Y(_08129_));
 sky130_fd_sc_hd__nand3_4 _18513_ (.A(_08124_),
    .B(_08127_),
    .C(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__or2_4 _18514_ (.A(_05983_),
    .B(_08114_),
    .X(_08132_));
 sky130_fd_sc_hd__inv_2 _18515_ (.A(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__a21oi_1 _18516_ (.A1(_08126_),
    .A2(_08130_),
    .B1(_08133_),
    .Y(_08134_));
 sky130_fd_sc_hd__nand2_1 _18517_ (.A(_07765_),
    .B(_07770_),
    .Y(_08135_));
 sky130_fd_sc_hd__nand2_1 _18518_ (.A(_08135_),
    .B(_07771_),
    .Y(_08136_));
 sky130_fd_sc_hd__inv_2 _18519_ (.A(_07823_),
    .Y(_08137_));
 sky130_fd_sc_hd__o21ai_1 _18520_ (.A1(_07819_),
    .A2(_08136_),
    .B1(_08137_),
    .Y(_08138_));
 sky130_fd_sc_hd__or2_1 _18521_ (.A(_07795_),
    .B(_08138_),
    .X(_08139_));
 sky130_fd_sc_hd__nand2_1 _18522_ (.A(_08138_),
    .B(_07795_),
    .Y(_08140_));
 sky130_fd_sc_hd__nand2_1 _18523_ (.A(_08139_),
    .B(_08140_),
    .Y(_08141_));
 sky130_fd_sc_hd__inv_2 _18524_ (.A(_08141_),
    .Y(_08143_));
 sky130_fd_sc_hd__nand2_1 _18525_ (.A(_08100_),
    .B(_08143_),
    .Y(_08144_));
 sky130_fd_sc_hd__nand2_1 _18526_ (.A(_08143_),
    .B(_07021_),
    .Y(_08145_));
 sky130_fd_sc_hd__nand2_1 _18527_ (.A(_08141_),
    .B(_07024_),
    .Y(_08146_));
 sky130_fd_sc_hd__nand2_1 _18528_ (.A(_08145_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__inv_2 _18529_ (.A(_08147_),
    .Y(_08148_));
 sky130_fd_sc_hd__nand2_1 _18530_ (.A(_07772_),
    .B(_07818_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand2_1 _18531_ (.A(_08136_),
    .B(_07817_),
    .Y(_08150_));
 sky130_fd_sc_hd__nand2_1 _18532_ (.A(_08149_),
    .B(_08150_),
    .Y(_08151_));
 sky130_fd_sc_hd__nand2_1 _18533_ (.A(_08151_),
    .B(_07031_),
    .Y(_08152_));
 sky130_fd_sc_hd__nand3_1 _18534_ (.A(_08149_),
    .B(_07034_),
    .C(_08150_),
    .Y(_08154_));
 sky130_fd_sc_hd__nand2_1 _18535_ (.A(_08152_),
    .B(_08154_),
    .Y(_08155_));
 sky130_fd_sc_hd__inv_2 _18536_ (.A(_08155_),
    .Y(_08156_));
 sky130_fd_sc_hd__inv_2 _18537_ (.A(_08110_),
    .Y(_08157_));
 sky130_fd_sc_hd__a21o_1 _18538_ (.A1(_08108_),
    .A2(_08107_),
    .B1(_08157_),
    .X(_08158_));
 sky130_fd_sc_hd__nand2_1 _18539_ (.A(_07771_),
    .B(_07754_),
    .Y(_08159_));
 sky130_fd_sc_hd__nand2_1 _18540_ (.A(_07770_),
    .B(_07763_),
    .Y(_08160_));
 sky130_fd_sc_hd__xor2_1 _18541_ (.A(_08159_),
    .B(_08160_),
    .X(_08161_));
 sky130_fd_sc_hd__nand2_1 _18542_ (.A(_08161_),
    .B(_07043_),
    .Y(_08162_));
 sky130_fd_sc_hd__nand2_1 _18543_ (.A(_08158_),
    .B(_08162_),
    .Y(_08163_));
 sky130_fd_sc_hd__inv_2 _18544_ (.A(_08161_),
    .Y(_08165_));
 sky130_fd_sc_hd__nand2_1 _18545_ (.A(_08165_),
    .B(_07048_),
    .Y(_08166_));
 sky130_fd_sc_hd__nand2_1 _18546_ (.A(_08163_),
    .B(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand2_1 _18547_ (.A(_08156_),
    .B(_08167_),
    .Y(_08168_));
 sky130_fd_sc_hd__nand2_1 _18548_ (.A(_08168_),
    .B(_08154_),
    .Y(_08169_));
 sky130_fd_sc_hd__nand2_1 _18549_ (.A(_08149_),
    .B(_07815_),
    .Y(_08170_));
 sky130_fd_sc_hd__xor2_1 _18550_ (.A(_07807_),
    .B(_08170_),
    .X(_08171_));
 sky130_fd_sc_hd__nand2_1 _18551_ (.A(_08171_),
    .B(_06465_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_1 _18552_ (.A(_08169_),
    .B(_08172_),
    .Y(_08173_));
 sky130_fd_sc_hd__inv_2 _18553_ (.A(_08171_),
    .Y(_08174_));
 sky130_fd_sc_hd__clkbuf_8 _18554_ (.A(_05211_),
    .X(_08176_));
 sky130_fd_sc_hd__nand2_1 _18555_ (.A(_08174_),
    .B(_08176_),
    .Y(_08177_));
 sky130_fd_sc_hd__nand2_1 _18556_ (.A(_08173_),
    .B(_08177_),
    .Y(_08178_));
 sky130_fd_sc_hd__or2_1 _18557_ (.A(_08148_),
    .B(_08178_),
    .X(_08179_));
 sky130_fd_sc_hd__nand2_1 _18558_ (.A(_08178_),
    .B(_08148_),
    .Y(_08180_));
 sky130_fd_sc_hd__nand2_1 _18559_ (.A(_08179_),
    .B(_08180_),
    .Y(_08181_));
 sky130_fd_sc_hd__inv_2 _18560_ (.A(_08181_),
    .Y(_08182_));
 sky130_fd_sc_hd__nand3_1 _18561_ (.A(_08096_),
    .B(_08098_),
    .C(_08182_),
    .Y(_08183_));
 sky130_fd_sc_hd__nand2_1 _18562_ (.A(_08144_),
    .B(_08183_),
    .Y(_08184_));
 sky130_fd_sc_hd__nand2_1 _18563_ (.A(_08184_),
    .B(_06636_),
    .Y(_08185_));
 sky130_fd_sc_hd__nand3_1 _18564_ (.A(_08144_),
    .B(_06639_),
    .C(_08183_),
    .Y(_08187_));
 sky130_fd_sc_hd__nand2_1 _18565_ (.A(_08185_),
    .B(_08187_),
    .Y(_08188_));
 sky130_fd_sc_hd__inv_2 _18566_ (.A(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__nand2_1 _18567_ (.A(_08100_),
    .B(_08174_),
    .Y(_08190_));
 sky130_fd_sc_hd__nand2_1 _18568_ (.A(_08177_),
    .B(_08172_),
    .Y(_08191_));
 sky130_fd_sc_hd__xnor2_1 _18569_ (.A(_08169_),
    .B(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__nand3_1 _18570_ (.A(_08096_),
    .B(_08098_),
    .C(_08192_),
    .Y(_08193_));
 sky130_fd_sc_hd__nand2_1 _18571_ (.A(_08190_),
    .B(_08193_),
    .Y(_08194_));
 sky130_fd_sc_hd__nand2_2 _18572_ (.A(_08194_),
    .B(_06651_),
    .Y(_08195_));
 sky130_fd_sc_hd__nand3_1 _18573_ (.A(_08190_),
    .B(_06648_),
    .C(_08193_),
    .Y(_08196_));
 sky130_fd_sc_hd__nand2_1 _18574_ (.A(_08195_),
    .B(_08196_),
    .Y(_08198_));
 sky130_fd_sc_hd__inv_2 _18575_ (.A(_08198_),
    .Y(_08199_));
 sky130_fd_sc_hd__nand2_1 _18576_ (.A(_08189_),
    .B(_08199_),
    .Y(_08200_));
 sky130_fd_sc_hd__inv_2 _18577_ (.A(_08151_),
    .Y(_08201_));
 sky130_fd_sc_hd__nand2_1 _18578_ (.A(_08100_),
    .B(_08201_),
    .Y(_08202_));
 sky130_fd_sc_hd__or2_1 _18579_ (.A(_08167_),
    .B(_08156_),
    .X(_08203_));
 sky130_fd_sc_hd__nand2_1 _18580_ (.A(_08203_),
    .B(_08168_),
    .Y(_08204_));
 sky130_fd_sc_hd__clkinvlp_2 _18581_ (.A(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__nand3_1 _18582_ (.A(_08096_),
    .B(_08098_),
    .C(_08205_),
    .Y(_08206_));
 sky130_fd_sc_hd__nand2_1 _18583_ (.A(_08202_),
    .B(_08206_),
    .Y(_08207_));
 sky130_fd_sc_hd__nand2_1 _18584_ (.A(_08207_),
    .B(_06033_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand3_1 _18585_ (.A(_08202_),
    .B(_07092_),
    .C(_08206_),
    .Y(_08210_));
 sky130_fd_sc_hd__nand2_2 _18586_ (.A(_08209_),
    .B(_08210_),
    .Y(_08211_));
 sky130_fd_sc_hd__inv_2 _18587_ (.A(_08211_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand2_1 _18588_ (.A(_08100_),
    .B(_08165_),
    .Y(_08213_));
 sky130_fd_sc_hd__nand2_1 _18589_ (.A(_08166_),
    .B(_08162_),
    .Y(_08214_));
 sky130_fd_sc_hd__xnor2_1 _18590_ (.A(_08158_),
    .B(_08214_),
    .Y(_08215_));
 sky130_fd_sc_hd__nand3_1 _18591_ (.A(_08096_),
    .B(_08098_),
    .C(_08215_),
    .Y(_08216_));
 sky130_fd_sc_hd__nand2_1 _18592_ (.A(_08213_),
    .B(_08216_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_1 _18593_ (.A(_08217_),
    .B(_07102_),
    .Y(_08218_));
 sky130_fd_sc_hd__nand3_1 _18594_ (.A(_08213_),
    .B(_06046_),
    .C(_08216_),
    .Y(_08220_));
 sky130_fd_sc_hd__nand2_1 _18595_ (.A(_08218_),
    .B(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__inv_2 _18596_ (.A(_08221_),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2_1 _18597_ (.A(_08212_),
    .B(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__nor2_1 _18598_ (.A(_08200_),
    .B(_08223_),
    .Y(_08224_));
 sky130_fd_sc_hd__nand2_1 _18599_ (.A(_08134_),
    .B(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__inv_2 _18600_ (.A(_08210_),
    .Y(_08226_));
 sky130_fd_sc_hd__o21ai_2 _18601_ (.A1(_08218_),
    .A2(_08226_),
    .B1(_08209_),
    .Y(_08227_));
 sky130_fd_sc_hd__nor2_1 _18602_ (.A(_08188_),
    .B(_08198_),
    .Y(_08228_));
 sky130_fd_sc_hd__inv_2 _18603_ (.A(_08187_),
    .Y(_08229_));
 sky130_fd_sc_hd__o21ai_1 _18604_ (.A1(_08195_),
    .A2(_08229_),
    .B1(_08185_),
    .Y(_08231_));
 sky130_fd_sc_hd__a21oi_1 _18605_ (.A1(_08227_),
    .A2(_08228_),
    .B1(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__nand2_2 _18606_ (.A(_08225_),
    .B(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__inv_2 _18607_ (.A(_07851_),
    .Y(_08234_));
 sky130_fd_sc_hd__nand2_1 _18608_ (.A(_07829_),
    .B(_08234_),
    .Y(_08235_));
 sky130_fd_sc_hd__inv_2 _18609_ (.A(_07875_),
    .Y(_08236_));
 sky130_fd_sc_hd__nand2_1 _18610_ (.A(_08235_),
    .B(_08236_),
    .Y(_08237_));
 sky130_fd_sc_hd__inv_2 _18611_ (.A(_07862_),
    .Y(_08238_));
 sky130_fd_sc_hd__nand2_1 _18612_ (.A(_08237_),
    .B(_08238_),
    .Y(_08239_));
 sky130_fd_sc_hd__nand3_1 _18613_ (.A(_08235_),
    .B(_07862_),
    .C(_08236_),
    .Y(_08240_));
 sky130_fd_sc_hd__nand2_1 _18614_ (.A(_08239_),
    .B(_08240_),
    .Y(_08242_));
 sky130_fd_sc_hd__inv_2 _18615_ (.A(_08242_),
    .Y(_08243_));
 sky130_fd_sc_hd__nand2_1 _18616_ (.A(_08243_),
    .B(_07128_),
    .Y(_08244_));
 sky130_fd_sc_hd__nand2_1 _18617_ (.A(_08242_),
    .B(_07130_),
    .Y(_08245_));
 sky130_fd_sc_hd__nand2_1 _18618_ (.A(_08244_),
    .B(_08245_),
    .Y(_08246_));
 sky130_fd_sc_hd__inv_2 _18619_ (.A(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__nand2_1 _18620_ (.A(_08140_),
    .B(_07793_),
    .Y(_08248_));
 sky130_fd_sc_hd__or2_1 _18621_ (.A(_07785_),
    .B(_08248_),
    .X(_08249_));
 sky130_fd_sc_hd__nand2_1 _18622_ (.A(_08248_),
    .B(_07785_),
    .Y(_08250_));
 sky130_fd_sc_hd__nand3_1 _18623_ (.A(_08249_),
    .B(_05896_),
    .C(_08250_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_1 _18624_ (.A(_08251_),
    .B(_08145_),
    .Y(_08253_));
 sky130_fd_sc_hd__inv_2 _18625_ (.A(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__nand2_2 _18626_ (.A(_08180_),
    .B(_08254_),
    .Y(_08255_));
 sky130_fd_sc_hd__nand2_1 _18627_ (.A(_07829_),
    .B(_07850_),
    .Y(_08256_));
 sky130_fd_sc_hd__nand2_2 _18628_ (.A(_08256_),
    .B(_07848_),
    .Y(_08257_));
 sky130_fd_sc_hd__xor2_2 _18629_ (.A(_07838_),
    .B(_08257_),
    .X(_08258_));
 sky130_fd_sc_hd__nand2_2 _18630_ (.A(_08258_),
    .B(_07146_),
    .Y(_08259_));
 sky130_fd_sc_hd__or2_1 _18631_ (.A(_07839_),
    .B(_08257_),
    .X(_08260_));
 sky130_fd_sc_hd__nand2_1 _18632_ (.A(_08257_),
    .B(_07839_),
    .Y(_08261_));
 sky130_fd_sc_hd__nand3_2 _18633_ (.A(_08260_),
    .B(_07149_),
    .C(_08261_),
    .Y(_08262_));
 sky130_fd_sc_hd__or2_1 _18634_ (.A(_07850_),
    .B(_07829_),
    .X(_08264_));
 sky130_fd_sc_hd__nand2_1 _18635_ (.A(_08264_),
    .B(_08256_),
    .Y(_08265_));
 sky130_fd_sc_hd__nand2_1 _18636_ (.A(_08265_),
    .B(_07155_),
    .Y(_08266_));
 sky130_fd_sc_hd__nand3_2 _18637_ (.A(_08264_),
    .B(_07157_),
    .C(_08256_),
    .Y(_08267_));
 sky130_fd_sc_hd__nand2_1 _18638_ (.A(_08266_),
    .B(_08267_),
    .Y(_08268_));
 sky130_fd_sc_hd__inv_2 _18639_ (.A(_08268_),
    .Y(_08269_));
 sky130_fd_sc_hd__nand3_1 _18640_ (.A(_08259_),
    .B(_08262_),
    .C(_08269_),
    .Y(_08270_));
 sky130_fd_sc_hd__inv_2 _18641_ (.A(_08270_),
    .Y(_08271_));
 sky130_fd_sc_hd__nand2_1 _18642_ (.A(_08249_),
    .B(_08250_),
    .Y(_08272_));
 sky130_fd_sc_hd__nand2_2 _18643_ (.A(_08272_),
    .B(_05255_),
    .Y(_08273_));
 sky130_fd_sc_hd__nand3_2 _18644_ (.A(_08255_),
    .B(_08271_),
    .C(_08273_),
    .Y(_08275_));
 sky130_fd_sc_hd__clkinvlp_2 _18645_ (.A(_08267_),
    .Y(_08276_));
 sky130_fd_sc_hd__a21boi_2 _18646_ (.A1(_08259_),
    .A2(_08276_),
    .B1_N(_08262_),
    .Y(_08277_));
 sky130_fd_sc_hd__nand2_1 _18647_ (.A(_08275_),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__or2_1 _18648_ (.A(_08247_),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__inv_6 _18649_ (.A(_08100_),
    .Y(_08280_));
 sky130_fd_sc_hd__nand2_1 _18650_ (.A(_08278_),
    .B(_08247_),
    .Y(_08281_));
 sky130_fd_sc_hd__nand3_1 _18651_ (.A(_08279_),
    .B(_08280_),
    .C(_08281_),
    .Y(_08282_));
 sky130_fd_sc_hd__nand2_1 _18652_ (.A(net221),
    .B(_08243_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand2_1 _18653_ (.A(_08282_),
    .B(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__nand2_1 _18654_ (.A(_08284_),
    .B(_06731_),
    .Y(_08286_));
 sky130_fd_sc_hd__nand3_1 _18655_ (.A(_08282_),
    .B(_06733_),
    .C(_08283_),
    .Y(_08287_));
 sky130_fd_sc_hd__nand2_2 _18656_ (.A(_08286_),
    .B(_08287_),
    .Y(_08288_));
 sky130_fd_sc_hd__nand3_1 _18657_ (.A(_08255_),
    .B(_08273_),
    .C(_08269_),
    .Y(_08289_));
 sky130_fd_sc_hd__nand2_1 _18658_ (.A(_08289_),
    .B(_08267_),
    .Y(_08290_));
 sky130_fd_sc_hd__nand3_1 _18659_ (.A(_08290_),
    .B(_08262_),
    .C(_08259_),
    .Y(_08291_));
 sky130_fd_sc_hd__nand2_1 _18660_ (.A(_08259_),
    .B(_08262_),
    .Y(_08292_));
 sky130_fd_sc_hd__nand3_1 _18661_ (.A(_08289_),
    .B(_08292_),
    .C(_08267_),
    .Y(_08293_));
 sky130_fd_sc_hd__a21o_1 _18662_ (.A1(_08291_),
    .A2(_08293_),
    .B1(_08101_),
    .X(_08294_));
 sky130_fd_sc_hd__nand2_2 _18663_ (.A(net221),
    .B(_08258_),
    .Y(_08295_));
 sky130_fd_sc_hd__nand2_1 _18664_ (.A(_08294_),
    .B(_08295_),
    .Y(_08297_));
 sky130_fd_sc_hd__nand2_1 _18665_ (.A(_08297_),
    .B(_06721_),
    .Y(_08298_));
 sky130_fd_sc_hd__nand3_2 _18666_ (.A(_08294_),
    .B(_06723_),
    .C(_08295_),
    .Y(_08299_));
 sky130_fd_sc_hd__nand2_2 _18667_ (.A(_08298_),
    .B(_08299_),
    .Y(_08300_));
 sky130_fd_sc_hd__nor2_2 _18668_ (.A(_08288_),
    .B(_08300_),
    .Y(_08301_));
 sky130_fd_sc_hd__a21o_1 _18669_ (.A1(_08255_),
    .A2(_08273_),
    .B1(_08269_),
    .X(_08302_));
 sky130_fd_sc_hd__nand3_1 _18670_ (.A(_08280_),
    .B(_08289_),
    .C(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__a21o_1 _18671_ (.A1(_08096_),
    .A2(_08098_),
    .B1(_08265_),
    .X(_08304_));
 sky130_fd_sc_hd__nand2_1 _18672_ (.A(_08303_),
    .B(_08304_),
    .Y(_08305_));
 sky130_fd_sc_hd__nand2_1 _18673_ (.A(_08305_),
    .B(_06695_),
    .Y(_08306_));
 sky130_fd_sc_hd__nand3_1 _18674_ (.A(_08303_),
    .B(_06697_),
    .C(_08304_),
    .Y(_08308_));
 sky130_fd_sc_hd__nand2_1 _18675_ (.A(_08306_),
    .B(_08308_),
    .Y(_08309_));
 sky130_fd_sc_hd__nand2_1 _18676_ (.A(_08273_),
    .B(_08251_),
    .Y(_08310_));
 sky130_fd_sc_hd__nand2_1 _18677_ (.A(_08180_),
    .B(_08145_),
    .Y(_08311_));
 sky130_fd_sc_hd__xor2_1 _18678_ (.A(_08310_),
    .B(_08311_),
    .X(_08312_));
 sky130_fd_sc_hd__nand2_1 _18679_ (.A(_08280_),
    .B(_08312_),
    .Y(_08313_));
 sky130_fd_sc_hd__nand2_1 _18680_ (.A(_08101_),
    .B(_08272_),
    .Y(_08314_));
 sky130_fd_sc_hd__nand2_1 _18681_ (.A(_08313_),
    .B(_08314_),
    .Y(_08315_));
 sky130_fd_sc_hd__or2_4 _18682_ (.A(_05915_),
    .B(_08315_),
    .X(_08316_));
 sky130_fd_sc_hd__nand2_1 _18683_ (.A(_08315_),
    .B(_05915_),
    .Y(_08317_));
 sky130_fd_sc_hd__nand2_1 _18684_ (.A(_08316_),
    .B(_08317_),
    .Y(_08319_));
 sky130_fd_sc_hd__nor2_2 _18685_ (.A(_08309_),
    .B(_08319_),
    .Y(_08320_));
 sky130_fd_sc_hd__nand2_1 _18686_ (.A(_08301_),
    .B(_08320_),
    .Y(_08321_));
 sky130_fd_sc_hd__inv_2 _18687_ (.A(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__nand2_1 _18688_ (.A(_08233_),
    .B(_08322_),
    .Y(_08323_));
 sky130_fd_sc_hd__o21ai_2 _18689_ (.A1(_08316_),
    .A2(_08309_),
    .B1(_08306_),
    .Y(_08324_));
 sky130_fd_sc_hd__o21ai_1 _18690_ (.A1(_08299_),
    .A2(_08288_),
    .B1(_08286_),
    .Y(_08325_));
 sky130_fd_sc_hd__a21oi_1 _18691_ (.A1(_08324_),
    .A2(_08301_),
    .B1(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__nand2_2 _18692_ (.A(_08323_),
    .B(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__inv_2 _18693_ (.A(_08275_),
    .Y(_08328_));
 sky130_fd_sc_hd__nand2_1 _18694_ (.A(_08239_),
    .B(_07861_),
    .Y(_08330_));
 sky130_fd_sc_hd__inv_2 _18695_ (.A(_07870_),
    .Y(_08331_));
 sky130_fd_sc_hd__nand2_1 _18696_ (.A(_08330_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__nand3_1 _18697_ (.A(_08239_),
    .B(_07861_),
    .C(_07870_),
    .Y(_08333_));
 sky130_fd_sc_hd__nand2_1 _18698_ (.A(_08332_),
    .B(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__nand2_1 _18699_ (.A(_08334_),
    .B(_07226_),
    .Y(_08335_));
 sky130_fd_sc_hd__nand3_1 _18700_ (.A(_08332_),
    .B(_07228_),
    .C(_08333_),
    .Y(_08336_));
 sky130_fd_sc_hd__nand3_1 _18701_ (.A(_08247_),
    .B(_08335_),
    .C(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__inv_2 _18702_ (.A(_08337_),
    .Y(_08338_));
 sky130_fd_sc_hd__nand2_1 _18703_ (.A(_08328_),
    .B(_08338_),
    .Y(_08339_));
 sky130_fd_sc_hd__nor2_1 _18704_ (.A(_08277_),
    .B(_08337_),
    .Y(_08341_));
 sky130_fd_sc_hd__nand2_1 _18705_ (.A(_08335_),
    .B(_08336_),
    .Y(_08342_));
 sky130_fd_sc_hd__o21ai_1 _18706_ (.A1(_08244_),
    .A2(_08342_),
    .B1(_08336_),
    .Y(_08343_));
 sky130_fd_sc_hd__nor2_1 _18707_ (.A(_08341_),
    .B(_08343_),
    .Y(_08344_));
 sky130_fd_sc_hd__nand2_2 _18708_ (.A(_08339_),
    .B(_08344_),
    .Y(_08345_));
 sky130_fd_sc_hd__inv_2 _18709_ (.A(_07884_),
    .Y(_08346_));
 sky130_fd_sc_hd__inv_2 _18710_ (.A(_07883_),
    .Y(_08347_));
 sky130_fd_sc_hd__nand2_1 _18711_ (.A(_07880_),
    .B(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nand2_1 _18712_ (.A(_08348_),
    .B(_07735_),
    .Y(_08349_));
 sky130_fd_sc_hd__or2_1 _18713_ (.A(_08346_),
    .B(_08349_),
    .X(_08350_));
 sky130_fd_sc_hd__nand2_1 _18714_ (.A(_08349_),
    .B(_08346_),
    .Y(_08352_));
 sky130_fd_sc_hd__nand2_1 _18715_ (.A(_08350_),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__nand2_1 _18716_ (.A(_08353_),
    .B(_07247_),
    .Y(_08354_));
 sky130_fd_sc_hd__nand3_1 _18717_ (.A(_08350_),
    .B(_07249_),
    .C(_08352_),
    .Y(_08355_));
 sky130_fd_sc_hd__nand2_1 _18718_ (.A(_08354_),
    .B(_08355_),
    .Y(_08356_));
 sky130_fd_sc_hd__inv_2 _18719_ (.A(_08356_),
    .Y(_08357_));
 sky130_fd_sc_hd__or2_1 _18720_ (.A(_08347_),
    .B(_07880_),
    .X(_08358_));
 sky130_fd_sc_hd__nand2_1 _18721_ (.A(_08358_),
    .B(_08348_),
    .Y(_08359_));
 sky130_fd_sc_hd__inv_2 _18722_ (.A(_08359_),
    .Y(_08360_));
 sky130_fd_sc_hd__nand2_1 _18723_ (.A(_08360_),
    .B(_06521_),
    .Y(_08361_));
 sky130_fd_sc_hd__nand2_1 _18724_ (.A(_08359_),
    .B(_07677_),
    .Y(_08363_));
 sky130_fd_sc_hd__nand2_2 _18725_ (.A(_08361_),
    .B(_08363_),
    .Y(_08364_));
 sky130_fd_sc_hd__inv_4 _18726_ (.A(_08364_),
    .Y(_08365_));
 sky130_fd_sc_hd__nand2_1 _18727_ (.A(_08357_),
    .B(_08365_),
    .Y(_08366_));
 sky130_fd_sc_hd__inv_2 _18728_ (.A(_08366_),
    .Y(_08367_));
 sky130_fd_sc_hd__nand2_1 _18729_ (.A(_08345_),
    .B(_08367_),
    .Y(_08368_));
 sky130_fd_sc_hd__inv_2 _18730_ (.A(_08361_),
    .Y(_08369_));
 sky130_fd_sc_hd__a21boi_2 _18731_ (.A1(_08354_),
    .A2(_08369_),
    .B1_N(_08355_),
    .Y(_08370_));
 sky130_fd_sc_hd__nand2_1 _18732_ (.A(_08368_),
    .B(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__nand2_1 _18733_ (.A(_07880_),
    .B(_07885_),
    .Y(_08372_));
 sky130_fd_sc_hd__inv_2 _18734_ (.A(_07743_),
    .Y(_08374_));
 sky130_fd_sc_hd__nand2_1 _18735_ (.A(_08372_),
    .B(_08374_),
    .Y(_08375_));
 sky130_fd_sc_hd__inv_2 _18736_ (.A(_07722_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand2_1 _18737_ (.A(_08375_),
    .B(_08376_),
    .Y(_08377_));
 sky130_fd_sc_hd__nand3_1 _18738_ (.A(_08372_),
    .B(_08374_),
    .C(_07722_),
    .Y(_08378_));
 sky130_fd_sc_hd__nand2_1 _18739_ (.A(_08377_),
    .B(_08378_),
    .Y(_08379_));
 sky130_fd_sc_hd__nand2_1 _18740_ (.A(_08379_),
    .B(_07276_),
    .Y(_08380_));
 sky130_fd_sc_hd__nand3_1 _18741_ (.A(_08377_),
    .B(_08378_),
    .C(_07278_),
    .Y(_08381_));
 sky130_fd_sc_hd__nand2_1 _18742_ (.A(_08380_),
    .B(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__inv_2 _18743_ (.A(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__nand2_1 _18744_ (.A(_08371_),
    .B(_08383_),
    .Y(_08385_));
 sky130_fd_sc_hd__nand3_1 _18745_ (.A(_08368_),
    .B(_08382_),
    .C(_08370_),
    .Y(_08386_));
 sky130_fd_sc_hd__nand3_1 _18746_ (.A(_08385_),
    .B(_08280_),
    .C(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__or2_1 _18747_ (.A(_08379_),
    .B(_08280_),
    .X(_08388_));
 sky130_fd_sc_hd__nand2_1 _18748_ (.A(_08387_),
    .B(_08388_),
    .Y(_08389_));
 sky130_fd_sc_hd__nand2_1 _18749_ (.A(_08389_),
    .B(_06554_),
    .Y(_08390_));
 sky130_fd_sc_hd__nand3_1 _18750_ (.A(_08387_),
    .B(_06556_),
    .C(_08388_),
    .Y(_08391_));
 sky130_fd_sc_hd__nand2_1 _18751_ (.A(_08390_),
    .B(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__nand2_1 _18752_ (.A(_08345_),
    .B(_08365_),
    .Y(_08393_));
 sky130_fd_sc_hd__nand2_1 _18753_ (.A(_08393_),
    .B(_08361_),
    .Y(_08394_));
 sky130_fd_sc_hd__nand2_1 _18754_ (.A(_08394_),
    .B(_08357_),
    .Y(_08396_));
 sky130_fd_sc_hd__nand3_1 _18755_ (.A(_08393_),
    .B(_08356_),
    .C(_08361_),
    .Y(_08397_));
 sky130_fd_sc_hd__nand2_1 _18756_ (.A(_08396_),
    .B(_08397_),
    .Y(_08398_));
 sky130_fd_sc_hd__nand2_1 _18757_ (.A(_08398_),
    .B(_08280_),
    .Y(_08399_));
 sky130_fd_sc_hd__nand2_1 _18758_ (.A(\div1i.quot[15] ),
    .B(_08353_),
    .Y(_08400_));
 sky130_fd_sc_hd__nand2_1 _18759_ (.A(_08399_),
    .B(_08400_),
    .Y(_08401_));
 sky130_fd_sc_hd__nand2_1 _18760_ (.A(_08401_),
    .B(_06568_),
    .Y(_08402_));
 sky130_fd_sc_hd__nand3_2 _18761_ (.A(_08399_),
    .B(_06570_),
    .C(_08400_),
    .Y(_08403_));
 sky130_fd_sc_hd__nand2_1 _18762_ (.A(_08402_),
    .B(_08403_),
    .Y(_08404_));
 sky130_fd_sc_hd__nor2_1 _18763_ (.A(_08392_),
    .B(_08404_),
    .Y(_08405_));
 sky130_fd_sc_hd__or2_1 _18764_ (.A(_08365_),
    .B(_08345_),
    .X(_08407_));
 sky130_fd_sc_hd__nand3_1 _18765_ (.A(_08407_),
    .B(_08280_),
    .C(_08393_),
    .Y(_08408_));
 sky130_fd_sc_hd__nand2_1 _18766_ (.A(net221),
    .B(_08360_),
    .Y(_08409_));
 sky130_fd_sc_hd__nand2_1 _18767_ (.A(_08408_),
    .B(_08409_),
    .Y(_08410_));
 sky130_fd_sc_hd__nand2_1 _18768_ (.A(_08410_),
    .B(_06149_),
    .Y(_08411_));
 sky130_fd_sc_hd__nand3_1 _18769_ (.A(_08408_),
    .B(_06592_),
    .C(_08409_),
    .Y(_08412_));
 sky130_fd_sc_hd__nand2_1 _18770_ (.A(_08411_),
    .B(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__nand2_1 _18771_ (.A(_08281_),
    .B(_08244_),
    .Y(_08414_));
 sky130_fd_sc_hd__xor2_1 _18772_ (.A(_08342_),
    .B(_08414_),
    .X(_08415_));
 sky130_fd_sc_hd__buf_6 _18773_ (.A(_08280_),
    .X(_08416_));
 sky130_fd_sc_hd__nand2_1 _18774_ (.A(_08415_),
    .B(_08416_),
    .Y(_08418_));
 sky130_fd_sc_hd__nand2_1 _18775_ (.A(\div1i.quot[15] ),
    .B(_08334_),
    .Y(_08419_));
 sky130_fd_sc_hd__nand2_1 _18776_ (.A(_08418_),
    .B(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__nand2_1 _18777_ (.A(_08420_),
    .B(_06159_),
    .Y(_08421_));
 sky130_fd_sc_hd__nand3_1 _18778_ (.A(_08418_),
    .B(_07318_),
    .C(_08419_),
    .Y(_08422_));
 sky130_fd_sc_hd__nand2_1 _18779_ (.A(_08421_),
    .B(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__nor2_2 _18780_ (.A(_08413_),
    .B(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__nand2_1 _18781_ (.A(_08405_),
    .B(_08424_),
    .Y(_08425_));
 sky130_fd_sc_hd__inv_2 _18782_ (.A(_08425_),
    .Y(_08426_));
 sky130_fd_sc_hd__nand2_2 _18783_ (.A(_08327_),
    .B(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__o21ai_1 _18784_ (.A1(_08422_),
    .A2(_08413_),
    .B1(_08411_),
    .Y(_08429_));
 sky130_fd_sc_hd__o21ai_1 _18785_ (.A1(_08403_),
    .A2(_08392_),
    .B1(_08390_),
    .Y(_08430_));
 sky130_fd_sc_hd__a21oi_1 _18786_ (.A1(_08405_),
    .A2(_08429_),
    .B1(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__nand2_4 _18787_ (.A(_08427_),
    .B(_08431_),
    .Y(_08432_));
 sky130_fd_sc_hd__nand2_1 _18788_ (.A(_08377_),
    .B(_07721_),
    .Y(_08433_));
 sky130_fd_sc_hd__inv_2 _18789_ (.A(_07710_),
    .Y(_08434_));
 sky130_fd_sc_hd__nand2_1 _18790_ (.A(_08433_),
    .B(_08434_),
    .Y(_08435_));
 sky130_fd_sc_hd__nand3_1 _18791_ (.A(_08377_),
    .B(_07710_),
    .C(_07721_),
    .Y(_08436_));
 sky130_fd_sc_hd__nand2_1 _18792_ (.A(_08435_),
    .B(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand2_1 _18793_ (.A(_08437_),
    .B(_07905_),
    .Y(_08438_));
 sky130_fd_sc_hd__nand3_1 _18794_ (.A(_08435_),
    .B(_06772_),
    .C(_08436_),
    .Y(_08440_));
 sky130_fd_sc_hd__nand3_1 _18795_ (.A(_08438_),
    .B(_08440_),
    .C(_08383_),
    .Y(_08441_));
 sky130_fd_sc_hd__nor2_1 _18796_ (.A(_08441_),
    .B(_08366_),
    .Y(_08442_));
 sky130_fd_sc_hd__nand2_2 _18797_ (.A(_08345_),
    .B(_08442_),
    .Y(_08443_));
 sky130_fd_sc_hd__nor2_1 _18798_ (.A(_08441_),
    .B(_08370_),
    .Y(_08444_));
 sky130_fd_sc_hd__nand2_1 _18799_ (.A(_08438_),
    .B(_08440_),
    .Y(_08445_));
 sky130_fd_sc_hd__o21ai_1 _18800_ (.A1(_08381_),
    .A2(_08445_),
    .B1(_08440_),
    .Y(_08446_));
 sky130_fd_sc_hd__nor2_2 _18801_ (.A(_08444_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__nand2_2 _18802_ (.A(_08447_),
    .B(_08443_),
    .Y(_08448_));
 sky130_fd_sc_hd__clkinvlp_2 _18803_ (.A(_07924_),
    .Y(_08449_));
 sky130_fd_sc_hd__inv_2 _18804_ (.A(_07933_),
    .Y(_08451_));
 sky130_fd_sc_hd__nand2_1 _18805_ (.A(_07887_),
    .B(_08451_),
    .Y(_08452_));
 sky130_fd_sc_hd__nand2_1 _18806_ (.A(_08452_),
    .B(_07932_),
    .Y(_08453_));
 sky130_fd_sc_hd__or2_1 _18807_ (.A(_08449_),
    .B(_08453_),
    .X(_08454_));
 sky130_fd_sc_hd__nand2_1 _18808_ (.A(_08453_),
    .B(_08449_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand2_1 _18809_ (.A(_08454_),
    .B(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__nand2_1 _18810_ (.A(_08456_),
    .B(_07957_),
    .Y(_08457_));
 sky130_fd_sc_hd__nand3_1 _18811_ (.A(_08454_),
    .B(_06827_),
    .C(_08455_),
    .Y(_08458_));
 sky130_fd_sc_hd__nand2_1 _18812_ (.A(_08457_),
    .B(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__or2_1 _18813_ (.A(_08451_),
    .B(_07887_),
    .X(_08460_));
 sky130_fd_sc_hd__nand2_1 _18814_ (.A(_08460_),
    .B(_08452_),
    .Y(_08462_));
 sky130_fd_sc_hd__inv_2 _18815_ (.A(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__nand2_1 _18816_ (.A(_08463_),
    .B(_06207_),
    .Y(_08464_));
 sky130_fd_sc_hd__buf_6 _18817_ (.A(_05408_),
    .X(_08465_));
 sky130_fd_sc_hd__nand2_1 _18818_ (.A(_08462_),
    .B(_08465_),
    .Y(_08466_));
 sky130_fd_sc_hd__nand2_1 _18819_ (.A(_08464_),
    .B(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__inv_2 _18820_ (.A(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__nand2b_1 _18821_ (.A_N(_08459_),
    .B(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__inv_4 _18822_ (.A(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__nand2_1 _18823_ (.A(_08448_),
    .B(_08470_),
    .Y(_08471_));
 sky130_fd_sc_hd__inv_2 _18824_ (.A(_08464_),
    .Y(_08473_));
 sky130_fd_sc_hd__a21boi_2 _18825_ (.A1(_08457_),
    .A2(_08473_),
    .B1_N(_08458_),
    .Y(_08474_));
 sky130_fd_sc_hd__nand2_1 _18826_ (.A(_08471_),
    .B(_08474_),
    .Y(_08475_));
 sky130_fd_sc_hd__inv_2 _18827_ (.A(_07981_),
    .Y(_08476_));
 sky130_fd_sc_hd__nand2_1 _18828_ (.A(_07939_),
    .B(_08476_),
    .Y(_08477_));
 sky130_fd_sc_hd__nand3_1 _18829_ (.A(_07936_),
    .B(_07938_),
    .C(_07981_),
    .Y(_08478_));
 sky130_fd_sc_hd__nand2_1 _18830_ (.A(_08477_),
    .B(_08478_),
    .Y(_08479_));
 sky130_fd_sc_hd__inv_2 _18831_ (.A(_08479_),
    .Y(_08480_));
 sky130_fd_sc_hd__nand2_1 _18832_ (.A(_08480_),
    .B(_06819_),
    .Y(_08481_));
 sky130_fd_sc_hd__nand2_1 _18833_ (.A(_08479_),
    .B(_07948_),
    .Y(_08482_));
 sky130_fd_sc_hd__nand2_1 _18834_ (.A(_08481_),
    .B(_08482_),
    .Y(_08484_));
 sky130_fd_sc_hd__inv_2 _18835_ (.A(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__nand2_1 _18836_ (.A(_08475_),
    .B(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__nand3_1 _18837_ (.A(_08471_),
    .B(_08484_),
    .C(_08474_),
    .Y(_08487_));
 sky130_fd_sc_hd__nand3_1 _18838_ (.A(_08486_),
    .B(_08416_),
    .C(_08487_),
    .Y(_08488_));
 sky130_fd_sc_hd__nand2_1 _18839_ (.A(\div1i.quot[15] ),
    .B(_08480_),
    .Y(_08489_));
 sky130_fd_sc_hd__nand2_1 _18840_ (.A(_08488_),
    .B(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_1 _18841_ (.A(_08490_),
    .B(_06856_),
    .Y(_08491_));
 sky130_fd_sc_hd__nand3_1 _18842_ (.A(_08488_),
    .B(_06809_),
    .C(_08489_),
    .Y(_08492_));
 sky130_fd_sc_hd__nand2_1 _18843_ (.A(_08491_),
    .B(_08492_),
    .Y(_08493_));
 sky130_fd_sc_hd__nand2_1 _18844_ (.A(_08448_),
    .B(_08468_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand2_1 _18845_ (.A(_08495_),
    .B(_08464_),
    .Y(_08496_));
 sky130_fd_sc_hd__xor2_1 _18846_ (.A(_08459_),
    .B(_08496_),
    .X(_08497_));
 sky130_fd_sc_hd__nand2_1 _18847_ (.A(_08497_),
    .B(_08416_),
    .Y(_08498_));
 sky130_fd_sc_hd__nand2_1 _18848_ (.A(\div1i.quot[15] ),
    .B(_08456_),
    .Y(_08499_));
 sky130_fd_sc_hd__nand2_1 _18849_ (.A(_08498_),
    .B(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2_1 _18850_ (.A(_08500_),
    .B(_06844_),
    .Y(_08501_));
 sky130_fd_sc_hd__nand3_2 _18851_ (.A(_08498_),
    .B(_07400_),
    .C(_08499_),
    .Y(_08502_));
 sky130_fd_sc_hd__nand2_1 _18852_ (.A(_08501_),
    .B(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__nor2_1 _18853_ (.A(_08493_),
    .B(_08503_),
    .Y(_08504_));
 sky130_fd_sc_hd__nand3_1 _18854_ (.A(_08443_),
    .B(_08447_),
    .C(_08467_),
    .Y(_08506_));
 sky130_fd_sc_hd__nand3_1 _18855_ (.A(_08495_),
    .B(_08280_),
    .C(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__nand2_1 _18856_ (.A(net221),
    .B(_08463_),
    .Y(_08508_));
 sky130_fd_sc_hd__nand2_1 _18857_ (.A(_08507_),
    .B(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__or2_1 _18858_ (.A(_06805_),
    .B(_08509_),
    .X(_08510_));
 sky130_fd_sc_hd__nand2_1 _18859_ (.A(_08509_),
    .B(_06805_),
    .Y(_08511_));
 sky130_fd_sc_hd__nand2_2 _18860_ (.A(_08510_),
    .B(_08511_),
    .Y(_08512_));
 sky130_fd_sc_hd__nand2_1 _18861_ (.A(_08385_),
    .B(_08381_),
    .Y(_08513_));
 sky130_fd_sc_hd__xor2_1 _18862_ (.A(_08445_),
    .B(_08513_),
    .X(_08514_));
 sky130_fd_sc_hd__nand2_1 _18863_ (.A(_08514_),
    .B(_08416_),
    .Y(_08515_));
 sky130_fd_sc_hd__nand2_1 _18864_ (.A(net222),
    .B(_08437_),
    .Y(_08517_));
 sky130_fd_sc_hd__nand2_1 _18865_ (.A(_08515_),
    .B(_08517_),
    .Y(_08518_));
 sky130_fd_sc_hd__nand2_1 _18866_ (.A(_08518_),
    .B(_06797_),
    .Y(_08519_));
 sky130_fd_sc_hd__nand3_2 _18867_ (.A(_08515_),
    .B(_06799_),
    .C(_08517_),
    .Y(_08520_));
 sky130_fd_sc_hd__nand3b_1 _18868_ (.A_N(_08512_),
    .B(_08519_),
    .C(_08520_),
    .Y(_08521_));
 sky130_fd_sc_hd__inv_2 _18869_ (.A(_08521_),
    .Y(_08522_));
 sky130_fd_sc_hd__nand3_4 _18870_ (.A(_08432_),
    .B(_08504_),
    .C(_08522_),
    .Y(_08523_));
 sky130_fd_sc_hd__inv_2 _18871_ (.A(_08511_),
    .Y(_08524_));
 sky130_fd_sc_hd__o21bai_2 _18872_ (.A1(_08512_),
    .A2(_08520_),
    .B1_N(_08524_),
    .Y(_08525_));
 sky130_fd_sc_hd__o21ai_1 _18873_ (.A1(_08493_),
    .A2(_08502_),
    .B1(_08491_),
    .Y(_08526_));
 sky130_fd_sc_hd__a21oi_1 _18874_ (.A1(_08504_),
    .A2(_08525_),
    .B1(_08526_),
    .Y(_08528_));
 sky130_fd_sc_hd__nand2_4 _18875_ (.A(_08523_),
    .B(_08528_),
    .Y(_08529_));
 sky130_fd_sc_hd__nand2_1 _18876_ (.A(_08477_),
    .B(_07979_),
    .Y(_08530_));
 sky130_fd_sc_hd__inv_2 _18877_ (.A(_07972_),
    .Y(_08531_));
 sky130_fd_sc_hd__nand2_1 _18878_ (.A(_08530_),
    .B(_08531_),
    .Y(_08532_));
 sky130_fd_sc_hd__nand3_1 _18879_ (.A(_08477_),
    .B(_07972_),
    .C(_07979_),
    .Y(_08533_));
 sky130_fd_sc_hd__nand2_1 _18880_ (.A(_08532_),
    .B(_08533_),
    .Y(_08534_));
 sky130_fd_sc_hd__nand2_1 _18881_ (.A(_08534_),
    .B(_08001_),
    .Y(_08535_));
 sky130_fd_sc_hd__nand3_1 _18882_ (.A(_08532_),
    .B(_06874_),
    .C(_08533_),
    .Y(_08536_));
 sky130_fd_sc_hd__nand3_1 _18883_ (.A(_08485_),
    .B(_08535_),
    .C(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__inv_2 _18884_ (.A(_08537_),
    .Y(_08539_));
 sky130_fd_sc_hd__nand3_2 _18885_ (.A(_08448_),
    .B(_08470_),
    .C(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__inv_2 _18886_ (.A(_08535_),
    .Y(_08541_));
 sky130_fd_sc_hd__o21ai_1 _18887_ (.A1(_08481_),
    .A2(_08541_),
    .B1(_08536_),
    .Y(_08542_));
 sky130_fd_sc_hd__nor2_1 _18888_ (.A(_08474_),
    .B(_08537_),
    .Y(_08543_));
 sky130_fd_sc_hd__nor2_1 _18889_ (.A(_08542_),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__nand2_1 _18890_ (.A(_08540_),
    .B(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__inv_2 _18891_ (.A(_07986_),
    .Y(_08546_));
 sky130_fd_sc_hd__nand2_1 _18892_ (.A(_08032_),
    .B(_08034_),
    .Y(_08547_));
 sky130_fd_sc_hd__nand2_1 _18893_ (.A(_08546_),
    .B(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__inv_2 _18894_ (.A(_08547_),
    .Y(_08550_));
 sky130_fd_sc_hd__nand2_1 _18895_ (.A(_07986_),
    .B(_08550_),
    .Y(_08551_));
 sky130_fd_sc_hd__nand2_1 _18896_ (.A(_08548_),
    .B(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand2_1 _18897_ (.A(_08552_),
    .B(_07450_),
    .Y(_08553_));
 sky130_fd_sc_hd__buf_6 _18898_ (.A(_06649_),
    .X(_08554_));
 sky130_fd_sc_hd__nand3_2 _18899_ (.A(_08548_),
    .B(_08554_),
    .C(_08551_),
    .Y(_08555_));
 sky130_fd_sc_hd__nand2_1 _18900_ (.A(_08553_),
    .B(_08555_),
    .Y(_08556_));
 sky130_fd_sc_hd__inv_2 _18901_ (.A(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__nand2_2 _18902_ (.A(_08545_),
    .B(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__nand3_1 _18903_ (.A(_08540_),
    .B(_08544_),
    .C(_08556_),
    .Y(_08559_));
 sky130_fd_sc_hd__nand3_1 _18904_ (.A(_08558_),
    .B(_08559_),
    .C(_08416_),
    .Y(_08561_));
 sky130_fd_sc_hd__or2_1 _18905_ (.A(_08552_),
    .B(_08280_),
    .X(_08562_));
 sky130_fd_sc_hd__nand2_1 _18906_ (.A(_08561_),
    .B(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__or2_1 _18907_ (.A(_06348_),
    .B(_08563_),
    .X(_08564_));
 sky130_fd_sc_hd__nand2_1 _18908_ (.A(_08563_),
    .B(_06348_),
    .Y(_08565_));
 sky130_fd_sc_hd__nand2_1 _18909_ (.A(_08564_),
    .B(_08565_),
    .Y(_08566_));
 sky130_fd_sc_hd__inv_2 _18910_ (.A(_08566_),
    .Y(_08567_));
 sky130_fd_sc_hd__nand2_1 _18911_ (.A(_08535_),
    .B(_08536_),
    .Y(_08568_));
 sky130_fd_sc_hd__nand2_1 _18912_ (.A(_08486_),
    .B(_08481_),
    .Y(_08569_));
 sky130_fd_sc_hd__xor2_1 _18913_ (.A(_08568_),
    .B(_08569_),
    .X(_08570_));
 sky130_fd_sc_hd__nand2_1 _18914_ (.A(_08570_),
    .B(_08416_),
    .Y(_08572_));
 sky130_fd_sc_hd__nand2_1 _18915_ (.A(net222),
    .B(_08534_),
    .Y(_08573_));
 sky130_fd_sc_hd__nand2_1 _18916_ (.A(_08572_),
    .B(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__nand2_1 _18917_ (.A(_08574_),
    .B(_06903_),
    .Y(_08575_));
 sky130_fd_sc_hd__nand3_2 _18918_ (.A(_08572_),
    .B(_06898_),
    .C(_08573_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand3_1 _18919_ (.A(_08567_),
    .B(_08575_),
    .C(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand2_1 _18920_ (.A(_08558_),
    .B(_08555_),
    .Y(_08578_));
 sky130_fd_sc_hd__nand2_1 _18921_ (.A(_08551_),
    .B(_08034_),
    .Y(_08579_));
 sky130_fd_sc_hd__xor2_2 _18922_ (.A(_08024_),
    .B(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__inv_2 _18923_ (.A(_08580_),
    .Y(_08581_));
 sky130_fd_sc_hd__nand2_1 _18924_ (.A(_08581_),
    .B(_07461_),
    .Y(_08583_));
 sky130_fd_sc_hd__nand2_1 _18925_ (.A(_08580_),
    .B(_08041_),
    .Y(_08584_));
 sky130_fd_sc_hd__nand2_1 _18926_ (.A(_08583_),
    .B(_08584_),
    .Y(_08585_));
 sky130_fd_sc_hd__inv_2 _18927_ (.A(_08585_),
    .Y(_08586_));
 sky130_fd_sc_hd__nand2_1 _18928_ (.A(_08578_),
    .B(_08586_),
    .Y(_08587_));
 sky130_fd_sc_hd__nand3_1 _18929_ (.A(_08558_),
    .B(_08585_),
    .C(_08555_),
    .Y(_08588_));
 sky130_fd_sc_hd__nand2_1 _18930_ (.A(_08587_),
    .B(_08588_),
    .Y(_08589_));
 sky130_fd_sc_hd__nand2_1 _18931_ (.A(_08589_),
    .B(_08416_),
    .Y(_08590_));
 sky130_fd_sc_hd__nand2_1 _18932_ (.A(_08580_),
    .B(net222),
    .Y(_08591_));
 sky130_fd_sc_hd__nand2_1 _18933_ (.A(_08590_),
    .B(_08591_),
    .Y(_08592_));
 sky130_fd_sc_hd__nand2_1 _18934_ (.A(_08592_),
    .B(_07474_),
    .Y(_08594_));
 sky130_fd_sc_hd__nand3_1 _18935_ (.A(_08590_),
    .B(_06366_),
    .C(_08591_),
    .Y(_08595_));
 sky130_fd_sc_hd__nand2_1 _18936_ (.A(_08594_),
    .B(_08595_),
    .Y(_08596_));
 sky130_fd_sc_hd__inv_2 _18937_ (.A(_08596_),
    .Y(_08597_));
 sky130_fd_sc_hd__nand3_1 _18938_ (.A(_08583_),
    .B(_08584_),
    .C(_08557_),
    .Y(_08598_));
 sky130_fd_sc_hd__inv_2 _18939_ (.A(_08598_),
    .Y(_08599_));
 sky130_fd_sc_hd__nand2_1 _18940_ (.A(_08599_),
    .B(_08545_),
    .Y(_08600_));
 sky130_fd_sc_hd__inv_2 _18941_ (.A(_08584_),
    .Y(_08601_));
 sky130_fd_sc_hd__o21a_1 _18942_ (.A1(_08555_),
    .A2(_08601_),
    .B1(_08583_),
    .X(_08602_));
 sky130_fd_sc_hd__nand2_1 _18943_ (.A(_08600_),
    .B(_08602_),
    .Y(_08603_));
 sky130_fd_sc_hd__o21bai_1 _18944_ (.A1(_08035_),
    .A2(_08546_),
    .B1_N(_08086_),
    .Y(_08605_));
 sky130_fd_sc_hd__or2_1 _18945_ (.A(_08056_),
    .B(_08605_),
    .X(_08606_));
 sky130_fd_sc_hd__nand2_1 _18946_ (.A(_08605_),
    .B(_08056_),
    .Y(_08607_));
 sky130_fd_sc_hd__nand2_1 _18947_ (.A(_08606_),
    .B(_08607_),
    .Y(_08608_));
 sky130_fd_sc_hd__inv_2 _18948_ (.A(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__nand2_1 _18949_ (.A(_08609_),
    .B(_06936_),
    .Y(_08610_));
 sky130_fd_sc_hd__buf_6 _18950_ (.A(_06594_),
    .X(_08611_));
 sky130_fd_sc_hd__nand2_1 _18951_ (.A(_08608_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__nand2_1 _18952_ (.A(_08610_),
    .B(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__inv_2 _18953_ (.A(_08613_),
    .Y(_08614_));
 sky130_fd_sc_hd__nand2_1 _18954_ (.A(_08603_),
    .B(_08614_),
    .Y(_08616_));
 sky130_fd_sc_hd__nand3_1 _18955_ (.A(_08600_),
    .B(_08602_),
    .C(_08613_),
    .Y(_08617_));
 sky130_fd_sc_hd__nand3_2 _18956_ (.A(_08616_),
    .B(_08617_),
    .C(_08416_),
    .Y(_08618_));
 sky130_fd_sc_hd__nand2_1 _18957_ (.A(_08609_),
    .B(\div1i.quot[15] ),
    .Y(_08619_));
 sky130_fd_sc_hd__nand2_1 _18958_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__nand2_1 _18959_ (.A(_08620_),
    .B(_06947_),
    .Y(_08621_));
 sky130_fd_sc_hd__nand3_2 _18960_ (.A(_08618_),
    .B(_06949_),
    .C(_08619_),
    .Y(_08622_));
 sky130_fd_sc_hd__nand2_2 _18961_ (.A(_08621_),
    .B(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__inv_2 _18962_ (.A(_08623_),
    .Y(_08624_));
 sky130_fd_sc_hd__nand2_1 _18963_ (.A(_08597_),
    .B(_08624_),
    .Y(_08625_));
 sky130_fd_sc_hd__nor2_1 _18964_ (.A(_08577_),
    .B(_08625_),
    .Y(_08627_));
 sky130_fd_sc_hd__nand2_4 _18965_ (.A(_08529_),
    .B(_08627_),
    .Y(_08628_));
 sky130_fd_sc_hd__o21ai_2 _18966_ (.A1(_08566_),
    .A2(_08576_),
    .B1(_08565_),
    .Y(_08629_));
 sky130_fd_sc_hd__nor2_1 _18967_ (.A(_08623_),
    .B(_08596_),
    .Y(_08630_));
 sky130_fd_sc_hd__inv_2 _18968_ (.A(_08622_),
    .Y(_08631_));
 sky130_fd_sc_hd__o21ai_1 _18969_ (.A1(_08595_),
    .A2(_08631_),
    .B1(_08621_),
    .Y(_08632_));
 sky130_fd_sc_hd__a21oi_2 _18970_ (.A1(_08629_),
    .A2(_08630_),
    .B1(_08632_),
    .Y(_08633_));
 sky130_fd_sc_hd__nand2_4 _18971_ (.A(_08633_),
    .B(_08628_),
    .Y(_08634_));
 sky130_fd_sc_hd__nand2_2 _18972_ (.A(_08607_),
    .B(_08053_),
    .Y(_08635_));
 sky130_fd_sc_hd__xor2_4 _18973_ (.A(_08081_),
    .B(_08635_),
    .X(_08636_));
 sky130_fd_sc_hd__nand3_2 _18974_ (.A(_08616_),
    .B(_08416_),
    .C(_08610_),
    .Y(_08638_));
 sky130_fd_sc_hd__xnor2_4 _18975_ (.A(_08636_),
    .B(_08638_),
    .Y(_08639_));
 sky130_fd_sc_hd__nand2_8 _18976_ (.A(_08634_),
    .B(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__clkinvlp_2 _18977_ (.A(_08639_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand3_4 _18978_ (.A(_08628_),
    .B(_08633_),
    .C(_08641_),
    .Y(_08642_));
 sky130_fd_sc_hd__nand2_8 _18979_ (.A(_08642_),
    .B(_08640_),
    .Y(_08643_));
 sky130_fd_sc_hd__buf_8 _18980_ (.A(_08643_),
    .X(_08644_));
 sky130_fd_sc_hd__buf_6 _18981_ (.A(net229),
    .X(\div1i.quot[14] ));
 sky130_fd_sc_hd__nand2_1 _18982_ (.A(_08233_),
    .B(_08320_),
    .Y(_08645_));
 sky130_fd_sc_hd__inv_2 _18983_ (.A(_08324_),
    .Y(_08646_));
 sky130_fd_sc_hd__nand2_1 _18984_ (.A(_08645_),
    .B(_08646_),
    .Y(_08648_));
 sky130_fd_sc_hd__inv_2 _18985_ (.A(_08300_),
    .Y(_08649_));
 sky130_fd_sc_hd__nand2_1 _18986_ (.A(_08648_),
    .B(_08649_),
    .Y(_08650_));
 sky130_fd_sc_hd__nand2_1 _18987_ (.A(_08650_),
    .B(_08299_),
    .Y(_08651_));
 sky130_fd_sc_hd__inv_2 _18988_ (.A(_08288_),
    .Y(_08652_));
 sky130_fd_sc_hd__nand2_1 _18989_ (.A(_08651_),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__nand3_1 _18990_ (.A(_08650_),
    .B(_08299_),
    .C(_08288_),
    .Y(_08654_));
 sky130_fd_sc_hd__nand2_1 _18991_ (.A(_08653_),
    .B(_08654_),
    .Y(_08655_));
 sky130_fd_sc_hd__nand2_1 _18992_ (.A(_08655_),
    .B(_07226_),
    .Y(_08656_));
 sky130_fd_sc_hd__nand3_1 _18993_ (.A(_08645_),
    .B(_08300_),
    .C(_08646_),
    .Y(_08657_));
 sky130_fd_sc_hd__nand3_2 _18994_ (.A(_08650_),
    .B(_07128_),
    .C(_08657_),
    .Y(_08659_));
 sky130_fd_sc_hd__inv_2 _18995_ (.A(_08659_),
    .Y(_08660_));
 sky130_fd_sc_hd__nand3_2 _18996_ (.A(_08653_),
    .B(_07228_),
    .C(_08654_),
    .Y(_08661_));
 sky130_fd_sc_hd__nand3_1 _18997_ (.A(_08656_),
    .B(_08660_),
    .C(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__nand2_1 _18998_ (.A(_08662_),
    .B(_08661_),
    .Y(_08663_));
 sky130_fd_sc_hd__inv_2 _18999_ (.A(_08319_),
    .Y(_08664_));
 sky130_fd_sc_hd__nand2_1 _19000_ (.A(_08233_),
    .B(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__nand2_1 _19001_ (.A(_08665_),
    .B(_08316_),
    .Y(_08666_));
 sky130_fd_sc_hd__inv_2 _19002_ (.A(_08309_),
    .Y(_08667_));
 sky130_fd_sc_hd__nand2_1 _19003_ (.A(_08666_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__nand3_1 _19004_ (.A(_08665_),
    .B(_08309_),
    .C(_08316_),
    .Y(_08670_));
 sky130_fd_sc_hd__nand2_1 _19005_ (.A(_08668_),
    .B(_08670_),
    .Y(_08671_));
 sky130_fd_sc_hd__nand2_1 _19006_ (.A(_08671_),
    .B(_07146_),
    .Y(_08672_));
 sky130_fd_sc_hd__or2_1 _19007_ (.A(_08664_),
    .B(_08233_),
    .X(_08673_));
 sky130_fd_sc_hd__nand2_1 _19008_ (.A(_08673_),
    .B(_08665_),
    .Y(_08674_));
 sky130_fd_sc_hd__inv_2 _19009_ (.A(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__nand2_1 _19010_ (.A(_08675_),
    .B(_07157_),
    .Y(_08676_));
 sky130_fd_sc_hd__inv_2 _19011_ (.A(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__inv_2 _19012_ (.A(_08671_),
    .Y(_08678_));
 sky130_fd_sc_hd__nand2_1 _19013_ (.A(_08678_),
    .B(_07149_),
    .Y(_08679_));
 sky130_fd_sc_hd__inv_2 _19014_ (.A(_08679_),
    .Y(_08681_));
 sky130_fd_sc_hd__a21oi_1 _19015_ (.A1(_08672_),
    .A2(_08677_),
    .B1(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__nand2_1 _19016_ (.A(_08650_),
    .B(_08657_),
    .Y(_08683_));
 sky130_fd_sc_hd__nand2_1 _19017_ (.A(_08683_),
    .B(_07130_),
    .Y(_08684_));
 sky130_fd_sc_hd__nand2_1 _19018_ (.A(_08684_),
    .B(_08659_),
    .Y(_08685_));
 sky130_fd_sc_hd__inv_2 _19019_ (.A(_08685_),
    .Y(_08686_));
 sky130_fd_sc_hd__nand3_1 _19020_ (.A(_08656_),
    .B(_08686_),
    .C(_08661_),
    .Y(_08687_));
 sky130_fd_sc_hd__nor2_1 _19021_ (.A(_08682_),
    .B(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__nor2_1 _19022_ (.A(_08663_),
    .B(_08688_),
    .Y(_08689_));
 sky130_fd_sc_hd__inv_2 _19023_ (.A(_08687_),
    .Y(_08690_));
 sky130_fd_sc_hd__nand2_1 _19024_ (.A(_08124_),
    .B(_08127_),
    .Y(_08692_));
 sky130_fd_sc_hd__nand2_1 _19025_ (.A(_08692_),
    .B(_08128_),
    .Y(_08693_));
 sky130_fd_sc_hd__nand2_1 _19026_ (.A(_08693_),
    .B(_08130_),
    .Y(_08694_));
 sky130_fd_sc_hd__nand2_1 _19027_ (.A(_08694_),
    .B(_06982_),
    .Y(_08695_));
 sky130_fd_sc_hd__o21ai_2 _19028_ (.A1(_06979_),
    .A2(net222),
    .B1(_06980_),
    .Y(_08696_));
 sky130_fd_sc_hd__nand3_1 _19029_ (.A(_08693_),
    .B(_06984_),
    .C(_08130_),
    .Y(_08697_));
 sky130_fd_sc_hd__inv_2 _19030_ (.A(_08697_),
    .Y(_08698_));
 sky130_fd_sc_hd__a21o_1 _19031_ (.A1(_08695_),
    .A2(_08696_),
    .B1(_08698_),
    .X(_08699_));
 sky130_fd_sc_hd__nand2_1 _19032_ (.A(_08132_),
    .B(_08115_),
    .Y(_08700_));
 sky130_fd_sc_hd__nand2_1 _19033_ (.A(_08130_),
    .B(_08124_),
    .Y(_08701_));
 sky130_fd_sc_hd__xor2_2 _19034_ (.A(_08700_),
    .B(_08701_),
    .X(_08703_));
 sky130_fd_sc_hd__nand2_1 _19035_ (.A(_08703_),
    .B(_07043_),
    .Y(_08704_));
 sky130_fd_sc_hd__nand2_1 _19036_ (.A(_08699_),
    .B(_08704_),
    .Y(_08705_));
 sky130_fd_sc_hd__inv_2 _19037_ (.A(_08703_),
    .Y(_08706_));
 sky130_fd_sc_hd__nand2_1 _19038_ (.A(_08706_),
    .B(_07048_),
    .Y(_08707_));
 sky130_fd_sc_hd__nand2_1 _19039_ (.A(_08705_),
    .B(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__nand2_1 _19040_ (.A(_08126_),
    .B(_08130_),
    .Y(_08709_));
 sky130_fd_sc_hd__nand2_1 _19041_ (.A(_08709_),
    .B(_08132_),
    .Y(_08710_));
 sky130_fd_sc_hd__nand2_1 _19042_ (.A(_08710_),
    .B(_08221_),
    .Y(_08711_));
 sky130_fd_sc_hd__nand3_2 _19043_ (.A(_08709_),
    .B(_08132_),
    .C(_08222_),
    .Y(_08712_));
 sky130_fd_sc_hd__nand2_1 _19044_ (.A(_08711_),
    .B(_08712_),
    .Y(_08714_));
 sky130_fd_sc_hd__nand2_1 _19045_ (.A(_08714_),
    .B(_07031_),
    .Y(_08715_));
 sky130_fd_sc_hd__nand3_1 _19046_ (.A(_08711_),
    .B(_07034_),
    .C(_08712_),
    .Y(_08716_));
 sky130_fd_sc_hd__nand2_1 _19047_ (.A(_08715_),
    .B(_08716_),
    .Y(_08717_));
 sky130_fd_sc_hd__inv_2 _19048_ (.A(_08717_),
    .Y(_08718_));
 sky130_fd_sc_hd__nand2_1 _19049_ (.A(_08708_),
    .B(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__nand2_1 _19050_ (.A(_08719_),
    .B(_08716_),
    .Y(_08720_));
 sky130_fd_sc_hd__nand2_1 _19051_ (.A(_08712_),
    .B(_08218_),
    .Y(_08721_));
 sky130_fd_sc_hd__xor2_2 _19052_ (.A(_08211_),
    .B(_08721_),
    .X(_08722_));
 sky130_fd_sc_hd__nand2_1 _19053_ (.A(_08722_),
    .B(_06465_),
    .Y(_08723_));
 sky130_fd_sc_hd__nand2_1 _19054_ (.A(_08720_),
    .B(_08723_),
    .Y(_08725_));
 sky130_fd_sc_hd__or2_1 _19055_ (.A(_06465_),
    .B(_08722_),
    .X(_08726_));
 sky130_fd_sc_hd__nand2_1 _19056_ (.A(_08725_),
    .B(_08726_),
    .Y(_08727_));
 sky130_fd_sc_hd__nor2_1 _19057_ (.A(_08211_),
    .B(_08221_),
    .Y(_08728_));
 sky130_fd_sc_hd__nand3_1 _19058_ (.A(_08709_),
    .B(_08728_),
    .C(_08132_),
    .Y(_08729_));
 sky130_fd_sc_hd__inv_2 _19059_ (.A(_08227_),
    .Y(_08730_));
 sky130_fd_sc_hd__nand2_1 _19060_ (.A(_08729_),
    .B(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__nand2_2 _19061_ (.A(_08731_),
    .B(_08199_),
    .Y(_08732_));
 sky130_fd_sc_hd__nand2_1 _19062_ (.A(_08732_),
    .B(_08195_),
    .Y(_08733_));
 sky130_fd_sc_hd__nand2_1 _19063_ (.A(_08733_),
    .B(_08189_),
    .Y(_08734_));
 sky130_fd_sc_hd__nand3_1 _19064_ (.A(_08732_),
    .B(_08188_),
    .C(_08195_),
    .Y(_08736_));
 sky130_fd_sc_hd__nand2_1 _19065_ (.A(_08734_),
    .B(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__buf_6 _19066_ (.A(_05255_),
    .X(_08738_));
 sky130_fd_sc_hd__nand2_1 _19067_ (.A(_08737_),
    .B(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__nand3_1 _19068_ (.A(_08729_),
    .B(_08198_),
    .C(_08730_),
    .Y(_08740_));
 sky130_fd_sc_hd__nand2_1 _19069_ (.A(_08732_),
    .B(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__nand2_1 _19070_ (.A(_08741_),
    .B(_07024_),
    .Y(_08742_));
 sky130_fd_sc_hd__nand3_2 _19071_ (.A(_08732_),
    .B(_07021_),
    .C(_08740_),
    .Y(_08743_));
 sky130_fd_sc_hd__nand2_1 _19072_ (.A(_08742_),
    .B(_08743_),
    .Y(_08744_));
 sky130_fd_sc_hd__inv_2 _19073_ (.A(_08744_),
    .Y(_08745_));
 sky130_fd_sc_hd__nand3_1 _19074_ (.A(_08734_),
    .B(_05896_),
    .C(_08736_),
    .Y(_08747_));
 sky130_fd_sc_hd__nand3_1 _19075_ (.A(_08739_),
    .B(_08745_),
    .C(_08747_),
    .Y(_08748_));
 sky130_fd_sc_hd__inv_2 _19076_ (.A(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand2_1 _19077_ (.A(_08727_),
    .B(_08749_),
    .Y(_08750_));
 sky130_fd_sc_hd__inv_2 _19078_ (.A(_08743_),
    .Y(_08751_));
 sky130_fd_sc_hd__a21boi_1 _19079_ (.A1(_08739_),
    .A2(_08751_),
    .B1_N(_08747_),
    .Y(_08752_));
 sky130_fd_sc_hd__nand2_1 _19080_ (.A(_08750_),
    .B(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__nand2_1 _19081_ (.A(_08679_),
    .B(_08672_),
    .Y(_08754_));
 sky130_fd_sc_hd__inv_2 _19082_ (.A(_08754_),
    .Y(_08755_));
 sky130_fd_sc_hd__nand2_1 _19083_ (.A(_08674_),
    .B(_07155_),
    .Y(_08756_));
 sky130_fd_sc_hd__nand2_1 _19084_ (.A(_08676_),
    .B(_08756_),
    .Y(_08758_));
 sky130_fd_sc_hd__inv_4 _19085_ (.A(_08758_),
    .Y(_08759_));
 sky130_fd_sc_hd__nand2_1 _19086_ (.A(_08755_),
    .B(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__inv_2 _19087_ (.A(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__nand3_1 _19088_ (.A(_08690_),
    .B(_08753_),
    .C(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__nand2_2 _19089_ (.A(_08689_),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__inv_2 _19090_ (.A(_08413_),
    .Y(_08764_));
 sky130_fd_sc_hd__inv_2 _19091_ (.A(_08423_),
    .Y(_08765_));
 sky130_fd_sc_hd__nand2_1 _19092_ (.A(_08327_),
    .B(_08765_),
    .Y(_08766_));
 sky130_fd_sc_hd__nand2_1 _19093_ (.A(_08766_),
    .B(_08422_),
    .Y(_08767_));
 sky130_fd_sc_hd__or2_1 _19094_ (.A(_08764_),
    .B(_08767_),
    .X(_08769_));
 sky130_fd_sc_hd__nand2_1 _19095_ (.A(_08767_),
    .B(_08764_),
    .Y(_08770_));
 sky130_fd_sc_hd__nand2_1 _19096_ (.A(_08769_),
    .B(_08770_),
    .Y(_08771_));
 sky130_fd_sc_hd__nand2_1 _19097_ (.A(_08771_),
    .B(_07247_),
    .Y(_08772_));
 sky130_fd_sc_hd__nand3_1 _19098_ (.A(_08769_),
    .B(_07249_),
    .C(_08770_),
    .Y(_08773_));
 sky130_fd_sc_hd__nand2_1 _19099_ (.A(_08772_),
    .B(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__inv_2 _19100_ (.A(_08774_),
    .Y(_08775_));
 sky130_fd_sc_hd__or2_1 _19101_ (.A(_08765_),
    .B(_08327_),
    .X(_08776_));
 sky130_fd_sc_hd__nand2_1 _19102_ (.A(_08776_),
    .B(_08766_),
    .Y(_08777_));
 sky130_fd_sc_hd__inv_2 _19103_ (.A(_08777_),
    .Y(_08778_));
 sky130_fd_sc_hd__nand2_1 _19104_ (.A(_08778_),
    .B(_06521_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand2_1 _19105_ (.A(_08777_),
    .B(_07677_),
    .Y(_08781_));
 sky130_fd_sc_hd__nand2_1 _19106_ (.A(_08780_),
    .B(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__inv_2 _19107_ (.A(_08782_),
    .Y(_08783_));
 sky130_fd_sc_hd__nand2_1 _19108_ (.A(_08775_),
    .B(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__inv_2 _19109_ (.A(_08784_),
    .Y(_08785_));
 sky130_fd_sc_hd__nand2_1 _19110_ (.A(_08763_),
    .B(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__inv_2 _19111_ (.A(_08780_),
    .Y(_08787_));
 sky130_fd_sc_hd__a21boi_2 _19112_ (.A1(_08772_),
    .A2(_08787_),
    .B1_N(_08773_),
    .Y(_08788_));
 sky130_fd_sc_hd__nand2_1 _19113_ (.A(_08786_),
    .B(_08788_),
    .Y(_08789_));
 sky130_fd_sc_hd__nand2_1 _19114_ (.A(_08327_),
    .B(_08424_),
    .Y(_08791_));
 sky130_fd_sc_hd__inv_2 _19115_ (.A(_08429_),
    .Y(_08792_));
 sky130_fd_sc_hd__nand2_1 _19116_ (.A(_08791_),
    .B(_08792_),
    .Y(_08793_));
 sky130_fd_sc_hd__inv_2 _19117_ (.A(_08404_),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_1 _19118_ (.A(_08793_),
    .B(_08794_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand3_1 _19119_ (.A(_08791_),
    .B(_08404_),
    .C(_08792_),
    .Y(_08796_));
 sky130_fd_sc_hd__nand2_1 _19120_ (.A(_08795_),
    .B(_08796_),
    .Y(_08797_));
 sky130_fd_sc_hd__inv_2 _19121_ (.A(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__nand2_1 _19122_ (.A(_08798_),
    .B(_07278_),
    .Y(_08799_));
 sky130_fd_sc_hd__nand2_1 _19123_ (.A(_08797_),
    .B(_07276_),
    .Y(_08800_));
 sky130_fd_sc_hd__nand2_1 _19124_ (.A(_08799_),
    .B(_08800_),
    .Y(_08802_));
 sky130_fd_sc_hd__inv_2 _19125_ (.A(_08802_),
    .Y(_08803_));
 sky130_fd_sc_hd__nand2_1 _19126_ (.A(_08789_),
    .B(_08803_),
    .Y(_08804_));
 sky130_fd_sc_hd__inv_6 _19127_ (.A(_08643_),
    .Y(_08805_));
 sky130_fd_sc_hd__nand3_1 _19128_ (.A(_08786_),
    .B(_08802_),
    .C(_08788_),
    .Y(_08806_));
 sky130_fd_sc_hd__nand3_1 _19129_ (.A(_08804_),
    .B(_08805_),
    .C(_08806_),
    .Y(_08807_));
 sky130_fd_sc_hd__nand2_1 _19130_ (.A(net229),
    .B(_08798_),
    .Y(_08808_));
 sky130_fd_sc_hd__nand2_1 _19131_ (.A(_08807_),
    .B(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__nand2_1 _19132_ (.A(_08809_),
    .B(_06554_),
    .Y(_08810_));
 sky130_fd_sc_hd__nand3_1 _19133_ (.A(_08807_),
    .B(_06556_),
    .C(_08808_),
    .Y(_08811_));
 sky130_fd_sc_hd__nand2_1 _19134_ (.A(_08810_),
    .B(_08811_),
    .Y(_08813_));
 sky130_fd_sc_hd__nand2_1 _19135_ (.A(_08763_),
    .B(_08783_),
    .Y(_08814_));
 sky130_fd_sc_hd__nand2_1 _19136_ (.A(_08814_),
    .B(_08780_),
    .Y(_08815_));
 sky130_fd_sc_hd__nand2_1 _19137_ (.A(_08815_),
    .B(_08775_),
    .Y(_08816_));
 sky130_fd_sc_hd__nand3_1 _19138_ (.A(_08814_),
    .B(_08774_),
    .C(_08780_),
    .Y(_08817_));
 sky130_fd_sc_hd__nand2_1 _19139_ (.A(_08816_),
    .B(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__nand2_1 _19140_ (.A(_08818_),
    .B(_08805_),
    .Y(_08819_));
 sky130_fd_sc_hd__nand2_1 _19141_ (.A(net229),
    .B(_08771_),
    .Y(_08820_));
 sky130_fd_sc_hd__nand2_1 _19142_ (.A(_08819_),
    .B(_08820_),
    .Y(_08821_));
 sky130_fd_sc_hd__nand2_1 _19143_ (.A(_08821_),
    .B(_06568_),
    .Y(_08822_));
 sky130_fd_sc_hd__nand3_2 _19144_ (.A(_08819_),
    .B(_06570_),
    .C(_08820_),
    .Y(_08824_));
 sky130_fd_sc_hd__nand2_1 _19145_ (.A(_08822_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__nor2_1 _19146_ (.A(_08813_),
    .B(_08825_),
    .Y(_08826_));
 sky130_fd_sc_hd__nand2_1 _19147_ (.A(_08761_),
    .B(_08753_),
    .Y(_08827_));
 sky130_fd_sc_hd__nand2_1 _19148_ (.A(_08827_),
    .B(_08682_),
    .Y(_08828_));
 sky130_fd_sc_hd__nand2_1 _19149_ (.A(_08828_),
    .B(_08686_),
    .Y(_08829_));
 sky130_fd_sc_hd__nand2_1 _19150_ (.A(_08829_),
    .B(_08659_),
    .Y(_08830_));
 sky130_fd_sc_hd__nand3_1 _19151_ (.A(_08830_),
    .B(_08661_),
    .C(_08656_),
    .Y(_08831_));
 sky130_fd_sc_hd__nand2_1 _19152_ (.A(_08656_),
    .B(_08661_),
    .Y(_08832_));
 sky130_fd_sc_hd__nand3_1 _19153_ (.A(_08829_),
    .B(_08659_),
    .C(_08832_),
    .Y(_08833_));
 sky130_fd_sc_hd__nand2_1 _19154_ (.A(_08831_),
    .B(_08833_),
    .Y(_08835_));
 sky130_fd_sc_hd__nand2_1 _19155_ (.A(_08835_),
    .B(_08805_),
    .Y(_08836_));
 sky130_fd_sc_hd__nand2_1 _19156_ (.A(net229),
    .B(_08655_),
    .Y(_08837_));
 sky130_fd_sc_hd__nand3_2 _19157_ (.A(_08836_),
    .B(_07318_),
    .C(_08837_),
    .Y(_08838_));
 sky130_fd_sc_hd__or2_1 _19158_ (.A(_08783_),
    .B(_08763_),
    .X(_08839_));
 sky130_fd_sc_hd__nand3_1 _19159_ (.A(_08839_),
    .B(_08805_),
    .C(_08814_),
    .Y(_08840_));
 sky130_fd_sc_hd__nand2_1 _19160_ (.A(net229),
    .B(_08778_),
    .Y(_08841_));
 sky130_fd_sc_hd__nand3_1 _19161_ (.A(_08840_),
    .B(_06592_),
    .C(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__inv_2 _19162_ (.A(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__a21o_1 _19163_ (.A1(_08840_),
    .A2(_08841_),
    .B1(_06592_),
    .X(_08844_));
 sky130_fd_sc_hd__o21ai_2 _19164_ (.A1(_08838_),
    .A2(_08843_),
    .B1(_08844_),
    .Y(_08846_));
 sky130_fd_sc_hd__inv_2 _19165_ (.A(_08811_),
    .Y(_08847_));
 sky130_fd_sc_hd__o21ai_1 _19166_ (.A1(_08824_),
    .A2(_08847_),
    .B1(_08810_),
    .Y(_08848_));
 sky130_fd_sc_hd__a21oi_1 _19167_ (.A1(_08826_),
    .A2(_08846_),
    .B1(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__inv_2 _19168_ (.A(_08694_),
    .Y(_08850_));
 sky130_fd_sc_hd__nand2_1 _19169_ (.A(_08644_),
    .B(_08850_),
    .Y(_08851_));
 sky130_fd_sc_hd__nand2_1 _19170_ (.A(_08695_),
    .B(_08697_),
    .Y(_08852_));
 sky130_fd_sc_hd__xor2_1 _19171_ (.A(_08696_),
    .B(_08852_),
    .X(_08853_));
 sky130_fd_sc_hd__nand3b_1 _19172_ (.A_N(_08853_),
    .B(_08640_),
    .C(_08642_),
    .Y(_08854_));
 sky130_fd_sc_hd__nand2_1 _19173_ (.A(_08851_),
    .B(_08854_),
    .Y(_08855_));
 sky130_fd_sc_hd__buf_6 _19174_ (.A(_05983_),
    .X(_08857_));
 sky130_fd_sc_hd__nand2_1 _19175_ (.A(_08855_),
    .B(_08857_),
    .Y(_08858_));
 sky130_fd_sc_hd__nor2_1 _19176_ (.A(_06979_),
    .B(_08416_),
    .Y(_08859_));
 sky130_fd_sc_hd__or2_1 _19177_ (.A(_06607_),
    .B(_08859_),
    .X(_08860_));
 sky130_fd_sc_hd__nand2_1 _19178_ (.A(_08860_),
    .B(_08128_),
    .Y(_08861_));
 sky130_fd_sc_hd__inv_2 _19179_ (.A(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__nand2_1 _19180_ (.A(_08643_),
    .B(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__nand3_1 _19181_ (.A(_08640_),
    .B(_08642_),
    .C(_08859_),
    .Y(_08864_));
 sky130_fd_sc_hd__nand2_1 _19182_ (.A(_08863_),
    .B(_08864_),
    .Y(_08865_));
 sky130_fd_sc_hd__nand2_1 _19183_ (.A(_08865_),
    .B(_06615_),
    .Y(_08866_));
 sky130_fd_sc_hd__nand2_1 _19184_ (.A(_08858_),
    .B(_08866_),
    .Y(_08868_));
 sky130_fd_sc_hd__inv_2 _19185_ (.A(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__nand3_1 _19186_ (.A(_08863_),
    .B(_06620_),
    .C(_08864_),
    .Y(_08870_));
 sky130_fd_sc_hd__nand3_2 _19187_ (.A(_08644_),
    .B(_06980_),
    .C(_07004_),
    .Y(_08871_));
 sky130_fd_sc_hd__inv_2 _19188_ (.A(_08871_),
    .Y(_08872_));
 sky130_fd_sc_hd__nand3_2 _19189_ (.A(_08866_),
    .B(_08870_),
    .C(_08872_),
    .Y(_08873_));
 sky130_fd_sc_hd__or2_4 _19190_ (.A(_08857_),
    .B(_08855_),
    .X(_08874_));
 sky130_fd_sc_hd__a21boi_1 _19191_ (.A1(_08869_),
    .A2(_08873_),
    .B1_N(_08874_),
    .Y(_08875_));
 sky130_fd_sc_hd__clkinvlp_2 _19192_ (.A(_08741_),
    .Y(_08876_));
 sky130_fd_sc_hd__nand2_1 _19193_ (.A(_08643_),
    .B(_08876_),
    .Y(_08877_));
 sky130_fd_sc_hd__nand2_1 _19194_ (.A(_08727_),
    .B(_08745_),
    .Y(_08879_));
 sky130_fd_sc_hd__nand3_1 _19195_ (.A(_08725_),
    .B(_08744_),
    .C(_08726_),
    .Y(_08880_));
 sky130_fd_sc_hd__nand2_1 _19196_ (.A(_08879_),
    .B(_08880_),
    .Y(_08881_));
 sky130_fd_sc_hd__inv_2 _19197_ (.A(_08881_),
    .Y(_08882_));
 sky130_fd_sc_hd__nand3_1 _19198_ (.A(_08640_),
    .B(_08642_),
    .C(_08882_),
    .Y(_08883_));
 sky130_fd_sc_hd__nand2_1 _19199_ (.A(_08877_),
    .B(_08883_),
    .Y(_08884_));
 sky130_fd_sc_hd__nand2_1 _19200_ (.A(_08884_),
    .B(_06636_),
    .Y(_08885_));
 sky130_fd_sc_hd__nand3_1 _19201_ (.A(_08877_),
    .B(_06639_),
    .C(_08883_),
    .Y(_08886_));
 sky130_fd_sc_hd__nand2_1 _19202_ (.A(_08885_),
    .B(_08886_),
    .Y(_08887_));
 sky130_fd_sc_hd__clkinvlp_2 _19203_ (.A(_08887_),
    .Y(_08888_));
 sky130_fd_sc_hd__nand2_1 _19204_ (.A(_08644_),
    .B(_08722_),
    .Y(_08890_));
 sky130_fd_sc_hd__nand2_1 _19205_ (.A(_08726_),
    .B(_08723_),
    .Y(_08891_));
 sky130_fd_sc_hd__xor2_1 _19206_ (.A(_08720_),
    .B(_08891_),
    .X(_08892_));
 sky130_fd_sc_hd__nand3_1 _19207_ (.A(_08640_),
    .B(_08642_),
    .C(_08892_),
    .Y(_08893_));
 sky130_fd_sc_hd__nand2_1 _19208_ (.A(_08890_),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__nand2_1 _19209_ (.A(_08894_),
    .B(_06648_),
    .Y(_08895_));
 sky130_fd_sc_hd__nand3_2 _19210_ (.A(_08890_),
    .B(_06651_),
    .C(_08893_),
    .Y(_08896_));
 sky130_fd_sc_hd__nand2_2 _19211_ (.A(_08896_),
    .B(_08895_),
    .Y(_08897_));
 sky130_fd_sc_hd__inv_2 _19212_ (.A(_08897_),
    .Y(_08898_));
 sky130_fd_sc_hd__nand2_1 _19213_ (.A(_08888_),
    .B(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__inv_2 _19214_ (.A(_08714_),
    .Y(_08901_));
 sky130_fd_sc_hd__nand2_1 _19215_ (.A(_08643_),
    .B(_08901_),
    .Y(_08902_));
 sky130_fd_sc_hd__or2_1 _19216_ (.A(_08718_),
    .B(_08708_),
    .X(_08903_));
 sky130_fd_sc_hd__nand2_1 _19217_ (.A(_08903_),
    .B(_08719_),
    .Y(_08904_));
 sky130_fd_sc_hd__clkinvlp_2 _19218_ (.A(_08904_),
    .Y(_08905_));
 sky130_fd_sc_hd__nand3_1 _19219_ (.A(_08640_),
    .B(_08642_),
    .C(_08905_),
    .Y(_08906_));
 sky130_fd_sc_hd__nand2_1 _19220_ (.A(_08902_),
    .B(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__nand2_1 _19221_ (.A(_08907_),
    .B(_06033_),
    .Y(_08908_));
 sky130_fd_sc_hd__nand3_1 _19222_ (.A(_08902_),
    .B(_07092_),
    .C(_08906_),
    .Y(_08909_));
 sky130_fd_sc_hd__nand2_1 _19223_ (.A(_08908_),
    .B(_08909_),
    .Y(_08910_));
 sky130_fd_sc_hd__clkinvlp_2 _19224_ (.A(_08910_),
    .Y(_08912_));
 sky130_fd_sc_hd__nand2_1 _19225_ (.A(_08643_),
    .B(_08706_),
    .Y(_08913_));
 sky130_fd_sc_hd__nand2_1 _19226_ (.A(_08707_),
    .B(_08704_),
    .Y(_08914_));
 sky130_fd_sc_hd__xnor2_1 _19227_ (.A(_08699_),
    .B(_08914_),
    .Y(_08915_));
 sky130_fd_sc_hd__nand3_1 _19228_ (.A(_08640_),
    .B(_08642_),
    .C(_08915_),
    .Y(_08916_));
 sky130_fd_sc_hd__nand2_1 _19229_ (.A(_08913_),
    .B(_08916_),
    .Y(_08917_));
 sky130_fd_sc_hd__nand2_1 _19230_ (.A(_08917_),
    .B(_07102_),
    .Y(_08918_));
 sky130_fd_sc_hd__nand3_1 _19231_ (.A(_08913_),
    .B(_06046_),
    .C(_08916_),
    .Y(_08919_));
 sky130_fd_sc_hd__nand2_1 _19232_ (.A(_08918_),
    .B(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__inv_2 _19233_ (.A(_08920_),
    .Y(_08921_));
 sky130_fd_sc_hd__nand2_1 _19234_ (.A(_08912_),
    .B(_08921_),
    .Y(_08923_));
 sky130_fd_sc_hd__nor2_1 _19235_ (.A(_08899_),
    .B(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__nand2_1 _19236_ (.A(_08875_),
    .B(_08924_),
    .Y(_08925_));
 sky130_fd_sc_hd__inv_2 _19237_ (.A(_08909_),
    .Y(_08926_));
 sky130_fd_sc_hd__o21ai_2 _19238_ (.A1(_08918_),
    .A2(_08926_),
    .B1(_08908_),
    .Y(_08927_));
 sky130_fd_sc_hd__nor2_1 _19239_ (.A(_08887_),
    .B(_08897_),
    .Y(_08928_));
 sky130_fd_sc_hd__clkinvlp_2 _19240_ (.A(_08886_),
    .Y(_08929_));
 sky130_fd_sc_hd__o21ai_1 _19241_ (.A1(_08896_),
    .A2(_08929_),
    .B1(_08885_),
    .Y(_08930_));
 sky130_fd_sc_hd__a21oi_1 _19242_ (.A1(_08927_),
    .A2(_08928_),
    .B1(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__nand2_2 _19243_ (.A(_08925_),
    .B(_08931_),
    .Y(_08932_));
 sky130_fd_sc_hd__nand2_1 _19244_ (.A(_08753_),
    .B(_08759_),
    .Y(_08934_));
 sky130_fd_sc_hd__or2_1 _19245_ (.A(_08759_),
    .B(_08753_),
    .X(_08935_));
 sky130_fd_sc_hd__nand3_1 _19246_ (.A(_08805_),
    .B(_08934_),
    .C(_08935_),
    .Y(_08936_));
 sky130_fd_sc_hd__nand2_1 _19247_ (.A(_08643_),
    .B(_08675_),
    .Y(_08937_));
 sky130_fd_sc_hd__nand2_1 _19248_ (.A(_08936_),
    .B(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__nand2_1 _19249_ (.A(_08938_),
    .B(_06695_),
    .Y(_08939_));
 sky130_fd_sc_hd__nand3_1 _19250_ (.A(_08936_),
    .B(_06697_),
    .C(_08937_),
    .Y(_08940_));
 sky130_fd_sc_hd__nand2_1 _19251_ (.A(_08939_),
    .B(_08940_),
    .Y(_08941_));
 sky130_fd_sc_hd__inv_2 _19252_ (.A(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__nand2_1 _19253_ (.A(_08739_),
    .B(_08747_),
    .Y(_08943_));
 sky130_fd_sc_hd__nand2_1 _19254_ (.A(_08879_),
    .B(_08743_),
    .Y(_08945_));
 sky130_fd_sc_hd__xor2_1 _19255_ (.A(_08943_),
    .B(_08945_),
    .X(_08946_));
 sky130_fd_sc_hd__nand2_1 _19256_ (.A(_08946_),
    .B(_08805_),
    .Y(_08947_));
 sky130_fd_sc_hd__nand2_1 _19257_ (.A(_08644_),
    .B(_08737_),
    .Y(_08948_));
 sky130_fd_sc_hd__nand2_1 _19258_ (.A(_08947_),
    .B(_08948_),
    .Y(_08949_));
 sky130_fd_sc_hd__nand2_1 _19259_ (.A(_08949_),
    .B(_05915_),
    .Y(_08950_));
 sky130_fd_sc_hd__buf_6 _19260_ (.A(_08834_),
    .X(_08951_));
 sky130_fd_sc_hd__nand3_2 _19261_ (.A(_08947_),
    .B(_08951_),
    .C(_08948_),
    .Y(_08952_));
 sky130_fd_sc_hd__nand2_1 _19262_ (.A(_08950_),
    .B(_08952_),
    .Y(_08953_));
 sky130_fd_sc_hd__inv_2 _19263_ (.A(_08953_),
    .Y(_08954_));
 sky130_fd_sc_hd__nand2_1 _19264_ (.A(_08942_),
    .B(_08954_),
    .Y(_08956_));
 sky130_fd_sc_hd__nand2_1 _19265_ (.A(_08934_),
    .B(_08676_),
    .Y(_08957_));
 sky130_fd_sc_hd__nand2_1 _19266_ (.A(_08957_),
    .B(_08755_),
    .Y(_08958_));
 sky130_fd_sc_hd__nand3_1 _19267_ (.A(_08934_),
    .B(_08754_),
    .C(_08676_),
    .Y(_08959_));
 sky130_fd_sc_hd__nand2_1 _19268_ (.A(_08958_),
    .B(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__nand2_1 _19269_ (.A(_08960_),
    .B(_08805_),
    .Y(_08961_));
 sky130_fd_sc_hd__nand2_1 _19270_ (.A(_08644_),
    .B(_08671_),
    .Y(_08962_));
 sky130_fd_sc_hd__nand2_1 _19271_ (.A(_08961_),
    .B(_08962_),
    .Y(_08963_));
 sky130_fd_sc_hd__nand2_1 _19272_ (.A(_08963_),
    .B(_06721_),
    .Y(_08964_));
 sky130_fd_sc_hd__nand3_2 _19273_ (.A(_08961_),
    .B(_06723_),
    .C(_08962_),
    .Y(_08965_));
 sky130_fd_sc_hd__nand2_1 _19274_ (.A(_08964_),
    .B(_08965_),
    .Y(_08967_));
 sky130_fd_sc_hd__or2_1 _19275_ (.A(_08683_),
    .B(_08805_),
    .X(_08968_));
 sky130_fd_sc_hd__nand3_1 _19276_ (.A(_08827_),
    .B(_08685_),
    .C(_08682_),
    .Y(_08969_));
 sky130_fd_sc_hd__nand3_1 _19277_ (.A(_08829_),
    .B(_08805_),
    .C(_08969_),
    .Y(_08970_));
 sky130_fd_sc_hd__nand2_1 _19278_ (.A(_08968_),
    .B(_08970_),
    .Y(_08971_));
 sky130_fd_sc_hd__nand2_1 _19279_ (.A(_08971_),
    .B(_06731_),
    .Y(_08972_));
 sky130_fd_sc_hd__nand3_1 _19280_ (.A(_08968_),
    .B(_08970_),
    .C(_06733_),
    .Y(_08973_));
 sky130_fd_sc_hd__nand2_2 _19281_ (.A(_08972_),
    .B(_08973_),
    .Y(_08974_));
 sky130_fd_sc_hd__nor2_1 _19282_ (.A(_08967_),
    .B(_08974_),
    .Y(_08975_));
 sky130_fd_sc_hd__nor2b_1 _19283_ (.A(_08956_),
    .B_N(_08975_),
    .Y(_08976_));
 sky130_fd_sc_hd__nand2_1 _19284_ (.A(_08932_),
    .B(_08976_),
    .Y(_08978_));
 sky130_fd_sc_hd__inv_2 _19285_ (.A(_08940_),
    .Y(_08979_));
 sky130_fd_sc_hd__o21ai_2 _19286_ (.A1(_08952_),
    .A2(_08979_),
    .B1(_08939_),
    .Y(_08980_));
 sky130_fd_sc_hd__inv_2 _19287_ (.A(_08973_),
    .Y(_08981_));
 sky130_fd_sc_hd__o21ai_1 _19288_ (.A1(_08965_),
    .A2(_08981_),
    .B1(_08972_),
    .Y(_08982_));
 sky130_fd_sc_hd__a21oi_1 _19289_ (.A1(_08975_),
    .A2(_08980_),
    .B1(_08982_),
    .Y(_08983_));
 sky130_fd_sc_hd__nand2_2 _19290_ (.A(_08978_),
    .B(_08983_),
    .Y(_08984_));
 sky130_fd_sc_hd__nand2_1 _19291_ (.A(_08836_),
    .B(_08837_),
    .Y(_08985_));
 sky130_fd_sc_hd__nand2_1 _19292_ (.A(_08985_),
    .B(_06159_),
    .Y(_08986_));
 sky130_fd_sc_hd__nand2_1 _19293_ (.A(_08986_),
    .B(_08838_),
    .Y(_08987_));
 sky130_fd_sc_hd__nand2_1 _19294_ (.A(_08844_),
    .B(_08842_),
    .Y(_08989_));
 sky130_fd_sc_hd__nor2_1 _19295_ (.A(_08987_),
    .B(_08989_),
    .Y(_08990_));
 sky130_fd_sc_hd__nand3_1 _19296_ (.A(_08984_),
    .B(_08826_),
    .C(_08990_),
    .Y(_08991_));
 sky130_fd_sc_hd__nand2_2 _19297_ (.A(_08849_),
    .B(_08991_),
    .Y(_08992_));
 sky130_fd_sc_hd__nand2_1 _19298_ (.A(_08519_),
    .B(_08520_),
    .Y(_08993_));
 sky130_fd_sc_hd__inv_4 _19299_ (.A(_08993_),
    .Y(_08994_));
 sky130_fd_sc_hd__or2_1 _19300_ (.A(_08994_),
    .B(_08432_),
    .X(_08995_));
 sky130_fd_sc_hd__nand2_1 _19301_ (.A(_08432_),
    .B(_08994_),
    .Y(_08996_));
 sky130_fd_sc_hd__nand2_1 _19302_ (.A(_08995_),
    .B(_08996_),
    .Y(_08997_));
 sky130_fd_sc_hd__inv_2 _19303_ (.A(_08997_),
    .Y(_08998_));
 sky130_fd_sc_hd__nand2_1 _19304_ (.A(_08998_),
    .B(_06207_),
    .Y(_09000_));
 sky130_fd_sc_hd__nand2_1 _19305_ (.A(_08997_),
    .B(_08465_),
    .Y(_09001_));
 sky130_fd_sc_hd__nand2_1 _19306_ (.A(_09000_),
    .B(_09001_),
    .Y(_09002_));
 sky130_fd_sc_hd__inv_2 _19307_ (.A(_09002_),
    .Y(_09003_));
 sky130_fd_sc_hd__nand2_1 _19308_ (.A(_08795_),
    .B(_08403_),
    .Y(_09004_));
 sky130_fd_sc_hd__inv_2 _19309_ (.A(_08392_),
    .Y(_09005_));
 sky130_fd_sc_hd__nand2_1 _19310_ (.A(_09004_),
    .B(_09005_),
    .Y(_09006_));
 sky130_fd_sc_hd__nand3_1 _19311_ (.A(_08795_),
    .B(_08392_),
    .C(_08403_),
    .Y(_09007_));
 sky130_fd_sc_hd__nand2_1 _19312_ (.A(_09006_),
    .B(_09007_),
    .Y(_09008_));
 sky130_fd_sc_hd__nand2_1 _19313_ (.A(_09008_),
    .B(_07905_),
    .Y(_09009_));
 sky130_fd_sc_hd__nand3_1 _19314_ (.A(_09006_),
    .B(_06772_),
    .C(_09007_),
    .Y(_09011_));
 sky130_fd_sc_hd__nand3_1 _19315_ (.A(_08803_),
    .B(_09009_),
    .C(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__inv_2 _19316_ (.A(_09012_),
    .Y(_09013_));
 sky130_fd_sc_hd__nand3_1 _19317_ (.A(_08763_),
    .B(_08785_),
    .C(_09013_),
    .Y(_09014_));
 sky130_fd_sc_hd__inv_2 _19318_ (.A(_09009_),
    .Y(_09015_));
 sky130_fd_sc_hd__o21ai_1 _19319_ (.A1(_08799_),
    .A2(_09015_),
    .B1(_09011_),
    .Y(_09016_));
 sky130_fd_sc_hd__nor2_1 _19320_ (.A(_08788_),
    .B(_09012_),
    .Y(_09017_));
 sky130_fd_sc_hd__nor2_1 _19321_ (.A(_09016_),
    .B(_09017_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand2_2 _19322_ (.A(_09014_),
    .B(_09018_),
    .Y(_09019_));
 sky130_fd_sc_hd__or2_1 _19323_ (.A(_09003_),
    .B(_09019_),
    .X(_09020_));
 sky130_fd_sc_hd__buf_6 _19324_ (.A(_08805_),
    .X(_09022_));
 sky130_fd_sc_hd__nand2_1 _19325_ (.A(_09019_),
    .B(_09003_),
    .Y(_09023_));
 sky130_fd_sc_hd__nand3_1 _19326_ (.A(_09020_),
    .B(_09022_),
    .C(_09023_),
    .Y(_09024_));
 sky130_fd_sc_hd__nand2_1 _19327_ (.A(\div1i.quot[14] ),
    .B(_08998_),
    .Y(_09025_));
 sky130_fd_sc_hd__nand2_1 _19328_ (.A(_09024_),
    .B(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__xor2_2 _19329_ (.A(_06754_),
    .B(_09026_),
    .X(_09027_));
 sky130_fd_sc_hd__nand2_1 _19330_ (.A(_09009_),
    .B(_09011_),
    .Y(_09028_));
 sky130_fd_sc_hd__nand2_1 _19331_ (.A(_08804_),
    .B(_08799_),
    .Y(_09029_));
 sky130_fd_sc_hd__xor2_1 _19332_ (.A(_09028_),
    .B(_09029_),
    .X(_09030_));
 sky130_fd_sc_hd__nand2_1 _19333_ (.A(_09030_),
    .B(_09022_),
    .Y(_09031_));
 sky130_fd_sc_hd__nand2_1 _19334_ (.A(\div1i.quot[14] ),
    .B(_09008_),
    .Y(_09033_));
 sky130_fd_sc_hd__nand2_1 _19335_ (.A(_09031_),
    .B(_09033_),
    .Y(_09034_));
 sky130_fd_sc_hd__nand2_1 _19336_ (.A(_09034_),
    .B(_06797_),
    .Y(_09035_));
 sky130_fd_sc_hd__nand3_1 _19337_ (.A(_09031_),
    .B(_06799_),
    .C(_09033_),
    .Y(_09036_));
 sky130_fd_sc_hd__nand2_1 _19338_ (.A(_09035_),
    .B(_09036_),
    .Y(_09037_));
 sky130_fd_sc_hd__nor2_1 _19339_ (.A(_09027_),
    .B(_09037_),
    .Y(_09038_));
 sky130_fd_sc_hd__nand2_2 _19340_ (.A(_08992_),
    .B(_09038_),
    .Y(_09039_));
 sky130_fd_sc_hd__nand2_1 _19341_ (.A(_09026_),
    .B(_06805_),
    .Y(_09040_));
 sky130_fd_sc_hd__o21a_1 _19342_ (.A1(_09036_),
    .A2(_09027_),
    .B1(_09040_),
    .X(_09041_));
 sky130_fd_sc_hd__nand2_1 _19343_ (.A(_09039_),
    .B(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__nand2_1 _19344_ (.A(_08432_),
    .B(_08522_),
    .Y(_09044_));
 sky130_fd_sc_hd__inv_2 _19345_ (.A(_08525_),
    .Y(_09045_));
 sky130_fd_sc_hd__a21o_1 _19346_ (.A1(_09044_),
    .A2(_09045_),
    .B1(_08503_),
    .X(_09046_));
 sky130_fd_sc_hd__nand3_1 _19347_ (.A(_09044_),
    .B(_08503_),
    .C(_09045_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_1 _19348_ (.A(_09046_),
    .B(_09047_),
    .Y(_09048_));
 sky130_fd_sc_hd__inv_2 _19349_ (.A(_09048_),
    .Y(_09049_));
 sky130_fd_sc_hd__nand2_1 _19350_ (.A(_09049_),
    .B(_06819_),
    .Y(_09050_));
 sky130_fd_sc_hd__nand2_1 _19351_ (.A(_09048_),
    .B(_07948_),
    .Y(_09051_));
 sky130_fd_sc_hd__nand2_1 _19352_ (.A(_09050_),
    .B(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__inv_4 _19353_ (.A(_09052_),
    .Y(_09053_));
 sky130_fd_sc_hd__nand2_1 _19354_ (.A(_08996_),
    .B(_08520_),
    .Y(_09055_));
 sky130_fd_sc_hd__xor2_2 _19355_ (.A(_08512_),
    .B(_09055_),
    .X(_09056_));
 sky130_fd_sc_hd__inv_2 _19356_ (.A(_09056_),
    .Y(_09057_));
 sky130_fd_sc_hd__nand2_1 _19357_ (.A(_09057_),
    .B(_06827_),
    .Y(_09058_));
 sky130_fd_sc_hd__nand2_1 _19358_ (.A(_09056_),
    .B(_07957_),
    .Y(_09059_));
 sky130_fd_sc_hd__nand2_1 _19359_ (.A(_09058_),
    .B(_09059_),
    .Y(_09060_));
 sky130_fd_sc_hd__or2_1 _19360_ (.A(_09002_),
    .B(_09060_),
    .X(_09061_));
 sky130_fd_sc_hd__inv_4 _19361_ (.A(_09061_),
    .Y(_09062_));
 sky130_fd_sc_hd__nand2_1 _19362_ (.A(_09019_),
    .B(_09062_),
    .Y(_09063_));
 sky130_fd_sc_hd__inv_2 _19363_ (.A(_09000_),
    .Y(_09064_));
 sky130_fd_sc_hd__a21boi_1 _19364_ (.A1(_09064_),
    .A2(_09059_),
    .B1_N(_09058_),
    .Y(_09066_));
 sky130_fd_sc_hd__nand2_1 _19365_ (.A(_09063_),
    .B(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__or2_1 _19366_ (.A(_09053_),
    .B(_09067_),
    .X(_09068_));
 sky130_fd_sc_hd__nand2_1 _19367_ (.A(_09067_),
    .B(_09053_),
    .Y(_09069_));
 sky130_fd_sc_hd__nand3_1 _19368_ (.A(_09068_),
    .B(_09022_),
    .C(_09069_),
    .Y(_09070_));
 sky130_fd_sc_hd__nand2_1 _19369_ (.A(\div1i.quot[14] ),
    .B(_09049_),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_1 _19370_ (.A(_09070_),
    .B(_09071_),
    .Y(_09072_));
 sky130_fd_sc_hd__xor2_2 _19371_ (.A(_06809_),
    .B(_09072_),
    .X(_09073_));
 sky130_fd_sc_hd__nand2_1 _19372_ (.A(_09023_),
    .B(_09000_),
    .Y(_09074_));
 sky130_fd_sc_hd__xor2_1 _19373_ (.A(_09060_),
    .B(_09074_),
    .X(_09075_));
 sky130_fd_sc_hd__nand2_1 _19374_ (.A(_09075_),
    .B(_09022_),
    .Y(_09077_));
 sky130_fd_sc_hd__nand2_1 _19375_ (.A(\div1i.quot[14] ),
    .B(_09056_),
    .Y(_09078_));
 sky130_fd_sc_hd__nand2_1 _19376_ (.A(_09077_),
    .B(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__or2_1 _19377_ (.A(_06844_),
    .B(_09079_),
    .X(_09080_));
 sky130_fd_sc_hd__nand2_1 _19378_ (.A(_09079_),
    .B(_06844_),
    .Y(_09081_));
 sky130_fd_sc_hd__nand2_1 _19379_ (.A(_09080_),
    .B(_09081_),
    .Y(_09082_));
 sky130_fd_sc_hd__nor2_1 _19380_ (.A(_09073_),
    .B(_09082_),
    .Y(_09083_));
 sky130_fd_sc_hd__nand2_1 _19381_ (.A(_09042_),
    .B(_09083_),
    .Y(_09084_));
 sky130_fd_sc_hd__nand2_1 _19382_ (.A(_09072_),
    .B(_06856_),
    .Y(_09085_));
 sky130_fd_sc_hd__o21a_1 _19383_ (.A1(_09080_),
    .A2(_09073_),
    .B1(_09085_),
    .X(_09086_));
 sky130_fd_sc_hd__nand2_2 _19384_ (.A(_09084_),
    .B(_09086_),
    .Y(_09088_));
 sky130_fd_sc_hd__nand2_1 _19385_ (.A(_08575_),
    .B(_08576_),
    .Y(_09089_));
 sky130_fd_sc_hd__nand2b_1 _19386_ (.A_N(_08529_),
    .B(_09089_),
    .Y(_09090_));
 sky130_fd_sc_hd__nand2b_1 _19387_ (.A_N(_09089_),
    .B(_08529_),
    .Y(_09091_));
 sky130_fd_sc_hd__nand2_1 _19388_ (.A(_09090_),
    .B(_09091_),
    .Y(_09092_));
 sky130_fd_sc_hd__or2_1 _19389_ (.A(_07450_),
    .B(_09092_),
    .X(_09093_));
 sky130_fd_sc_hd__nand2_1 _19390_ (.A(_09092_),
    .B(_07450_),
    .Y(_09094_));
 sky130_fd_sc_hd__nand2_1 _19391_ (.A(_09093_),
    .B(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__inv_4 _19392_ (.A(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__nand2_1 _19393_ (.A(_09046_),
    .B(_08502_),
    .Y(_09097_));
 sky130_fd_sc_hd__inv_2 _19394_ (.A(_08493_),
    .Y(_09099_));
 sky130_fd_sc_hd__nand2_1 _19395_ (.A(_09097_),
    .B(_09099_),
    .Y(_09100_));
 sky130_fd_sc_hd__nand3_1 _19396_ (.A(_09046_),
    .B(_08493_),
    .C(_08502_),
    .Y(_09101_));
 sky130_fd_sc_hd__nand2_1 _19397_ (.A(_09100_),
    .B(_09101_),
    .Y(_09102_));
 sky130_fd_sc_hd__nand2_1 _19398_ (.A(_09102_),
    .B(_08001_),
    .Y(_09103_));
 sky130_fd_sc_hd__nand3_2 _19399_ (.A(_09100_),
    .B(_06874_),
    .C(_09101_),
    .Y(_09104_));
 sky130_fd_sc_hd__nand3_1 _19400_ (.A(_09053_),
    .B(_09103_),
    .C(_09104_),
    .Y(_09105_));
 sky130_fd_sc_hd__inv_2 _19401_ (.A(_09105_),
    .Y(_09106_));
 sky130_fd_sc_hd__nand3_1 _19402_ (.A(_09019_),
    .B(_09062_),
    .C(_09106_),
    .Y(_09107_));
 sky130_fd_sc_hd__inv_2 _19403_ (.A(_09050_),
    .Y(_09108_));
 sky130_fd_sc_hd__inv_2 _19404_ (.A(_09104_),
    .Y(_09110_));
 sky130_fd_sc_hd__a21o_1 _19405_ (.A1(_09103_),
    .A2(_09108_),
    .B1(_09110_),
    .X(_09111_));
 sky130_fd_sc_hd__nor2_1 _19406_ (.A(_09066_),
    .B(_09105_),
    .Y(_09112_));
 sky130_fd_sc_hd__nor2_1 _19407_ (.A(_09111_),
    .B(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__nand2_2 _19408_ (.A(_09107_),
    .B(_09113_),
    .Y(_09114_));
 sky130_fd_sc_hd__or2_1 _19409_ (.A(_09096_),
    .B(_09114_),
    .X(_09115_));
 sky130_fd_sc_hd__nand2_1 _19410_ (.A(_09114_),
    .B(_09096_),
    .Y(_09116_));
 sky130_fd_sc_hd__nand2_1 _19411_ (.A(_09115_),
    .B(_09116_),
    .Y(_09117_));
 sky130_fd_sc_hd__nand2_1 _19412_ (.A(_09117_),
    .B(_09022_),
    .Y(_09118_));
 sky130_fd_sc_hd__nand2_1 _19413_ (.A(\div1i.quot[14] ),
    .B(_09092_),
    .Y(_09119_));
 sky130_fd_sc_hd__nand2_1 _19414_ (.A(_09118_),
    .B(_09119_),
    .Y(_09121_));
 sky130_fd_sc_hd__nand2_1 _19415_ (.A(_09121_),
    .B(_08020_),
    .Y(_09122_));
 sky130_fd_sc_hd__nand3_1 _19416_ (.A(_09118_),
    .B(_06348_),
    .C(_09119_),
    .Y(_09123_));
 sky130_fd_sc_hd__nand2_2 _19417_ (.A(_09122_),
    .B(_09123_),
    .Y(_09124_));
 sky130_fd_sc_hd__inv_2 _19418_ (.A(_09124_),
    .Y(_09125_));
 sky130_fd_sc_hd__nand2_1 _19419_ (.A(_09103_),
    .B(_09104_),
    .Y(_09126_));
 sky130_fd_sc_hd__nand2_1 _19420_ (.A(_09069_),
    .B(_09050_),
    .Y(_09127_));
 sky130_fd_sc_hd__xor2_1 _19421_ (.A(_09126_),
    .B(_09127_),
    .X(_09128_));
 sky130_fd_sc_hd__nand2_1 _19422_ (.A(_09128_),
    .B(_09022_),
    .Y(_09129_));
 sky130_fd_sc_hd__nand2_1 _19423_ (.A(_09102_),
    .B(\div1i.quot[14] ),
    .Y(_09130_));
 sky130_fd_sc_hd__nand2_1 _19424_ (.A(_09129_),
    .B(_09130_),
    .Y(_09132_));
 sky130_fd_sc_hd__nand2_1 _19425_ (.A(_09132_),
    .B(_06903_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand3_2 _19426_ (.A(_09129_),
    .B(_06898_),
    .C(_09130_),
    .Y(_09134_));
 sky130_fd_sc_hd__nand3_1 _19427_ (.A(_09125_),
    .B(_09133_),
    .C(_09134_),
    .Y(_09135_));
 sky130_fd_sc_hd__nand2_1 _19428_ (.A(_09116_),
    .B(_09093_),
    .Y(_09136_));
 sky130_fd_sc_hd__nand2_1 _19429_ (.A(_09091_),
    .B(_08576_),
    .Y(_09137_));
 sky130_fd_sc_hd__or2_1 _19430_ (.A(_08567_),
    .B(_09137_),
    .X(_09138_));
 sky130_fd_sc_hd__nand2_1 _19431_ (.A(_09137_),
    .B(_08567_),
    .Y(_09139_));
 sky130_fd_sc_hd__nand2_1 _19432_ (.A(_09138_),
    .B(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__nand2_1 _19433_ (.A(_09140_),
    .B(_08041_),
    .Y(_09141_));
 sky130_fd_sc_hd__nand3_1 _19434_ (.A(_09138_),
    .B(_07461_),
    .C(_09139_),
    .Y(_09143_));
 sky130_fd_sc_hd__nand2_1 _19435_ (.A(_09141_),
    .B(_09143_),
    .Y(_09144_));
 sky130_fd_sc_hd__inv_2 _19436_ (.A(_09144_),
    .Y(_09145_));
 sky130_fd_sc_hd__nand2_1 _19437_ (.A(_09136_),
    .B(_09145_),
    .Y(_09146_));
 sky130_fd_sc_hd__nand3_1 _19438_ (.A(_09116_),
    .B(_09144_),
    .C(_09093_),
    .Y(_09147_));
 sky130_fd_sc_hd__nand2_1 _19439_ (.A(_09146_),
    .B(_09147_),
    .Y(_09148_));
 sky130_fd_sc_hd__nand2_1 _19440_ (.A(_09148_),
    .B(_09022_),
    .Y(_09149_));
 sky130_fd_sc_hd__nand2_1 _19441_ (.A(_09140_),
    .B(\div1i.quot[14] ),
    .Y(_09150_));
 sky130_fd_sc_hd__nand2_1 _19442_ (.A(_09149_),
    .B(_09150_),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_1 _19443_ (.A(_09151_),
    .B(_07474_),
    .Y(_09152_));
 sky130_fd_sc_hd__nand3_1 _19444_ (.A(_09149_),
    .B(_06366_),
    .C(_09150_),
    .Y(_09154_));
 sky130_fd_sc_hd__nand2_1 _19445_ (.A(_09152_),
    .B(_09154_),
    .Y(_09155_));
 sky130_fd_sc_hd__inv_2 _19446_ (.A(_09155_),
    .Y(_09156_));
 sky130_fd_sc_hd__nand2_1 _19447_ (.A(_09145_),
    .B(_09096_),
    .Y(_09157_));
 sky130_fd_sc_hd__inv_2 _19448_ (.A(_09157_),
    .Y(_09158_));
 sky130_fd_sc_hd__nand2_1 _19449_ (.A(_09114_),
    .B(_09158_),
    .Y(_09159_));
 sky130_fd_sc_hd__o21a_1 _19450_ (.A1(_09093_),
    .A2(_09144_),
    .B1(_09143_),
    .X(_09160_));
 sky130_fd_sc_hd__nand2_1 _19451_ (.A(_09159_),
    .B(_09160_),
    .Y(_09161_));
 sky130_fd_sc_hd__a41o_1 _19452_ (.A1(_08529_),
    .A2(_08567_),
    .A3(_08576_),
    .A4(_08575_),
    .B1(_08629_),
    .X(_09162_));
 sky130_fd_sc_hd__or2_1 _19453_ (.A(_08597_),
    .B(_09162_),
    .X(_09163_));
 sky130_fd_sc_hd__nand2_1 _19454_ (.A(_09162_),
    .B(_08597_),
    .Y(_09165_));
 sky130_fd_sc_hd__nand2_1 _19455_ (.A(_09163_),
    .B(_09165_),
    .Y(_09166_));
 sky130_fd_sc_hd__inv_2 _19456_ (.A(_09166_),
    .Y(_09167_));
 sky130_fd_sc_hd__nand2_1 _19457_ (.A(_09167_),
    .B(_06936_),
    .Y(_09168_));
 sky130_fd_sc_hd__nand2_1 _19458_ (.A(_09166_),
    .B(_08611_),
    .Y(_09169_));
 sky130_fd_sc_hd__nand2_1 _19459_ (.A(_09168_),
    .B(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__inv_2 _19460_ (.A(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__nand2_1 _19461_ (.A(_09161_),
    .B(_09171_),
    .Y(_09172_));
 sky130_fd_sc_hd__nand3_1 _19462_ (.A(_09159_),
    .B(_09170_),
    .C(_09160_),
    .Y(_09173_));
 sky130_fd_sc_hd__nand3_2 _19463_ (.A(_09172_),
    .B(_09173_),
    .C(_09022_),
    .Y(_09174_));
 sky130_fd_sc_hd__nand2_1 _19464_ (.A(_09167_),
    .B(\div1i.quot[14] ),
    .Y(_09176_));
 sky130_fd_sc_hd__nand2_1 _19465_ (.A(_09174_),
    .B(_09176_),
    .Y(_09177_));
 sky130_fd_sc_hd__nand2_1 _19466_ (.A(_09177_),
    .B(_06947_),
    .Y(_09178_));
 sky130_fd_sc_hd__nand3_2 _19467_ (.A(_09174_),
    .B(_06949_),
    .C(_09176_),
    .Y(_09179_));
 sky130_fd_sc_hd__nand2_4 _19468_ (.A(_09178_),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__inv_2 _19469_ (.A(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__nand2_1 _19470_ (.A(_09156_),
    .B(_09181_),
    .Y(_09182_));
 sky130_fd_sc_hd__nor2_1 _19471_ (.A(_09135_),
    .B(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand2_4 _19472_ (.A(_09088_),
    .B(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__o21ai_1 _19473_ (.A1(_09134_),
    .A2(_09124_),
    .B1(_09123_),
    .Y(_09185_));
 sky130_fd_sc_hd__nor2_1 _19474_ (.A(_09180_),
    .B(_09155_),
    .Y(_09187_));
 sky130_fd_sc_hd__o21ai_1 _19475_ (.A1(_09154_),
    .A2(_09180_),
    .B1(_09178_),
    .Y(_09188_));
 sky130_fd_sc_hd__a21oi_2 _19476_ (.A1(_09185_),
    .A2(_09187_),
    .B1(_09188_),
    .Y(_09189_));
 sky130_fd_sc_hd__nand2_2 _19477_ (.A(_09184_),
    .B(_09189_),
    .Y(_09190_));
 sky130_fd_sc_hd__nand2_1 _19478_ (.A(_09165_),
    .B(_08595_),
    .Y(_09191_));
 sky130_fd_sc_hd__xor2_1 _19479_ (.A(_08623_),
    .B(_09191_),
    .X(_09192_));
 sky130_fd_sc_hd__nand3_1 _19480_ (.A(_09172_),
    .B(_09022_),
    .C(_09168_),
    .Y(_09193_));
 sky130_fd_sc_hd__xnor2_2 _19481_ (.A(_09192_),
    .B(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__nand2_8 _19482_ (.A(_09190_),
    .B(_09194_),
    .Y(_09195_));
 sky130_fd_sc_hd__inv_2 _19483_ (.A(_09194_),
    .Y(_09196_));
 sky130_fd_sc_hd__nand3_4 _19484_ (.A(_09184_),
    .B(_09189_),
    .C(_09196_),
    .Y(_09198_));
 sky130_fd_sc_hd__nand2_8 _19485_ (.A(_09195_),
    .B(_09198_),
    .Y(_09199_));
 sky130_fd_sc_hd__buf_12 _19486_ (.A(_09199_),
    .X(_09200_));
 sky130_fd_sc_hd__buf_8 _19487_ (.A(net238),
    .X(\div1i.quot[13] ));
 sky130_fd_sc_hd__nand2_1 _19488_ (.A(_08866_),
    .B(_08870_),
    .Y(_09201_));
 sky130_fd_sc_hd__nand2_1 _19489_ (.A(_09201_),
    .B(_08871_),
    .Y(_09202_));
 sky130_fd_sc_hd__nand2_1 _19490_ (.A(_09202_),
    .B(_08873_),
    .Y(_09203_));
 sky130_fd_sc_hd__inv_2 _19491_ (.A(_09203_),
    .Y(_09204_));
 sky130_fd_sc_hd__nand2_1 _19492_ (.A(_09200_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__o21ai_1 _19493_ (.A1(_06979_),
    .A2(\div1i.quot[14] ),
    .B1(_06980_),
    .Y(_09206_));
 sky130_fd_sc_hd__nand2_1 _19494_ (.A(_09203_),
    .B(_06982_),
    .Y(_09208_));
 sky130_fd_sc_hd__nand3_1 _19495_ (.A(_09202_),
    .B(_06984_),
    .C(_08873_),
    .Y(_09209_));
 sky130_fd_sc_hd__nand2_1 _19496_ (.A(_09208_),
    .B(_09209_),
    .Y(_09210_));
 sky130_fd_sc_hd__xor2_1 _19497_ (.A(_09206_),
    .B(_09210_),
    .X(_09211_));
 sky130_fd_sc_hd__nand3b_1 _19498_ (.A_N(_09211_),
    .B(_09195_),
    .C(_09198_),
    .Y(_09212_));
 sky130_fd_sc_hd__nand2_1 _19499_ (.A(_09205_),
    .B(_09212_),
    .Y(_09213_));
 sky130_fd_sc_hd__nand2_1 _19500_ (.A(_09213_),
    .B(_08857_),
    .Y(_09214_));
 sky130_fd_sc_hd__buf_6 _19501_ (.A(_06979_),
    .X(_09215_));
 sky130_fd_sc_hd__nor2_1 _19502_ (.A(_09215_),
    .B(_09022_),
    .Y(_09216_));
 sky130_fd_sc_hd__or2_1 _19503_ (.A(_06607_),
    .B(_09216_),
    .X(_09217_));
 sky130_fd_sc_hd__nand2_1 _19504_ (.A(_09217_),
    .B(_08871_),
    .Y(_09219_));
 sky130_fd_sc_hd__inv_2 _19505_ (.A(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__nand2_1 _19506_ (.A(_09200_),
    .B(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__nand3_1 _19507_ (.A(_09195_),
    .B(_09198_),
    .C(_09216_),
    .Y(_09222_));
 sky130_fd_sc_hd__nand2_1 _19508_ (.A(_09221_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__nand2_2 _19509_ (.A(_09223_),
    .B(_06615_),
    .Y(_09224_));
 sky130_fd_sc_hd__nand2_1 _19510_ (.A(_09214_),
    .B(_09224_),
    .Y(_09225_));
 sky130_fd_sc_hd__inv_2 _19511_ (.A(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__nand3_1 _19512_ (.A(_09221_),
    .B(_06620_),
    .C(_09222_),
    .Y(_09227_));
 sky130_fd_sc_hd__buf_6 _19513_ (.A(_06980_),
    .X(_09228_));
 sky130_fd_sc_hd__nand3_2 _19514_ (.A(_09200_),
    .B(_09228_),
    .C(_07004_),
    .Y(_09230_));
 sky130_fd_sc_hd__inv_2 _19515_ (.A(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__nand3_4 _19516_ (.A(_09224_),
    .B(_09227_),
    .C(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__or2_4 _19517_ (.A(_08857_),
    .B(_09213_),
    .X(_09233_));
 sky130_fd_sc_hd__inv_2 _19518_ (.A(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__a21oi_2 _19519_ (.A1(_09226_),
    .A2(_09232_),
    .B1(_09234_),
    .Y(_09235_));
 sky130_fd_sc_hd__nand2_1 _19520_ (.A(_08869_),
    .B(_08873_),
    .Y(_09236_));
 sky130_fd_sc_hd__nand2_1 _19521_ (.A(_09236_),
    .B(_08874_),
    .Y(_09237_));
 sky130_fd_sc_hd__inv_2 _19522_ (.A(_08927_),
    .Y(_09238_));
 sky130_fd_sc_hd__o21ai_1 _19523_ (.A1(_08923_),
    .A2(_09237_),
    .B1(_09238_),
    .Y(_09239_));
 sky130_fd_sc_hd__or2_1 _19524_ (.A(_08898_),
    .B(_09239_),
    .X(_09241_));
 sky130_fd_sc_hd__nand2_1 _19525_ (.A(_09239_),
    .B(_08898_),
    .Y(_09242_));
 sky130_fd_sc_hd__nand2_1 _19526_ (.A(_09241_),
    .B(_09242_),
    .Y(_09243_));
 sky130_fd_sc_hd__inv_2 _19527_ (.A(_09243_),
    .Y(_09244_));
 sky130_fd_sc_hd__nand2_1 _19528_ (.A(_09199_),
    .B(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__nand2_1 _19529_ (.A(_09244_),
    .B(_07021_),
    .Y(_09246_));
 sky130_fd_sc_hd__nand2_1 _19530_ (.A(_09243_),
    .B(_07024_),
    .Y(_09247_));
 sky130_fd_sc_hd__nand2_1 _19531_ (.A(_09246_),
    .B(_09247_),
    .Y(_09248_));
 sky130_fd_sc_hd__inv_2 _19532_ (.A(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__nand2_1 _19533_ (.A(_08875_),
    .B(_08921_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand2_1 _19534_ (.A(_09237_),
    .B(_08920_),
    .Y(_09252_));
 sky130_fd_sc_hd__nand2_1 _19535_ (.A(_09250_),
    .B(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__nand2_1 _19536_ (.A(_09253_),
    .B(_07031_),
    .Y(_09254_));
 sky130_fd_sc_hd__nand3_1 _19537_ (.A(_09250_),
    .B(_07034_),
    .C(_09252_),
    .Y(_09255_));
 sky130_fd_sc_hd__nand2_1 _19538_ (.A(_09254_),
    .B(_09255_),
    .Y(_09256_));
 sky130_fd_sc_hd__inv_2 _19539_ (.A(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__inv_2 _19540_ (.A(_09209_),
    .Y(_09258_));
 sky130_fd_sc_hd__a21o_1 _19541_ (.A1(_09208_),
    .A2(_09206_),
    .B1(_09258_),
    .X(_09259_));
 sky130_fd_sc_hd__nand2_1 _19542_ (.A(_08874_),
    .B(_08858_),
    .Y(_09260_));
 sky130_fd_sc_hd__nand2_1 _19543_ (.A(_08873_),
    .B(_08866_),
    .Y(_09261_));
 sky130_fd_sc_hd__xor2_2 _19544_ (.A(_09260_),
    .B(_09261_),
    .X(_09263_));
 sky130_fd_sc_hd__nand2_1 _19545_ (.A(_09263_),
    .B(_07043_),
    .Y(_09264_));
 sky130_fd_sc_hd__nand2_1 _19546_ (.A(_09259_),
    .B(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__inv_2 _19547_ (.A(_09263_),
    .Y(_09266_));
 sky130_fd_sc_hd__nand2_1 _19548_ (.A(_09266_),
    .B(_07048_),
    .Y(_09267_));
 sky130_fd_sc_hd__nand2_1 _19549_ (.A(_09265_),
    .B(_09267_),
    .Y(_09268_));
 sky130_fd_sc_hd__nand2_1 _19550_ (.A(_09257_),
    .B(_09268_),
    .Y(_09269_));
 sky130_fd_sc_hd__nand2_1 _19551_ (.A(_09269_),
    .B(_09255_),
    .Y(_09270_));
 sky130_fd_sc_hd__nand2_1 _19552_ (.A(_09250_),
    .B(_08918_),
    .Y(_09271_));
 sky130_fd_sc_hd__xor2_1 _19553_ (.A(_08910_),
    .B(_09271_),
    .X(_09272_));
 sky130_fd_sc_hd__nand2_1 _19554_ (.A(_09272_),
    .B(_06465_),
    .Y(_09274_));
 sky130_fd_sc_hd__nand2_1 _19555_ (.A(_09270_),
    .B(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__inv_2 _19556_ (.A(_09272_),
    .Y(_09276_));
 sky130_fd_sc_hd__nand2_1 _19557_ (.A(_09276_),
    .B(_08176_),
    .Y(_09277_));
 sky130_fd_sc_hd__nand2_1 _19558_ (.A(_09275_),
    .B(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__or2_1 _19559_ (.A(_09249_),
    .B(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__nand2_1 _19560_ (.A(_09278_),
    .B(_09249_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_1 _19561_ (.A(_09279_),
    .B(_09280_),
    .Y(_09281_));
 sky130_fd_sc_hd__inv_2 _19562_ (.A(_09281_),
    .Y(_09282_));
 sky130_fd_sc_hd__nand3_1 _19563_ (.A(_09195_),
    .B(_09198_),
    .C(_09282_),
    .Y(_09283_));
 sky130_fd_sc_hd__nand2_1 _19564_ (.A(_09245_),
    .B(_09283_),
    .Y(_09285_));
 sky130_fd_sc_hd__nand2_1 _19565_ (.A(_09285_),
    .B(_06636_),
    .Y(_09286_));
 sky130_fd_sc_hd__nand3_1 _19566_ (.A(_09245_),
    .B(_06639_),
    .C(_09283_),
    .Y(_09287_));
 sky130_fd_sc_hd__nand2_1 _19567_ (.A(_09286_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__inv_2 _19568_ (.A(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nand2_1 _19569_ (.A(_09199_),
    .B(_09276_),
    .Y(_09290_));
 sky130_fd_sc_hd__nand2_1 _19570_ (.A(_09277_),
    .B(_09274_),
    .Y(_09291_));
 sky130_fd_sc_hd__xnor2_1 _19571_ (.A(_09270_),
    .B(_09291_),
    .Y(_09292_));
 sky130_fd_sc_hd__nand3_1 _19572_ (.A(_09195_),
    .B(_09198_),
    .C(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__nand2_1 _19573_ (.A(_09290_),
    .B(_09293_),
    .Y(_09294_));
 sky130_fd_sc_hd__nand2_2 _19574_ (.A(_09294_),
    .B(_06651_),
    .Y(_09296_));
 sky130_fd_sc_hd__nand3_1 _19575_ (.A(_09290_),
    .B(_06648_),
    .C(_09293_),
    .Y(_09297_));
 sky130_fd_sc_hd__nand2_1 _19576_ (.A(_09296_),
    .B(_09297_),
    .Y(_09298_));
 sky130_fd_sc_hd__inv_2 _19577_ (.A(_09298_),
    .Y(_09299_));
 sky130_fd_sc_hd__nand2_1 _19578_ (.A(_09289_),
    .B(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__inv_2 _19579_ (.A(_09253_),
    .Y(_09301_));
 sky130_fd_sc_hd__nand2_1 _19580_ (.A(_09199_),
    .B(_09301_),
    .Y(_09302_));
 sky130_fd_sc_hd__or2_1 _19581_ (.A(_09268_),
    .B(_09257_),
    .X(_09303_));
 sky130_fd_sc_hd__nand2_1 _19582_ (.A(_09303_),
    .B(_09269_),
    .Y(_09304_));
 sky130_fd_sc_hd__clkinvlp_2 _19583_ (.A(_09304_),
    .Y(_09305_));
 sky130_fd_sc_hd__nand3_1 _19584_ (.A(_09195_),
    .B(_09198_),
    .C(_09305_),
    .Y(_09307_));
 sky130_fd_sc_hd__nand2_1 _19585_ (.A(_09302_),
    .B(_09307_),
    .Y(_09308_));
 sky130_fd_sc_hd__nand2_1 _19586_ (.A(_09308_),
    .B(_06033_),
    .Y(_09309_));
 sky130_fd_sc_hd__nand3_1 _19587_ (.A(_09302_),
    .B(_07092_),
    .C(_09307_),
    .Y(_09310_));
 sky130_fd_sc_hd__nand2_2 _19588_ (.A(_09309_),
    .B(_09310_),
    .Y(_09311_));
 sky130_fd_sc_hd__inv_2 _19589_ (.A(_09311_),
    .Y(_09312_));
 sky130_fd_sc_hd__nand2_1 _19590_ (.A(_09199_),
    .B(_09266_),
    .Y(_09313_));
 sky130_fd_sc_hd__nand2_1 _19591_ (.A(_09267_),
    .B(_09264_),
    .Y(_09314_));
 sky130_fd_sc_hd__xnor2_1 _19592_ (.A(_09259_),
    .B(_09314_),
    .Y(_09315_));
 sky130_fd_sc_hd__nand3_1 _19593_ (.A(_09195_),
    .B(_09198_),
    .C(_09315_),
    .Y(_09316_));
 sky130_fd_sc_hd__nand2_1 _19594_ (.A(_09313_),
    .B(_09316_),
    .Y(_09318_));
 sky130_fd_sc_hd__nand2_1 _19595_ (.A(_09318_),
    .B(_07102_),
    .Y(_09319_));
 sky130_fd_sc_hd__nand3_1 _19596_ (.A(_09313_),
    .B(_06046_),
    .C(_09316_),
    .Y(_09320_));
 sky130_fd_sc_hd__nand2_1 _19597_ (.A(_09319_),
    .B(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__inv_2 _19598_ (.A(_09321_),
    .Y(_09322_));
 sky130_fd_sc_hd__nand2_1 _19599_ (.A(_09312_),
    .B(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__nor2_1 _19600_ (.A(_09300_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__nand2_1 _19601_ (.A(_09235_),
    .B(_09324_),
    .Y(_09325_));
 sky130_fd_sc_hd__inv_2 _19602_ (.A(_09310_),
    .Y(_09326_));
 sky130_fd_sc_hd__o21ai_2 _19603_ (.A1(_09319_),
    .A2(_09326_),
    .B1(_09309_),
    .Y(_09327_));
 sky130_fd_sc_hd__nor2_1 _19604_ (.A(_09288_),
    .B(_09298_),
    .Y(_09329_));
 sky130_fd_sc_hd__inv_2 _19605_ (.A(_09287_),
    .Y(_09330_));
 sky130_fd_sc_hd__o21ai_1 _19606_ (.A1(_09296_),
    .A2(_09330_),
    .B1(_09286_),
    .Y(_09331_));
 sky130_fd_sc_hd__a21oi_1 _19607_ (.A1(_09327_),
    .A2(_09329_),
    .B1(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__nand2_2 _19608_ (.A(_09325_),
    .B(_09332_),
    .Y(_09333_));
 sky130_fd_sc_hd__inv_2 _19609_ (.A(_08956_),
    .Y(_09334_));
 sky130_fd_sc_hd__nand2_1 _19610_ (.A(_08932_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__inv_2 _19611_ (.A(_08980_),
    .Y(_09336_));
 sky130_fd_sc_hd__nand2_1 _19612_ (.A(_09335_),
    .B(_09336_),
    .Y(_09337_));
 sky130_fd_sc_hd__inv_2 _19613_ (.A(_08967_),
    .Y(_09338_));
 sky130_fd_sc_hd__nand2_1 _19614_ (.A(_09337_),
    .B(_09338_),
    .Y(_09340_));
 sky130_fd_sc_hd__nand3_1 _19615_ (.A(_09335_),
    .B(_08967_),
    .C(_09336_),
    .Y(_09341_));
 sky130_fd_sc_hd__nand2_1 _19616_ (.A(_09340_),
    .B(_09341_),
    .Y(_09342_));
 sky130_fd_sc_hd__inv_2 _19617_ (.A(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__nand2_1 _19618_ (.A(_09343_),
    .B(_07128_),
    .Y(_09344_));
 sky130_fd_sc_hd__nand2_1 _19619_ (.A(_09342_),
    .B(_07130_),
    .Y(_09345_));
 sky130_fd_sc_hd__nand2_1 _19620_ (.A(_09344_),
    .B(_09345_),
    .Y(_09346_));
 sky130_fd_sc_hd__inv_2 _19621_ (.A(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__nand2_1 _19622_ (.A(_09242_),
    .B(_08896_),
    .Y(_09348_));
 sky130_fd_sc_hd__or2_1 _19623_ (.A(_08888_),
    .B(_09348_),
    .X(_09349_));
 sky130_fd_sc_hd__nand2_1 _19624_ (.A(_09348_),
    .B(_08888_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand3_1 _19625_ (.A(_09349_),
    .B(_05896_),
    .C(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_1 _19626_ (.A(_09352_),
    .B(_09246_),
    .Y(_09353_));
 sky130_fd_sc_hd__inv_2 _19627_ (.A(_09353_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_1 _19628_ (.A(_09280_),
    .B(_09354_),
    .Y(_09355_));
 sky130_fd_sc_hd__nand2_1 _19629_ (.A(_08932_),
    .B(_08954_),
    .Y(_09356_));
 sky130_fd_sc_hd__nand2_1 _19630_ (.A(_09356_),
    .B(_08952_),
    .Y(_09357_));
 sky130_fd_sc_hd__xor2_1 _19631_ (.A(_08941_),
    .B(_09357_),
    .X(_09358_));
 sky130_fd_sc_hd__nand2_2 _19632_ (.A(_09358_),
    .B(_07146_),
    .Y(_09359_));
 sky130_fd_sc_hd__or2_1 _19633_ (.A(_08942_),
    .B(_09357_),
    .X(_09360_));
 sky130_fd_sc_hd__nand2_1 _19634_ (.A(_09357_),
    .B(_08942_),
    .Y(_09362_));
 sky130_fd_sc_hd__nand3_2 _19635_ (.A(_09360_),
    .B(_07149_),
    .C(_09362_),
    .Y(_09363_));
 sky130_fd_sc_hd__or2_1 _19636_ (.A(_08954_),
    .B(_08932_),
    .X(_09364_));
 sky130_fd_sc_hd__nand2_1 _19637_ (.A(_09364_),
    .B(_09356_),
    .Y(_09365_));
 sky130_fd_sc_hd__nand2_1 _19638_ (.A(_09365_),
    .B(_07155_),
    .Y(_09366_));
 sky130_fd_sc_hd__nand3_2 _19639_ (.A(_09364_),
    .B(_07157_),
    .C(_09356_),
    .Y(_09367_));
 sky130_fd_sc_hd__nand2_1 _19640_ (.A(_09366_),
    .B(_09367_),
    .Y(_09368_));
 sky130_fd_sc_hd__inv_2 _19641_ (.A(_09368_),
    .Y(_09369_));
 sky130_fd_sc_hd__nand3_1 _19642_ (.A(_09359_),
    .B(_09363_),
    .C(_09369_),
    .Y(_09370_));
 sky130_fd_sc_hd__inv_2 _19643_ (.A(_09370_),
    .Y(_09371_));
 sky130_fd_sc_hd__nand2_1 _19644_ (.A(_09349_),
    .B(_09351_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand2_2 _19645_ (.A(_09373_),
    .B(_08738_),
    .Y(_09374_));
 sky130_fd_sc_hd__nand3_2 _19646_ (.A(_09355_),
    .B(_09371_),
    .C(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__inv_2 _19647_ (.A(_09367_),
    .Y(_09376_));
 sky130_fd_sc_hd__a21boi_2 _19648_ (.A1(_09359_),
    .A2(_09376_),
    .B1_N(_09363_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand2_1 _19649_ (.A(_09375_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__or2_1 _19650_ (.A(_09347_),
    .B(_09378_),
    .X(_09379_));
 sky130_fd_sc_hd__inv_6 _19651_ (.A(_09199_),
    .Y(_09380_));
 sky130_fd_sc_hd__nand2_1 _19652_ (.A(_09378_),
    .B(_09347_),
    .Y(_09381_));
 sky130_fd_sc_hd__nand3_1 _19653_ (.A(_09379_),
    .B(_09380_),
    .C(_09381_),
    .Y(_09382_));
 sky130_fd_sc_hd__nand2_1 _19654_ (.A(_09200_),
    .B(_09343_),
    .Y(_09384_));
 sky130_fd_sc_hd__nand2_1 _19655_ (.A(_09382_),
    .B(_09384_),
    .Y(_09385_));
 sky130_fd_sc_hd__nand2_1 _19656_ (.A(_09385_),
    .B(_06731_),
    .Y(_09386_));
 sky130_fd_sc_hd__nand3_1 _19657_ (.A(_09382_),
    .B(_06733_),
    .C(_09384_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand2_1 _19658_ (.A(_09386_),
    .B(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__nand3_1 _19659_ (.A(_09355_),
    .B(_09374_),
    .C(_09369_),
    .Y(_09389_));
 sky130_fd_sc_hd__nand2_1 _19660_ (.A(_09389_),
    .B(_09367_),
    .Y(_09390_));
 sky130_fd_sc_hd__nand3_1 _19661_ (.A(_09390_),
    .B(_09363_),
    .C(_09359_),
    .Y(_09391_));
 sky130_fd_sc_hd__nand2_1 _19662_ (.A(_09359_),
    .B(_09363_),
    .Y(_09392_));
 sky130_fd_sc_hd__nand3_1 _19663_ (.A(_09389_),
    .B(_09392_),
    .C(_09367_),
    .Y(_09393_));
 sky130_fd_sc_hd__a21o_1 _19664_ (.A1(_09391_),
    .A2(_09393_),
    .B1(net238),
    .X(_09395_));
 sky130_fd_sc_hd__nand2_1 _19665_ (.A(net238),
    .B(_09358_),
    .Y(_09396_));
 sky130_fd_sc_hd__nand2_1 _19666_ (.A(_09395_),
    .B(_09396_),
    .Y(_09397_));
 sky130_fd_sc_hd__nand2_1 _19667_ (.A(_09397_),
    .B(_06721_),
    .Y(_09398_));
 sky130_fd_sc_hd__nand3_4 _19668_ (.A(_09395_),
    .B(_06723_),
    .C(_09396_),
    .Y(_09399_));
 sky130_fd_sc_hd__nand2_2 _19669_ (.A(_09398_),
    .B(_09399_),
    .Y(_09400_));
 sky130_fd_sc_hd__nor2_2 _19670_ (.A(_09400_),
    .B(_09388_),
    .Y(_09401_));
 sky130_fd_sc_hd__a21o_1 _19671_ (.A1(_09355_),
    .A2(_09374_),
    .B1(_09369_),
    .X(_09402_));
 sky130_fd_sc_hd__nand3_1 _19672_ (.A(_09380_),
    .B(_09389_),
    .C(_09402_),
    .Y(_09403_));
 sky130_fd_sc_hd__a21o_1 _19673_ (.A1(_09195_),
    .A2(_09198_),
    .B1(_09365_),
    .X(_09404_));
 sky130_fd_sc_hd__nand2_1 _19674_ (.A(_09403_),
    .B(_09404_),
    .Y(_09406_));
 sky130_fd_sc_hd__nand2_1 _19675_ (.A(_09406_),
    .B(_06695_),
    .Y(_09407_));
 sky130_fd_sc_hd__nand3_1 _19676_ (.A(_09403_),
    .B(_06697_),
    .C(_09404_),
    .Y(_09408_));
 sky130_fd_sc_hd__nand2_1 _19677_ (.A(_09407_),
    .B(_09408_),
    .Y(_09409_));
 sky130_fd_sc_hd__buf_6 _19678_ (.A(_05915_),
    .X(_09410_));
 sky130_fd_sc_hd__nand2_1 _19679_ (.A(_09374_),
    .B(_09352_),
    .Y(_09411_));
 sky130_fd_sc_hd__nand2_1 _19680_ (.A(_09280_),
    .B(_09246_),
    .Y(_09412_));
 sky130_fd_sc_hd__xor2_1 _19681_ (.A(_09411_),
    .B(_09412_),
    .X(_09413_));
 sky130_fd_sc_hd__nand2_1 _19682_ (.A(_09380_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__nand2_1 _19683_ (.A(_09200_),
    .B(_09373_),
    .Y(_09415_));
 sky130_fd_sc_hd__nand2_1 _19684_ (.A(_09414_),
    .B(_09415_),
    .Y(_09417_));
 sky130_fd_sc_hd__or2_4 _19685_ (.A(_09410_),
    .B(_09417_),
    .X(_09418_));
 sky130_fd_sc_hd__nand2_1 _19686_ (.A(_09417_),
    .B(_09410_),
    .Y(_09419_));
 sky130_fd_sc_hd__nand2_1 _19687_ (.A(_09418_),
    .B(_09419_),
    .Y(_09420_));
 sky130_fd_sc_hd__nor2_1 _19688_ (.A(_09409_),
    .B(_09420_),
    .Y(_09421_));
 sky130_fd_sc_hd__nand2_1 _19689_ (.A(_09401_),
    .B(_09421_),
    .Y(_09422_));
 sky130_fd_sc_hd__inv_2 _19690_ (.A(_09422_),
    .Y(_09423_));
 sky130_fd_sc_hd__nand2_1 _19691_ (.A(_09333_),
    .B(_09423_),
    .Y(_09424_));
 sky130_fd_sc_hd__o21ai_2 _19692_ (.A1(_09418_),
    .A2(_09409_),
    .B1(_09407_),
    .Y(_09425_));
 sky130_fd_sc_hd__o21ai_1 _19693_ (.A1(_09399_),
    .A2(_09388_),
    .B1(_09386_),
    .Y(_09426_));
 sky130_fd_sc_hd__a21oi_1 _19694_ (.A1(_09425_),
    .A2(_09401_),
    .B1(_09426_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand2_2 _19695_ (.A(_09424_),
    .B(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__inv_2 _19696_ (.A(_09375_),
    .Y(_09430_));
 sky130_fd_sc_hd__nand2_1 _19697_ (.A(_09340_),
    .B(_08965_),
    .Y(_09431_));
 sky130_fd_sc_hd__inv_2 _19698_ (.A(_08974_),
    .Y(_09432_));
 sky130_fd_sc_hd__nand2_1 _19699_ (.A(_09431_),
    .B(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__nand3_1 _19700_ (.A(_09340_),
    .B(_08965_),
    .C(_08974_),
    .Y(_09434_));
 sky130_fd_sc_hd__nand2_1 _19701_ (.A(_09433_),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__nand2_1 _19702_ (.A(_09435_),
    .B(_07226_),
    .Y(_09436_));
 sky130_fd_sc_hd__nand3_1 _19703_ (.A(_09433_),
    .B(_07228_),
    .C(_09434_),
    .Y(_09437_));
 sky130_fd_sc_hd__nand3_1 _19704_ (.A(_09347_),
    .B(_09436_),
    .C(_09437_),
    .Y(_09439_));
 sky130_fd_sc_hd__inv_2 _19705_ (.A(_09439_),
    .Y(_09440_));
 sky130_fd_sc_hd__nand2_1 _19706_ (.A(_09430_),
    .B(_09440_),
    .Y(_09441_));
 sky130_fd_sc_hd__nor2_1 _19707_ (.A(_09377_),
    .B(_09439_),
    .Y(_09442_));
 sky130_fd_sc_hd__nand2_1 _19708_ (.A(_09436_),
    .B(_09437_),
    .Y(_09443_));
 sky130_fd_sc_hd__o21ai_1 _19709_ (.A1(_09344_),
    .A2(_09443_),
    .B1(_09437_),
    .Y(_09444_));
 sky130_fd_sc_hd__nor2_1 _19710_ (.A(_09442_),
    .B(_09444_),
    .Y(_09445_));
 sky130_fd_sc_hd__nand2_2 _19711_ (.A(_09441_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__inv_2 _19712_ (.A(_08989_),
    .Y(_09447_));
 sky130_fd_sc_hd__inv_2 _19713_ (.A(_08987_),
    .Y(_09448_));
 sky130_fd_sc_hd__nand2_1 _19714_ (.A(_08984_),
    .B(_09448_),
    .Y(_09450_));
 sky130_fd_sc_hd__nand2_1 _19715_ (.A(_09450_),
    .B(_08838_),
    .Y(_09451_));
 sky130_fd_sc_hd__or2_1 _19716_ (.A(_09447_),
    .B(_09451_),
    .X(_09452_));
 sky130_fd_sc_hd__nand2_1 _19717_ (.A(_09451_),
    .B(_09447_),
    .Y(_09453_));
 sky130_fd_sc_hd__nand2_1 _19718_ (.A(_09452_),
    .B(_09453_),
    .Y(_09454_));
 sky130_fd_sc_hd__nand2_1 _19719_ (.A(_09454_),
    .B(_07247_),
    .Y(_09455_));
 sky130_fd_sc_hd__nand3_1 _19720_ (.A(_09452_),
    .B(_07249_),
    .C(_09453_),
    .Y(_09456_));
 sky130_fd_sc_hd__nand2_1 _19721_ (.A(_09455_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__inv_2 _19722_ (.A(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__or2_1 _19723_ (.A(_09448_),
    .B(_08984_),
    .X(_09459_));
 sky130_fd_sc_hd__nand2_1 _19724_ (.A(_09459_),
    .B(_09450_),
    .Y(_09461_));
 sky130_fd_sc_hd__inv_2 _19725_ (.A(_09461_),
    .Y(_09462_));
 sky130_fd_sc_hd__nand2_1 _19726_ (.A(_09462_),
    .B(_06521_),
    .Y(_09463_));
 sky130_fd_sc_hd__nand2_1 _19727_ (.A(_09461_),
    .B(_07677_),
    .Y(_09464_));
 sky130_fd_sc_hd__nand2_1 _19728_ (.A(_09463_),
    .B(_09464_),
    .Y(_09465_));
 sky130_fd_sc_hd__inv_4 _19729_ (.A(_09465_),
    .Y(_09466_));
 sky130_fd_sc_hd__nand2_1 _19730_ (.A(_09458_),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__inv_2 _19731_ (.A(_09467_),
    .Y(_09468_));
 sky130_fd_sc_hd__nand2_1 _19732_ (.A(_09446_),
    .B(_09468_),
    .Y(_09469_));
 sky130_fd_sc_hd__inv_2 _19733_ (.A(_09463_),
    .Y(_09470_));
 sky130_fd_sc_hd__a21boi_2 _19734_ (.A1(_09455_),
    .A2(_09470_),
    .B1_N(_09456_),
    .Y(_09472_));
 sky130_fd_sc_hd__nand2_1 _19735_ (.A(_09469_),
    .B(_09472_),
    .Y(_09473_));
 sky130_fd_sc_hd__nand2_1 _19736_ (.A(_08984_),
    .B(_08990_),
    .Y(_09474_));
 sky130_fd_sc_hd__inv_2 _19737_ (.A(_08846_),
    .Y(_09475_));
 sky130_fd_sc_hd__nand2_1 _19738_ (.A(_09474_),
    .B(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__inv_2 _19739_ (.A(_08825_),
    .Y(_09477_));
 sky130_fd_sc_hd__nand2_1 _19740_ (.A(_09476_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__nand3_1 _19741_ (.A(_09474_),
    .B(_09475_),
    .C(_08825_),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2_1 _19742_ (.A(_09478_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__nand2_1 _19743_ (.A(_09480_),
    .B(_07276_),
    .Y(_09481_));
 sky130_fd_sc_hd__nand3_1 _19744_ (.A(_09478_),
    .B(_09479_),
    .C(_07278_),
    .Y(_09483_));
 sky130_fd_sc_hd__nand2_1 _19745_ (.A(_09481_),
    .B(_09483_),
    .Y(_09484_));
 sky130_fd_sc_hd__inv_2 _19746_ (.A(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__nand2_1 _19747_ (.A(_09473_),
    .B(_09485_),
    .Y(_09486_));
 sky130_fd_sc_hd__nand3_1 _19748_ (.A(_09469_),
    .B(_09484_),
    .C(_09472_),
    .Y(_09487_));
 sky130_fd_sc_hd__nand3_1 _19749_ (.A(_09486_),
    .B(_09380_),
    .C(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__or2_1 _19750_ (.A(_09480_),
    .B(_09380_),
    .X(_09489_));
 sky130_fd_sc_hd__nand2_1 _19751_ (.A(_09488_),
    .B(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__nand2_1 _19752_ (.A(_09490_),
    .B(_06554_),
    .Y(_09491_));
 sky130_fd_sc_hd__nand3_1 _19753_ (.A(_09488_),
    .B(_06556_),
    .C(_09489_),
    .Y(_09492_));
 sky130_fd_sc_hd__nand2_1 _19754_ (.A(_09491_),
    .B(_09492_),
    .Y(_09494_));
 sky130_fd_sc_hd__nand2_1 _19755_ (.A(_09446_),
    .B(_09466_),
    .Y(_09495_));
 sky130_fd_sc_hd__nand2_1 _19756_ (.A(_09495_),
    .B(_09463_),
    .Y(_09496_));
 sky130_fd_sc_hd__nand2_1 _19757_ (.A(_09496_),
    .B(_09458_),
    .Y(_09497_));
 sky130_fd_sc_hd__nand3_1 _19758_ (.A(_09495_),
    .B(_09457_),
    .C(_09463_),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_1 _19759_ (.A(_09497_),
    .B(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__nand2_1 _19760_ (.A(_09499_),
    .B(_09380_),
    .Y(_09500_));
 sky130_fd_sc_hd__nand2_1 _19761_ (.A(\div1i.quot[13] ),
    .B(_09454_),
    .Y(_09501_));
 sky130_fd_sc_hd__nand2_1 _19762_ (.A(_09500_),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__nand2_1 _19763_ (.A(_09502_),
    .B(_06568_),
    .Y(_09503_));
 sky130_fd_sc_hd__nand3_2 _19764_ (.A(_09500_),
    .B(_06570_),
    .C(_09501_),
    .Y(_09505_));
 sky130_fd_sc_hd__nand2_1 _19765_ (.A(_09503_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__nor2_2 _19766_ (.A(_09494_),
    .B(_09506_),
    .Y(_09507_));
 sky130_fd_sc_hd__or2_1 _19767_ (.A(_09466_),
    .B(_09446_),
    .X(_09508_));
 sky130_fd_sc_hd__nand3_1 _19768_ (.A(_09508_),
    .B(_09380_),
    .C(_09495_),
    .Y(_09509_));
 sky130_fd_sc_hd__nand2_1 _19769_ (.A(net238),
    .B(_09462_),
    .Y(_09510_));
 sky130_fd_sc_hd__nand2_1 _19770_ (.A(_09509_),
    .B(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__nand2_1 _19771_ (.A(_09511_),
    .B(_06149_),
    .Y(_09512_));
 sky130_fd_sc_hd__nand3_1 _19772_ (.A(_09509_),
    .B(_06592_),
    .C(_09510_),
    .Y(_09513_));
 sky130_fd_sc_hd__nand2_1 _19773_ (.A(_09512_),
    .B(_09513_),
    .Y(_09514_));
 sky130_fd_sc_hd__nand2_1 _19774_ (.A(_09381_),
    .B(_09344_),
    .Y(_09516_));
 sky130_fd_sc_hd__xor2_1 _19775_ (.A(_09443_),
    .B(_09516_),
    .X(_09517_));
 sky130_fd_sc_hd__buf_6 _19776_ (.A(_09380_),
    .X(_09518_));
 sky130_fd_sc_hd__nand2_1 _19777_ (.A(_09517_),
    .B(_09518_),
    .Y(_09519_));
 sky130_fd_sc_hd__nand2_1 _19778_ (.A(\div1i.quot[13] ),
    .B(_09435_),
    .Y(_09520_));
 sky130_fd_sc_hd__nand2_1 _19779_ (.A(_09519_),
    .B(_09520_),
    .Y(_09521_));
 sky130_fd_sc_hd__nand2_1 _19780_ (.A(_09521_),
    .B(_06159_),
    .Y(_09522_));
 sky130_fd_sc_hd__nand3_1 _19781_ (.A(_09519_),
    .B(_07318_),
    .C(_09520_),
    .Y(_09523_));
 sky130_fd_sc_hd__nand2_1 _19782_ (.A(_09522_),
    .B(_09523_),
    .Y(_09524_));
 sky130_fd_sc_hd__nor2_1 _19783_ (.A(_09514_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__nand2_1 _19784_ (.A(_09507_),
    .B(_09525_),
    .Y(_09527_));
 sky130_fd_sc_hd__inv_2 _19785_ (.A(_09527_),
    .Y(_09528_));
 sky130_fd_sc_hd__nand2_2 _19786_ (.A(_09429_),
    .B(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__o21ai_1 _19787_ (.A1(_09523_),
    .A2(_09514_),
    .B1(_09512_),
    .Y(_09530_));
 sky130_fd_sc_hd__o21ai_1 _19788_ (.A1(_09505_),
    .A2(_09494_),
    .B1(_09491_),
    .Y(_09531_));
 sky130_fd_sc_hd__a21oi_2 _19789_ (.A1(_09507_),
    .A2(_09530_),
    .B1(_09531_),
    .Y(_09532_));
 sky130_fd_sc_hd__nand2_4 _19790_ (.A(_09529_),
    .B(_09532_),
    .Y(_09533_));
 sky130_fd_sc_hd__nand2_1 _19791_ (.A(_09478_),
    .B(_08824_),
    .Y(_09534_));
 sky130_fd_sc_hd__inv_2 _19792_ (.A(_08813_),
    .Y(_09535_));
 sky130_fd_sc_hd__nand2_1 _19793_ (.A(_09534_),
    .B(_09535_),
    .Y(_09536_));
 sky130_fd_sc_hd__nand3_1 _19794_ (.A(_09478_),
    .B(_08813_),
    .C(_08824_),
    .Y(_09538_));
 sky130_fd_sc_hd__nand2_1 _19795_ (.A(_09536_),
    .B(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__nand2_1 _19796_ (.A(_09539_),
    .B(_07905_),
    .Y(_09540_));
 sky130_fd_sc_hd__nand3_1 _19797_ (.A(_09536_),
    .B(_06772_),
    .C(_09538_),
    .Y(_09541_));
 sky130_fd_sc_hd__nand3_1 _19798_ (.A(_09540_),
    .B(_09541_),
    .C(_09485_),
    .Y(_09542_));
 sky130_fd_sc_hd__nor2_1 _19799_ (.A(_09542_),
    .B(_09467_),
    .Y(_09543_));
 sky130_fd_sc_hd__nand2_2 _19800_ (.A(_09446_),
    .B(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nor2_1 _19801_ (.A(_09542_),
    .B(_09472_),
    .Y(_09545_));
 sky130_fd_sc_hd__nand2_1 _19802_ (.A(_09540_),
    .B(_09541_),
    .Y(_09546_));
 sky130_fd_sc_hd__o21ai_1 _19803_ (.A1(_09483_),
    .A2(_09546_),
    .B1(_09541_),
    .Y(_09547_));
 sky130_fd_sc_hd__nor2_2 _19804_ (.A(_09545_),
    .B(_09547_),
    .Y(_09549_));
 sky130_fd_sc_hd__nand2_2 _19805_ (.A(_09544_),
    .B(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__clkinvlp_2 _19806_ (.A(_09027_),
    .Y(_09551_));
 sky130_fd_sc_hd__inv_2 _19807_ (.A(_09037_),
    .Y(_09552_));
 sky130_fd_sc_hd__nand2_1 _19808_ (.A(_08992_),
    .B(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__nand2_1 _19809_ (.A(_09553_),
    .B(_09036_),
    .Y(_09554_));
 sky130_fd_sc_hd__or2_1 _19810_ (.A(_09551_),
    .B(_09554_),
    .X(_09555_));
 sky130_fd_sc_hd__nand2_1 _19811_ (.A(_09554_),
    .B(_09551_),
    .Y(_09556_));
 sky130_fd_sc_hd__nand2_1 _19812_ (.A(_09555_),
    .B(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__nand2_1 _19813_ (.A(_09557_),
    .B(_07957_),
    .Y(_09558_));
 sky130_fd_sc_hd__nand3_1 _19814_ (.A(_09555_),
    .B(_06827_),
    .C(_09556_),
    .Y(_09560_));
 sky130_fd_sc_hd__nand2_1 _19815_ (.A(_09558_),
    .B(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__or2_1 _19816_ (.A(_09552_),
    .B(_08992_),
    .X(_09562_));
 sky130_fd_sc_hd__nand2_1 _19817_ (.A(_09562_),
    .B(_09553_),
    .Y(_09563_));
 sky130_fd_sc_hd__inv_2 _19818_ (.A(_09563_),
    .Y(_09564_));
 sky130_fd_sc_hd__nand2_1 _19819_ (.A(_09564_),
    .B(_06207_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand2_1 _19820_ (.A(_09563_),
    .B(_08465_),
    .Y(_09566_));
 sky130_fd_sc_hd__nand2_1 _19821_ (.A(_09565_),
    .B(_09566_),
    .Y(_09567_));
 sky130_fd_sc_hd__inv_2 _19822_ (.A(_09567_),
    .Y(_09568_));
 sky130_fd_sc_hd__nand2b_1 _19823_ (.A_N(_09561_),
    .B(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__inv_4 _19824_ (.A(_09569_),
    .Y(_09571_));
 sky130_fd_sc_hd__nand2_1 _19825_ (.A(_09550_),
    .B(_09571_),
    .Y(_09572_));
 sky130_fd_sc_hd__inv_2 _19826_ (.A(_09565_),
    .Y(_09573_));
 sky130_fd_sc_hd__a21boi_2 _19827_ (.A1(_09558_),
    .A2(_09573_),
    .B1_N(_09560_),
    .Y(_09574_));
 sky130_fd_sc_hd__nand2_1 _19828_ (.A(_09572_),
    .B(_09574_),
    .Y(_09575_));
 sky130_fd_sc_hd__inv_2 _19829_ (.A(_09082_),
    .Y(_09576_));
 sky130_fd_sc_hd__nand2_1 _19830_ (.A(_09042_),
    .B(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__nand3_1 _19831_ (.A(_09039_),
    .B(_09041_),
    .C(_09082_),
    .Y(_09578_));
 sky130_fd_sc_hd__nand2_1 _19832_ (.A(_09577_),
    .B(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__inv_2 _19833_ (.A(_09579_),
    .Y(_09580_));
 sky130_fd_sc_hd__nand2_1 _19834_ (.A(_09580_),
    .B(_06819_),
    .Y(_09582_));
 sky130_fd_sc_hd__nand2_1 _19835_ (.A(_09579_),
    .B(_07948_),
    .Y(_09583_));
 sky130_fd_sc_hd__nand2_1 _19836_ (.A(_09582_),
    .B(_09583_),
    .Y(_09584_));
 sky130_fd_sc_hd__inv_2 _19837_ (.A(_09584_),
    .Y(_09585_));
 sky130_fd_sc_hd__nand2_1 _19838_ (.A(_09575_),
    .B(_09585_),
    .Y(_09586_));
 sky130_fd_sc_hd__nand3_1 _19839_ (.A(_09572_),
    .B(_09584_),
    .C(_09574_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand3_1 _19840_ (.A(_09586_),
    .B(_09518_),
    .C(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__nand2_1 _19841_ (.A(\div1i.quot[13] ),
    .B(_09580_),
    .Y(_09589_));
 sky130_fd_sc_hd__nand2_1 _19842_ (.A(_09588_),
    .B(_09589_),
    .Y(_09590_));
 sky130_fd_sc_hd__nand2_1 _19843_ (.A(_09590_),
    .B(_06856_),
    .Y(_09591_));
 sky130_fd_sc_hd__nand3_1 _19844_ (.A(_09588_),
    .B(_06809_),
    .C(_09589_),
    .Y(_09593_));
 sky130_fd_sc_hd__nand2_1 _19845_ (.A(_09591_),
    .B(_09593_),
    .Y(_09594_));
 sky130_fd_sc_hd__nand2_1 _19846_ (.A(_09550_),
    .B(_09568_),
    .Y(_09595_));
 sky130_fd_sc_hd__nand2_1 _19847_ (.A(_09595_),
    .B(_09565_),
    .Y(_09596_));
 sky130_fd_sc_hd__xor2_1 _19848_ (.A(_09561_),
    .B(_09596_),
    .X(_09597_));
 sky130_fd_sc_hd__nand2_1 _19849_ (.A(_09597_),
    .B(_09518_),
    .Y(_09598_));
 sky130_fd_sc_hd__nand2_1 _19850_ (.A(\div1i.quot[13] ),
    .B(_09557_),
    .Y(_09599_));
 sky130_fd_sc_hd__nand2_1 _19851_ (.A(_09598_),
    .B(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__nand2_1 _19852_ (.A(_09600_),
    .B(_06844_),
    .Y(_09601_));
 sky130_fd_sc_hd__nand3_2 _19853_ (.A(_09598_),
    .B(_07400_),
    .C(_09599_),
    .Y(_09602_));
 sky130_fd_sc_hd__nand2_1 _19854_ (.A(_09601_),
    .B(_09602_),
    .Y(_09604_));
 sky130_fd_sc_hd__nor2_1 _19855_ (.A(_09594_),
    .B(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nand3_1 _19856_ (.A(_09544_),
    .B(_09549_),
    .C(_09567_),
    .Y(_09606_));
 sky130_fd_sc_hd__nand3_1 _19857_ (.A(_09595_),
    .B(_09380_),
    .C(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__nand2_1 _19858_ (.A(net238),
    .B(_09564_),
    .Y(_09608_));
 sky130_fd_sc_hd__nand2_1 _19859_ (.A(_09607_),
    .B(_09608_),
    .Y(_09609_));
 sky130_fd_sc_hd__or2_1 _19860_ (.A(_06805_),
    .B(_09609_),
    .X(_09610_));
 sky130_fd_sc_hd__nand2_1 _19861_ (.A(_09609_),
    .B(_06805_),
    .Y(_09611_));
 sky130_fd_sc_hd__nand2_2 _19862_ (.A(_09610_),
    .B(_09611_),
    .Y(_09612_));
 sky130_fd_sc_hd__nand2_1 _19863_ (.A(_09486_),
    .B(_09483_),
    .Y(_09613_));
 sky130_fd_sc_hd__xor2_1 _19864_ (.A(_09546_),
    .B(_09613_),
    .X(_09615_));
 sky130_fd_sc_hd__nand2_1 _19865_ (.A(_09615_),
    .B(_09518_),
    .Y(_09616_));
 sky130_fd_sc_hd__nand2_1 _19866_ (.A(\div1i.quot[13] ),
    .B(_09539_),
    .Y(_09617_));
 sky130_fd_sc_hd__nand2_1 _19867_ (.A(_09616_),
    .B(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__nand2_1 _19868_ (.A(_09618_),
    .B(_06797_),
    .Y(_09619_));
 sky130_fd_sc_hd__nand3_2 _19869_ (.A(_09616_),
    .B(_06799_),
    .C(_09617_),
    .Y(_09620_));
 sky130_fd_sc_hd__nand3b_1 _19870_ (.A_N(_09612_),
    .B(_09619_),
    .C(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__inv_2 _19871_ (.A(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__nand3_4 _19872_ (.A(_09533_),
    .B(_09605_),
    .C(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__inv_2 _19873_ (.A(_09611_),
    .Y(_09624_));
 sky130_fd_sc_hd__o21bai_2 _19874_ (.A1(_09612_),
    .A2(_09620_),
    .B1_N(_09624_),
    .Y(_09626_));
 sky130_fd_sc_hd__o21ai_1 _19875_ (.A1(_09594_),
    .A2(_09602_),
    .B1(_09591_),
    .Y(_09627_));
 sky130_fd_sc_hd__a21oi_1 _19876_ (.A1(_09605_),
    .A2(_09626_),
    .B1(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__nand2_4 _19877_ (.A(_09623_),
    .B(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__nand2_1 _19878_ (.A(_09577_),
    .B(_09080_),
    .Y(_09630_));
 sky130_fd_sc_hd__inv_2 _19879_ (.A(_09073_),
    .Y(_09631_));
 sky130_fd_sc_hd__nand2_1 _19880_ (.A(_09630_),
    .B(_09631_),
    .Y(_09632_));
 sky130_fd_sc_hd__nand3_1 _19881_ (.A(_09577_),
    .B(_09073_),
    .C(_09080_),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2_1 _19882_ (.A(_09632_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__nand2_1 _19883_ (.A(_09634_),
    .B(_08001_),
    .Y(_09635_));
 sky130_fd_sc_hd__nand3_1 _19884_ (.A(_09632_),
    .B(_06874_),
    .C(_09633_),
    .Y(_09637_));
 sky130_fd_sc_hd__nand3_1 _19885_ (.A(_09585_),
    .B(_09635_),
    .C(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__inv_2 _19886_ (.A(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__nand3_2 _19887_ (.A(_09550_),
    .B(_09571_),
    .C(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__inv_2 _19888_ (.A(_09635_),
    .Y(_09641_));
 sky130_fd_sc_hd__o21ai_1 _19889_ (.A1(_09582_),
    .A2(_09641_),
    .B1(_09637_),
    .Y(_09642_));
 sky130_fd_sc_hd__nor2_1 _19890_ (.A(_09574_),
    .B(_09638_),
    .Y(_09643_));
 sky130_fd_sc_hd__nor2_1 _19891_ (.A(_09642_),
    .B(_09643_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand2_1 _19892_ (.A(_09640_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__inv_2 _19893_ (.A(_09088_),
    .Y(_09646_));
 sky130_fd_sc_hd__nand2_1 _19894_ (.A(_09133_),
    .B(_09134_),
    .Y(_09648_));
 sky130_fd_sc_hd__nand2_1 _19895_ (.A(_09646_),
    .B(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__inv_2 _19896_ (.A(_09648_),
    .Y(_09650_));
 sky130_fd_sc_hd__nand2_1 _19897_ (.A(_09088_),
    .B(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__nand2_1 _19898_ (.A(_09649_),
    .B(_09651_),
    .Y(_09652_));
 sky130_fd_sc_hd__nand2_1 _19899_ (.A(_09652_),
    .B(_07450_),
    .Y(_09653_));
 sky130_fd_sc_hd__nand3_2 _19900_ (.A(_09649_),
    .B(_08554_),
    .C(_09651_),
    .Y(_09654_));
 sky130_fd_sc_hd__nand2_1 _19901_ (.A(_09653_),
    .B(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__inv_2 _19902_ (.A(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_1 _19903_ (.A(_09645_),
    .B(_09656_),
    .Y(_09657_));
 sky130_fd_sc_hd__nand3_1 _19904_ (.A(_09640_),
    .B(_09644_),
    .C(_09655_),
    .Y(_09659_));
 sky130_fd_sc_hd__nand3_1 _19905_ (.A(_09657_),
    .B(_09659_),
    .C(_09518_),
    .Y(_09660_));
 sky130_fd_sc_hd__or2_1 _19906_ (.A(_09652_),
    .B(_09380_),
    .X(_09661_));
 sky130_fd_sc_hd__nand2_1 _19907_ (.A(_09660_),
    .B(_09661_),
    .Y(_09662_));
 sky130_fd_sc_hd__or2_1 _19908_ (.A(_06348_),
    .B(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__buf_6 _19909_ (.A(_06348_),
    .X(_09664_));
 sky130_fd_sc_hd__nand2_1 _19910_ (.A(_09662_),
    .B(_09664_),
    .Y(_09665_));
 sky130_fd_sc_hd__nand2_1 _19911_ (.A(_09663_),
    .B(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__inv_2 _19912_ (.A(_09666_),
    .Y(_09667_));
 sky130_fd_sc_hd__nand2_1 _19913_ (.A(_09635_),
    .B(_09637_),
    .Y(_09668_));
 sky130_fd_sc_hd__nand2_1 _19914_ (.A(_09586_),
    .B(_09582_),
    .Y(_09670_));
 sky130_fd_sc_hd__xor2_1 _19915_ (.A(_09668_),
    .B(_09670_),
    .X(_09671_));
 sky130_fd_sc_hd__nand2_1 _19916_ (.A(_09671_),
    .B(_09518_),
    .Y(_09672_));
 sky130_fd_sc_hd__nand2_1 _19917_ (.A(\div1i.quot[13] ),
    .B(_09634_),
    .Y(_09673_));
 sky130_fd_sc_hd__nand2_1 _19918_ (.A(_09672_),
    .B(_09673_),
    .Y(_09674_));
 sky130_fd_sc_hd__nand2_1 _19919_ (.A(_09674_),
    .B(_06903_),
    .Y(_09675_));
 sky130_fd_sc_hd__nand3_2 _19920_ (.A(_09672_),
    .B(_06898_),
    .C(_09673_),
    .Y(_09676_));
 sky130_fd_sc_hd__nand3_1 _19921_ (.A(_09667_),
    .B(_09675_),
    .C(_09676_),
    .Y(_09677_));
 sky130_fd_sc_hd__nand2_1 _19922_ (.A(_09657_),
    .B(_09654_),
    .Y(_09678_));
 sky130_fd_sc_hd__nand2_1 _19923_ (.A(_09651_),
    .B(_09134_),
    .Y(_09679_));
 sky130_fd_sc_hd__xor2_2 _19924_ (.A(_09124_),
    .B(_09679_),
    .X(_09681_));
 sky130_fd_sc_hd__inv_2 _19925_ (.A(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__nand2_1 _19926_ (.A(_09682_),
    .B(_07461_),
    .Y(_09683_));
 sky130_fd_sc_hd__nand2_1 _19927_ (.A(_09681_),
    .B(_08041_),
    .Y(_09684_));
 sky130_fd_sc_hd__nand2_1 _19928_ (.A(_09683_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__inv_2 _19929_ (.A(_09685_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand2_1 _19930_ (.A(_09678_),
    .B(_09686_),
    .Y(_09687_));
 sky130_fd_sc_hd__nand3_1 _19931_ (.A(_09657_),
    .B(_09685_),
    .C(_09654_),
    .Y(_09688_));
 sky130_fd_sc_hd__nand2_1 _19932_ (.A(_09687_),
    .B(_09688_),
    .Y(_09689_));
 sky130_fd_sc_hd__nand2_1 _19933_ (.A(_09689_),
    .B(_09518_),
    .Y(_09690_));
 sky130_fd_sc_hd__nand2_1 _19934_ (.A(_09681_),
    .B(\div1i.quot[13] ),
    .Y(_09692_));
 sky130_fd_sc_hd__nand2_1 _19935_ (.A(_09690_),
    .B(_09692_),
    .Y(_09693_));
 sky130_fd_sc_hd__nand2_1 _19936_ (.A(_09693_),
    .B(_07474_),
    .Y(_09694_));
 sky130_fd_sc_hd__nand3_2 _19937_ (.A(_09690_),
    .B(_06366_),
    .C(_09692_),
    .Y(_09695_));
 sky130_fd_sc_hd__nand2_1 _19938_ (.A(_09694_),
    .B(_09695_),
    .Y(_09696_));
 sky130_fd_sc_hd__inv_2 _19939_ (.A(_09696_),
    .Y(_09697_));
 sky130_fd_sc_hd__nand3_1 _19940_ (.A(_09683_),
    .B(_09684_),
    .C(_09656_),
    .Y(_09698_));
 sky130_fd_sc_hd__inv_2 _19941_ (.A(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__nand2_1 _19942_ (.A(_09699_),
    .B(_09645_),
    .Y(_09700_));
 sky130_fd_sc_hd__inv_2 _19943_ (.A(_09684_),
    .Y(_09701_));
 sky130_fd_sc_hd__o21a_1 _19944_ (.A1(_09654_),
    .A2(_09701_),
    .B1(_09683_),
    .X(_09703_));
 sky130_fd_sc_hd__nand2_1 _19945_ (.A(_09700_),
    .B(_09703_),
    .Y(_09704_));
 sky130_fd_sc_hd__o21bai_1 _19946_ (.A1(_09135_),
    .A2(_09646_),
    .B1_N(_09185_),
    .Y(_09705_));
 sky130_fd_sc_hd__or2_1 _19947_ (.A(_09156_),
    .B(_09705_),
    .X(_09706_));
 sky130_fd_sc_hd__nand2_1 _19948_ (.A(_09705_),
    .B(_09156_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand2_1 _19949_ (.A(_09706_),
    .B(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__inv_2 _19950_ (.A(_09708_),
    .Y(_09709_));
 sky130_fd_sc_hd__nand2_1 _19951_ (.A(_09709_),
    .B(_06936_),
    .Y(_09710_));
 sky130_fd_sc_hd__nand2_1 _19952_ (.A(_09708_),
    .B(_08611_),
    .Y(_09711_));
 sky130_fd_sc_hd__nand2_1 _19953_ (.A(_09710_),
    .B(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__inv_2 _19954_ (.A(_09712_),
    .Y(_09714_));
 sky130_fd_sc_hd__nand2_1 _19955_ (.A(_09704_),
    .B(_09714_),
    .Y(_09715_));
 sky130_fd_sc_hd__nand3_1 _19956_ (.A(_09700_),
    .B(_09703_),
    .C(_09712_),
    .Y(_09716_));
 sky130_fd_sc_hd__nand3_2 _19957_ (.A(_09715_),
    .B(_09716_),
    .C(_09518_),
    .Y(_09717_));
 sky130_fd_sc_hd__nand2_1 _19958_ (.A(_09709_),
    .B(\div1i.quot[13] ),
    .Y(_09718_));
 sky130_fd_sc_hd__nand2_1 _19959_ (.A(_09717_),
    .B(_09718_),
    .Y(_09719_));
 sky130_fd_sc_hd__nand2_1 _19960_ (.A(_09719_),
    .B(_06947_),
    .Y(_09720_));
 sky130_fd_sc_hd__nand3_2 _19961_ (.A(_09717_),
    .B(_06949_),
    .C(_09718_),
    .Y(_09721_));
 sky130_fd_sc_hd__nand2_4 _19962_ (.A(_09721_),
    .B(_09720_),
    .Y(_09722_));
 sky130_fd_sc_hd__inv_2 _19963_ (.A(_09722_),
    .Y(_09723_));
 sky130_fd_sc_hd__nand2_1 _19964_ (.A(_09697_),
    .B(_09723_),
    .Y(_09725_));
 sky130_fd_sc_hd__nor2_1 _19965_ (.A(_09677_),
    .B(_09725_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand2_4 _19966_ (.A(_09629_),
    .B(_09726_),
    .Y(_09727_));
 sky130_fd_sc_hd__o21ai_1 _19967_ (.A1(_09666_),
    .A2(_09676_),
    .B1(_09665_),
    .Y(_09728_));
 sky130_fd_sc_hd__nor2_1 _19968_ (.A(_09722_),
    .B(_09696_),
    .Y(_09729_));
 sky130_fd_sc_hd__inv_2 _19969_ (.A(_09721_),
    .Y(_09730_));
 sky130_fd_sc_hd__o21ai_1 _19970_ (.A1(_09695_),
    .A2(_09730_),
    .B1(_09720_),
    .Y(_09731_));
 sky130_fd_sc_hd__a21oi_2 _19971_ (.A1(_09728_),
    .A2(_09729_),
    .B1(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__nand2_2 _19972_ (.A(_09727_),
    .B(_09732_),
    .Y(_09733_));
 sky130_fd_sc_hd__nand2_2 _19973_ (.A(_09707_),
    .B(_09154_),
    .Y(_09734_));
 sky130_fd_sc_hd__xor2_4 _19974_ (.A(_09180_),
    .B(_09734_),
    .X(_09736_));
 sky130_fd_sc_hd__nand3_2 _19975_ (.A(_09715_),
    .B(_09518_),
    .C(_09710_),
    .Y(_09737_));
 sky130_fd_sc_hd__xor2_4 _19976_ (.A(_09736_),
    .B(_09737_),
    .X(_09738_));
 sky130_fd_sc_hd__clkinvlp_2 _19977_ (.A(_09738_),
    .Y(_09739_));
 sky130_fd_sc_hd__nand2_4 _19978_ (.A(_09733_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nand3_4 _19979_ (.A(_09727_),
    .B(_09732_),
    .C(_09738_),
    .Y(_09741_));
 sky130_fd_sc_hd__nand2_8 _19980_ (.A(_09740_),
    .B(_09741_),
    .Y(_09742_));
 sky130_fd_sc_hd__buf_8 _19981_ (.A(_09742_),
    .X(_09743_));
 sky130_fd_sc_hd__buf_6 _19982_ (.A(net224),
    .X(\div1i.quot[12] ));
 sky130_fd_sc_hd__nand2_1 _19983_ (.A(_09333_),
    .B(_09421_),
    .Y(_09744_));
 sky130_fd_sc_hd__inv_2 _19984_ (.A(_09425_),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_1 _19985_ (.A(_09744_),
    .B(_09746_),
    .Y(_09747_));
 sky130_fd_sc_hd__inv_2 _19986_ (.A(_09400_),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_2 _19987_ (.A(_09747_),
    .B(_09748_),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_1 _19988_ (.A(_09749_),
    .B(_09399_),
    .Y(_09750_));
 sky130_fd_sc_hd__inv_2 _19989_ (.A(_09388_),
    .Y(_09751_));
 sky130_fd_sc_hd__nand2_1 _19990_ (.A(_09750_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__nand3_1 _19991_ (.A(_09749_),
    .B(_09388_),
    .C(_09399_),
    .Y(_09753_));
 sky130_fd_sc_hd__nand2_1 _19992_ (.A(_09752_),
    .B(_09753_),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_1 _19993_ (.A(_09754_),
    .B(_07226_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand3_1 _19994_ (.A(_09744_),
    .B(_09400_),
    .C(_09746_),
    .Y(_09757_));
 sky130_fd_sc_hd__nand3_2 _19995_ (.A(_09749_),
    .B(_07128_),
    .C(_09757_),
    .Y(_09758_));
 sky130_fd_sc_hd__inv_2 _19996_ (.A(_09758_),
    .Y(_09759_));
 sky130_fd_sc_hd__nand3_2 _19997_ (.A(_09752_),
    .B(_07228_),
    .C(_09753_),
    .Y(_09760_));
 sky130_fd_sc_hd__nand3_1 _19998_ (.A(_09755_),
    .B(_09759_),
    .C(_09760_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_1 _19999_ (.A(_09761_),
    .B(_09760_),
    .Y(_09762_));
 sky130_fd_sc_hd__inv_2 _20000_ (.A(_09420_),
    .Y(_09763_));
 sky130_fd_sc_hd__nand2_1 _20001_ (.A(_09333_),
    .B(_09763_),
    .Y(_09764_));
 sky130_fd_sc_hd__nand2_1 _20002_ (.A(_09764_),
    .B(_09418_),
    .Y(_09765_));
 sky130_fd_sc_hd__inv_2 _20003_ (.A(_09409_),
    .Y(_09766_));
 sky130_fd_sc_hd__nand2_1 _20004_ (.A(_09765_),
    .B(_09766_),
    .Y(_09768_));
 sky130_fd_sc_hd__nand3_1 _20005_ (.A(_09764_),
    .B(_09409_),
    .C(_09418_),
    .Y(_09769_));
 sky130_fd_sc_hd__nand2_1 _20006_ (.A(_09768_),
    .B(_09769_),
    .Y(_09770_));
 sky130_fd_sc_hd__nand2_1 _20007_ (.A(_09770_),
    .B(_07146_),
    .Y(_09771_));
 sky130_fd_sc_hd__or2_1 _20008_ (.A(_09763_),
    .B(_09333_),
    .X(_09772_));
 sky130_fd_sc_hd__nand2_1 _20009_ (.A(_09772_),
    .B(_09764_),
    .Y(_09773_));
 sky130_fd_sc_hd__inv_2 _20010_ (.A(_09773_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand2_1 _20011_ (.A(_09774_),
    .B(_07157_),
    .Y(_09775_));
 sky130_fd_sc_hd__inv_2 _20012_ (.A(_09775_),
    .Y(_09776_));
 sky130_fd_sc_hd__inv_2 _20013_ (.A(_09770_),
    .Y(_09777_));
 sky130_fd_sc_hd__nand2_1 _20014_ (.A(_09777_),
    .B(_07149_),
    .Y(_09779_));
 sky130_fd_sc_hd__inv_2 _20015_ (.A(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__a21oi_2 _20016_ (.A1(_09771_),
    .A2(_09776_),
    .B1(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__nand2_1 _20017_ (.A(_09749_),
    .B(_09757_),
    .Y(_09782_));
 sky130_fd_sc_hd__nand2_1 _20018_ (.A(_09782_),
    .B(_07130_),
    .Y(_09783_));
 sky130_fd_sc_hd__nand2_1 _20019_ (.A(_09783_),
    .B(_09758_),
    .Y(_09784_));
 sky130_fd_sc_hd__inv_2 _20020_ (.A(_09784_),
    .Y(_09785_));
 sky130_fd_sc_hd__nand3_1 _20021_ (.A(_09755_),
    .B(_09785_),
    .C(_09760_),
    .Y(_09786_));
 sky130_fd_sc_hd__nor2_1 _20022_ (.A(_09781_),
    .B(_09786_),
    .Y(_09787_));
 sky130_fd_sc_hd__nor2_1 _20023_ (.A(_09762_),
    .B(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__inv_2 _20024_ (.A(_09786_),
    .Y(_09790_));
 sky130_fd_sc_hd__nand2_1 _20025_ (.A(_09224_),
    .B(_09227_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand2_1 _20026_ (.A(_09791_),
    .B(_09230_),
    .Y(_09792_));
 sky130_fd_sc_hd__nand2_1 _20027_ (.A(_09792_),
    .B(_09232_),
    .Y(_09793_));
 sky130_fd_sc_hd__nand2_1 _20028_ (.A(_09793_),
    .B(_06982_),
    .Y(_09794_));
 sky130_fd_sc_hd__o21ai_1 _20029_ (.A1(_09215_),
    .A2(\div1i.quot[13] ),
    .B1(_09228_),
    .Y(_09795_));
 sky130_fd_sc_hd__nand3_1 _20030_ (.A(_09792_),
    .B(_06984_),
    .C(_09232_),
    .Y(_09796_));
 sky130_fd_sc_hd__inv_2 _20031_ (.A(_09796_),
    .Y(_09797_));
 sky130_fd_sc_hd__a21o_1 _20032_ (.A1(_09794_),
    .A2(_09795_),
    .B1(_09797_),
    .X(_09798_));
 sky130_fd_sc_hd__nand2_1 _20033_ (.A(_09233_),
    .B(_09214_),
    .Y(_09799_));
 sky130_fd_sc_hd__nand2_1 _20034_ (.A(_09232_),
    .B(_09224_),
    .Y(_09801_));
 sky130_fd_sc_hd__xor2_2 _20035_ (.A(_09799_),
    .B(_09801_),
    .X(_09802_));
 sky130_fd_sc_hd__nand2_1 _20036_ (.A(_09802_),
    .B(_07043_),
    .Y(_09803_));
 sky130_fd_sc_hd__nand2_1 _20037_ (.A(_09798_),
    .B(_09803_),
    .Y(_09804_));
 sky130_fd_sc_hd__inv_2 _20038_ (.A(_09802_),
    .Y(_09805_));
 sky130_fd_sc_hd__nand2_1 _20039_ (.A(_09805_),
    .B(_07048_),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_1 _20040_ (.A(_09804_),
    .B(_09806_),
    .Y(_09807_));
 sky130_fd_sc_hd__nand2_1 _20041_ (.A(_09226_),
    .B(_09232_),
    .Y(_09808_));
 sky130_fd_sc_hd__nand2_1 _20042_ (.A(_09808_),
    .B(_09233_),
    .Y(_09809_));
 sky130_fd_sc_hd__nand2_1 _20043_ (.A(_09809_),
    .B(_09321_),
    .Y(_09810_));
 sky130_fd_sc_hd__nand3_2 _20044_ (.A(_09808_),
    .B(_09233_),
    .C(_09322_),
    .Y(_09812_));
 sky130_fd_sc_hd__nand2_1 _20045_ (.A(_09810_),
    .B(_09812_),
    .Y(_09813_));
 sky130_fd_sc_hd__nand2_1 _20046_ (.A(_09813_),
    .B(_07031_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand3_1 _20047_ (.A(_09810_),
    .B(_07034_),
    .C(_09812_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand2_1 _20048_ (.A(_09814_),
    .B(_09815_),
    .Y(_09816_));
 sky130_fd_sc_hd__inv_2 _20049_ (.A(_09816_),
    .Y(_09817_));
 sky130_fd_sc_hd__nand2_1 _20050_ (.A(_09807_),
    .B(_09817_),
    .Y(_09818_));
 sky130_fd_sc_hd__nand2_1 _20051_ (.A(_09818_),
    .B(_09815_),
    .Y(_09819_));
 sky130_fd_sc_hd__nand2_1 _20052_ (.A(_09812_),
    .B(_09319_),
    .Y(_09820_));
 sky130_fd_sc_hd__xor2_2 _20053_ (.A(_09311_),
    .B(_09820_),
    .X(_09821_));
 sky130_fd_sc_hd__buf_6 _20054_ (.A(_06465_),
    .X(_09823_));
 sky130_fd_sc_hd__nand2_1 _20055_ (.A(_09821_),
    .B(_09823_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_1 _20056_ (.A(_09819_),
    .B(_09824_),
    .Y(_09825_));
 sky130_fd_sc_hd__or2_1 _20057_ (.A(_06465_),
    .B(_09821_),
    .X(_09826_));
 sky130_fd_sc_hd__nand2_1 _20058_ (.A(_09825_),
    .B(_09826_),
    .Y(_09827_));
 sky130_fd_sc_hd__nor2_1 _20059_ (.A(_09311_),
    .B(_09321_),
    .Y(_09828_));
 sky130_fd_sc_hd__nand3_1 _20060_ (.A(_09808_),
    .B(_09828_),
    .C(_09233_),
    .Y(_09829_));
 sky130_fd_sc_hd__inv_2 _20061_ (.A(_09327_),
    .Y(_09830_));
 sky130_fd_sc_hd__nand2_1 _20062_ (.A(_09829_),
    .B(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__nand2_2 _20063_ (.A(_09831_),
    .B(_09299_),
    .Y(_09832_));
 sky130_fd_sc_hd__nand2_1 _20064_ (.A(_09832_),
    .B(_09296_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_1 _20065_ (.A(_09834_),
    .B(_09289_),
    .Y(_09835_));
 sky130_fd_sc_hd__nand3_1 _20066_ (.A(_09832_),
    .B(_09288_),
    .C(_09296_),
    .Y(_09836_));
 sky130_fd_sc_hd__nand2_1 _20067_ (.A(_09835_),
    .B(_09836_),
    .Y(_09837_));
 sky130_fd_sc_hd__nand2_1 _20068_ (.A(_09837_),
    .B(_08738_),
    .Y(_09838_));
 sky130_fd_sc_hd__nand3_1 _20069_ (.A(_09829_),
    .B(_09298_),
    .C(_09830_),
    .Y(_09839_));
 sky130_fd_sc_hd__nand2_1 _20070_ (.A(_09832_),
    .B(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__nand2_1 _20071_ (.A(_09840_),
    .B(_07024_),
    .Y(_09841_));
 sky130_fd_sc_hd__nand3_2 _20072_ (.A(_09832_),
    .B(_07021_),
    .C(_09839_),
    .Y(_09842_));
 sky130_fd_sc_hd__nand2_1 _20073_ (.A(_09841_),
    .B(_09842_),
    .Y(_09843_));
 sky130_fd_sc_hd__inv_2 _20074_ (.A(_09843_),
    .Y(_09845_));
 sky130_fd_sc_hd__nand3_1 _20075_ (.A(_09835_),
    .B(_05896_),
    .C(_09836_),
    .Y(_09846_));
 sky130_fd_sc_hd__nand3_1 _20076_ (.A(_09838_),
    .B(_09845_),
    .C(_09846_),
    .Y(_09847_));
 sky130_fd_sc_hd__inv_2 _20077_ (.A(_09847_),
    .Y(_09848_));
 sky130_fd_sc_hd__nand2_1 _20078_ (.A(_09827_),
    .B(_09848_),
    .Y(_09849_));
 sky130_fd_sc_hd__inv_2 _20079_ (.A(_09842_),
    .Y(_09850_));
 sky130_fd_sc_hd__a21boi_1 _20080_ (.A1(_09838_),
    .A2(_09850_),
    .B1_N(_09846_),
    .Y(_09851_));
 sky130_fd_sc_hd__nand2_1 _20081_ (.A(_09849_),
    .B(_09851_),
    .Y(_09852_));
 sky130_fd_sc_hd__nand2_1 _20082_ (.A(_09779_),
    .B(_09771_),
    .Y(_09853_));
 sky130_fd_sc_hd__inv_2 _20083_ (.A(_09853_),
    .Y(_09854_));
 sky130_fd_sc_hd__nand2_1 _20084_ (.A(_09773_),
    .B(_07155_),
    .Y(_09856_));
 sky130_fd_sc_hd__nand2_1 _20085_ (.A(_09775_),
    .B(_09856_),
    .Y(_09857_));
 sky130_fd_sc_hd__inv_4 _20086_ (.A(_09857_),
    .Y(_09858_));
 sky130_fd_sc_hd__nand2_1 _20087_ (.A(_09854_),
    .B(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__inv_2 _20088_ (.A(_09859_),
    .Y(_09860_));
 sky130_fd_sc_hd__nand3_1 _20089_ (.A(_09790_),
    .B(_09852_),
    .C(_09860_),
    .Y(_09861_));
 sky130_fd_sc_hd__nand2_2 _20090_ (.A(_09788_),
    .B(_09861_),
    .Y(_09862_));
 sky130_fd_sc_hd__inv_2 _20091_ (.A(_09514_),
    .Y(_09863_));
 sky130_fd_sc_hd__inv_2 _20092_ (.A(_09524_),
    .Y(_09864_));
 sky130_fd_sc_hd__nand2_1 _20093_ (.A(_09429_),
    .B(_09864_),
    .Y(_09865_));
 sky130_fd_sc_hd__nand2_1 _20094_ (.A(_09865_),
    .B(_09523_),
    .Y(_09867_));
 sky130_fd_sc_hd__or2_1 _20095_ (.A(_09863_),
    .B(_09867_),
    .X(_09868_));
 sky130_fd_sc_hd__nand2_1 _20096_ (.A(_09867_),
    .B(_09863_),
    .Y(_09869_));
 sky130_fd_sc_hd__nand2_1 _20097_ (.A(_09868_),
    .B(_09869_),
    .Y(_09870_));
 sky130_fd_sc_hd__nand2_1 _20098_ (.A(_09870_),
    .B(_07247_),
    .Y(_09871_));
 sky130_fd_sc_hd__nand3_1 _20099_ (.A(_09868_),
    .B(_07249_),
    .C(_09869_),
    .Y(_09872_));
 sky130_fd_sc_hd__nand2_1 _20100_ (.A(_09871_),
    .B(_09872_),
    .Y(_09873_));
 sky130_fd_sc_hd__inv_2 _20101_ (.A(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__or2_1 _20102_ (.A(_09864_),
    .B(_09429_),
    .X(_09875_));
 sky130_fd_sc_hd__nand2_1 _20103_ (.A(_09875_),
    .B(_09865_),
    .Y(_09876_));
 sky130_fd_sc_hd__inv_2 _20104_ (.A(_09876_),
    .Y(_09878_));
 sky130_fd_sc_hd__nand2_2 _20105_ (.A(_09878_),
    .B(_06521_),
    .Y(_09879_));
 sky130_fd_sc_hd__nand2_1 _20106_ (.A(_09876_),
    .B(_07677_),
    .Y(_09880_));
 sky130_fd_sc_hd__nand2_1 _20107_ (.A(_09879_),
    .B(_09880_),
    .Y(_09881_));
 sky130_fd_sc_hd__inv_2 _20108_ (.A(_09881_),
    .Y(_09882_));
 sky130_fd_sc_hd__nand2_1 _20109_ (.A(_09874_),
    .B(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__inv_2 _20110_ (.A(_09883_),
    .Y(_09884_));
 sky130_fd_sc_hd__nand2_1 _20111_ (.A(_09862_),
    .B(_09884_),
    .Y(_09885_));
 sky130_fd_sc_hd__inv_2 _20112_ (.A(_09879_),
    .Y(_09886_));
 sky130_fd_sc_hd__a21boi_2 _20113_ (.A1(_09871_),
    .A2(_09886_),
    .B1_N(_09872_),
    .Y(_09887_));
 sky130_fd_sc_hd__nand2_1 _20114_ (.A(_09885_),
    .B(_09887_),
    .Y(_09889_));
 sky130_fd_sc_hd__nand2_1 _20115_ (.A(_09429_),
    .B(_09525_),
    .Y(_09890_));
 sky130_fd_sc_hd__inv_2 _20116_ (.A(_09530_),
    .Y(_09891_));
 sky130_fd_sc_hd__nand2_1 _20117_ (.A(_09890_),
    .B(_09891_),
    .Y(_09892_));
 sky130_fd_sc_hd__inv_2 _20118_ (.A(_09506_),
    .Y(_09893_));
 sky130_fd_sc_hd__nand2_1 _20119_ (.A(_09892_),
    .B(_09893_),
    .Y(_09894_));
 sky130_fd_sc_hd__nand3_1 _20120_ (.A(_09890_),
    .B(_09506_),
    .C(_09891_),
    .Y(_09895_));
 sky130_fd_sc_hd__nand2_1 _20121_ (.A(_09894_),
    .B(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__inv_2 _20122_ (.A(_09896_),
    .Y(_09897_));
 sky130_fd_sc_hd__nand2_1 _20123_ (.A(_09897_),
    .B(_07278_),
    .Y(_09898_));
 sky130_fd_sc_hd__nand2_1 _20124_ (.A(_09896_),
    .B(_07276_),
    .Y(_09900_));
 sky130_fd_sc_hd__nand2_1 _20125_ (.A(_09898_),
    .B(_09900_),
    .Y(_09901_));
 sky130_fd_sc_hd__inv_2 _20126_ (.A(_09901_),
    .Y(_09902_));
 sky130_fd_sc_hd__nand2_1 _20127_ (.A(_09889_),
    .B(_09902_),
    .Y(_09903_));
 sky130_fd_sc_hd__inv_6 _20128_ (.A(_09742_),
    .Y(_09904_));
 sky130_fd_sc_hd__nand3_1 _20129_ (.A(_09885_),
    .B(_09901_),
    .C(_09887_),
    .Y(_09905_));
 sky130_fd_sc_hd__nand3_1 _20130_ (.A(_09903_),
    .B(_09904_),
    .C(_09905_),
    .Y(_09906_));
 sky130_fd_sc_hd__nand2_1 _20131_ (.A(net224),
    .B(_09897_),
    .Y(_09907_));
 sky130_fd_sc_hd__nand2_1 _20132_ (.A(_09906_),
    .B(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__nand2_1 _20133_ (.A(_09908_),
    .B(_06554_),
    .Y(_09909_));
 sky130_fd_sc_hd__nand3_1 _20134_ (.A(_09906_),
    .B(_06556_),
    .C(_09907_),
    .Y(_09911_));
 sky130_fd_sc_hd__nand2_1 _20135_ (.A(_09909_),
    .B(_09911_),
    .Y(_09912_));
 sky130_fd_sc_hd__nand2_1 _20136_ (.A(_09862_),
    .B(_09882_),
    .Y(_09913_));
 sky130_fd_sc_hd__nand2_1 _20137_ (.A(_09913_),
    .B(_09879_),
    .Y(_09914_));
 sky130_fd_sc_hd__nand2_1 _20138_ (.A(_09914_),
    .B(_09874_),
    .Y(_09915_));
 sky130_fd_sc_hd__nand3_1 _20139_ (.A(_09913_),
    .B(_09873_),
    .C(_09879_),
    .Y(_09916_));
 sky130_fd_sc_hd__nand2_1 _20140_ (.A(_09915_),
    .B(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__nand2_1 _20141_ (.A(_09917_),
    .B(_09904_),
    .Y(_09918_));
 sky130_fd_sc_hd__nand2_1 _20142_ (.A(net224),
    .B(_09870_),
    .Y(_09919_));
 sky130_fd_sc_hd__nand2_1 _20143_ (.A(_09918_),
    .B(_09919_),
    .Y(_09920_));
 sky130_fd_sc_hd__nand2_1 _20144_ (.A(_09920_),
    .B(_06568_),
    .Y(_09922_));
 sky130_fd_sc_hd__nand3_2 _20145_ (.A(_09918_),
    .B(_06570_),
    .C(_09919_),
    .Y(_09923_));
 sky130_fd_sc_hd__nand2_1 _20146_ (.A(_09922_),
    .B(_09923_),
    .Y(_09924_));
 sky130_fd_sc_hd__nor2_1 _20147_ (.A(_09912_),
    .B(_09924_),
    .Y(_09925_));
 sky130_fd_sc_hd__nand2_1 _20148_ (.A(_09860_),
    .B(_09852_),
    .Y(_09926_));
 sky130_fd_sc_hd__nand2_1 _20149_ (.A(_09926_),
    .B(_09781_),
    .Y(_09927_));
 sky130_fd_sc_hd__nand2_1 _20150_ (.A(_09927_),
    .B(_09785_),
    .Y(_09928_));
 sky130_fd_sc_hd__nand2_1 _20151_ (.A(_09928_),
    .B(_09758_),
    .Y(_09929_));
 sky130_fd_sc_hd__nand3_1 _20152_ (.A(_09929_),
    .B(_09760_),
    .C(_09755_),
    .Y(_09930_));
 sky130_fd_sc_hd__nand2_1 _20153_ (.A(_09755_),
    .B(_09760_),
    .Y(_09931_));
 sky130_fd_sc_hd__nand3_1 _20154_ (.A(_09928_),
    .B(_09758_),
    .C(_09931_),
    .Y(_09933_));
 sky130_fd_sc_hd__nand2_1 _20155_ (.A(_09930_),
    .B(_09933_),
    .Y(_09934_));
 sky130_fd_sc_hd__nand2_1 _20156_ (.A(_09934_),
    .B(_09904_),
    .Y(_09935_));
 sky130_fd_sc_hd__nand2_1 _20157_ (.A(net224),
    .B(_09754_),
    .Y(_09936_));
 sky130_fd_sc_hd__nand3_2 _20158_ (.A(_09935_),
    .B(_07318_),
    .C(_09936_),
    .Y(_09937_));
 sky130_fd_sc_hd__or2_1 _20159_ (.A(_09882_),
    .B(_09862_),
    .X(_09938_));
 sky130_fd_sc_hd__nand3_1 _20160_ (.A(_09938_),
    .B(_09904_),
    .C(_09913_),
    .Y(_09939_));
 sky130_fd_sc_hd__nand2_1 _20161_ (.A(net224),
    .B(_09878_),
    .Y(_09940_));
 sky130_fd_sc_hd__nand3_1 _20162_ (.A(_09939_),
    .B(_06592_),
    .C(_09940_),
    .Y(_09941_));
 sky130_fd_sc_hd__inv_2 _20163_ (.A(_09941_),
    .Y(_09942_));
 sky130_fd_sc_hd__buf_6 _20164_ (.A(_06592_),
    .X(_09944_));
 sky130_fd_sc_hd__a21o_1 _20165_ (.A1(_09939_),
    .A2(_09940_),
    .B1(_09944_),
    .X(_09945_));
 sky130_fd_sc_hd__o21ai_2 _20166_ (.A1(_09937_),
    .A2(_09942_),
    .B1(_09945_),
    .Y(_09946_));
 sky130_fd_sc_hd__inv_2 _20167_ (.A(_09911_),
    .Y(_09947_));
 sky130_fd_sc_hd__o21ai_1 _20168_ (.A1(_09923_),
    .A2(_09947_),
    .B1(_09909_),
    .Y(_09948_));
 sky130_fd_sc_hd__a21oi_1 _20169_ (.A1(_09925_),
    .A2(_09946_),
    .B1(_09948_),
    .Y(_09949_));
 sky130_fd_sc_hd__inv_2 _20170_ (.A(_09793_),
    .Y(_09950_));
 sky130_fd_sc_hd__nand2_1 _20171_ (.A(_09743_),
    .B(_09950_),
    .Y(_09951_));
 sky130_fd_sc_hd__nand2_1 _20172_ (.A(_09794_),
    .B(_09796_),
    .Y(_09952_));
 sky130_fd_sc_hd__xor2_1 _20173_ (.A(_09795_),
    .B(_09952_),
    .X(_09953_));
 sky130_fd_sc_hd__nand3b_1 _20174_ (.A_N(_09953_),
    .B(_09740_),
    .C(_09741_),
    .Y(_09955_));
 sky130_fd_sc_hd__nand2_1 _20175_ (.A(_09951_),
    .B(_09955_),
    .Y(_09956_));
 sky130_fd_sc_hd__nand2_1 _20176_ (.A(_09956_),
    .B(_08857_),
    .Y(_09957_));
 sky130_fd_sc_hd__nor2_1 _20177_ (.A(_09215_),
    .B(_09518_),
    .Y(_09958_));
 sky130_fd_sc_hd__or2_1 _20178_ (.A(_06607_),
    .B(_09958_),
    .X(_09959_));
 sky130_fd_sc_hd__nand2_1 _20179_ (.A(_09959_),
    .B(_09230_),
    .Y(_09960_));
 sky130_fd_sc_hd__inv_2 _20180_ (.A(_09960_),
    .Y(_09961_));
 sky130_fd_sc_hd__nand2_1 _20181_ (.A(_09742_),
    .B(_09961_),
    .Y(_09962_));
 sky130_fd_sc_hd__nand3_1 _20182_ (.A(_09740_),
    .B(_09741_),
    .C(_09958_),
    .Y(_09963_));
 sky130_fd_sc_hd__nand2_1 _20183_ (.A(_09962_),
    .B(_09963_),
    .Y(_09964_));
 sky130_fd_sc_hd__nand2_2 _20184_ (.A(_09964_),
    .B(_06615_),
    .Y(_09966_));
 sky130_fd_sc_hd__nand2_1 _20185_ (.A(_09957_),
    .B(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__inv_2 _20186_ (.A(_09967_),
    .Y(_09968_));
 sky130_fd_sc_hd__nand3_1 _20187_ (.A(_09962_),
    .B(_06620_),
    .C(_09963_),
    .Y(_09969_));
 sky130_fd_sc_hd__nand3_2 _20188_ (.A(_09743_),
    .B(_09228_),
    .C(_07004_),
    .Y(_09970_));
 sky130_fd_sc_hd__inv_2 _20189_ (.A(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__nand3_4 _20190_ (.A(_09966_),
    .B(_09969_),
    .C(_09971_),
    .Y(_09972_));
 sky130_fd_sc_hd__or2_1 _20191_ (.A(_08857_),
    .B(_09956_),
    .X(_09973_));
 sky130_fd_sc_hd__a21boi_2 _20192_ (.A1(_09968_),
    .A2(_09972_),
    .B1_N(_09973_),
    .Y(_09974_));
 sky130_fd_sc_hd__clkinvlp_2 _20193_ (.A(_09840_),
    .Y(_09975_));
 sky130_fd_sc_hd__nand2_1 _20194_ (.A(_09742_),
    .B(_09975_),
    .Y(_09977_));
 sky130_fd_sc_hd__nand2_1 _20195_ (.A(_09827_),
    .B(_09845_),
    .Y(_09978_));
 sky130_fd_sc_hd__nand3_1 _20196_ (.A(_09825_),
    .B(_09843_),
    .C(_09826_),
    .Y(_09979_));
 sky130_fd_sc_hd__nand2_1 _20197_ (.A(_09978_),
    .B(_09979_),
    .Y(_09980_));
 sky130_fd_sc_hd__inv_2 _20198_ (.A(_09980_),
    .Y(_09981_));
 sky130_fd_sc_hd__nand3_1 _20199_ (.A(_09740_),
    .B(_09741_),
    .C(_09981_),
    .Y(_09982_));
 sky130_fd_sc_hd__nand2_1 _20200_ (.A(_09977_),
    .B(_09982_),
    .Y(_09983_));
 sky130_fd_sc_hd__nand2_1 _20201_ (.A(_09983_),
    .B(_06636_),
    .Y(_09984_));
 sky130_fd_sc_hd__nand3_1 _20202_ (.A(_09977_),
    .B(_06639_),
    .C(_09982_),
    .Y(_09985_));
 sky130_fd_sc_hd__nand2_1 _20203_ (.A(_09984_),
    .B(_09985_),
    .Y(_09986_));
 sky130_fd_sc_hd__clkinvlp_2 _20204_ (.A(_09986_),
    .Y(_09988_));
 sky130_fd_sc_hd__nand2_1 _20205_ (.A(_09743_),
    .B(_09821_),
    .Y(_09989_));
 sky130_fd_sc_hd__nand2_1 _20206_ (.A(_09826_),
    .B(_09824_),
    .Y(_09990_));
 sky130_fd_sc_hd__xor2_1 _20207_ (.A(_09819_),
    .B(_09990_),
    .X(_09991_));
 sky130_fd_sc_hd__nand3_1 _20208_ (.A(_09740_),
    .B(_09741_),
    .C(_09991_),
    .Y(_09992_));
 sky130_fd_sc_hd__nand2_1 _20209_ (.A(_09989_),
    .B(_09992_),
    .Y(_09993_));
 sky130_fd_sc_hd__nand2_1 _20210_ (.A(_09993_),
    .B(_06648_),
    .Y(_09994_));
 sky130_fd_sc_hd__nand3_2 _20211_ (.A(_09989_),
    .B(_06651_),
    .C(_09992_),
    .Y(_09995_));
 sky130_fd_sc_hd__nand2_2 _20212_ (.A(_09994_),
    .B(_09995_),
    .Y(_09996_));
 sky130_fd_sc_hd__inv_2 _20213_ (.A(_09996_),
    .Y(_09997_));
 sky130_fd_sc_hd__nand2_1 _20214_ (.A(_09988_),
    .B(_09997_),
    .Y(_09999_));
 sky130_fd_sc_hd__inv_2 _20215_ (.A(_09813_),
    .Y(_10000_));
 sky130_fd_sc_hd__nand2_1 _20216_ (.A(_09742_),
    .B(_10000_),
    .Y(_10001_));
 sky130_fd_sc_hd__or2_1 _20217_ (.A(_09817_),
    .B(_09807_),
    .X(_10002_));
 sky130_fd_sc_hd__nand2_1 _20218_ (.A(_10002_),
    .B(_09818_),
    .Y(_10003_));
 sky130_fd_sc_hd__clkinvlp_2 _20219_ (.A(_10003_),
    .Y(_10004_));
 sky130_fd_sc_hd__nand3_1 _20220_ (.A(_09740_),
    .B(_09741_),
    .C(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__nand2_1 _20221_ (.A(_10001_),
    .B(_10005_),
    .Y(_10006_));
 sky130_fd_sc_hd__nand2_1 _20222_ (.A(_10006_),
    .B(_06033_),
    .Y(_10007_));
 sky130_fd_sc_hd__nand3_1 _20223_ (.A(_10001_),
    .B(_07092_),
    .C(_10005_),
    .Y(_10008_));
 sky130_fd_sc_hd__nand2_1 _20224_ (.A(_10007_),
    .B(_10008_),
    .Y(_10010_));
 sky130_fd_sc_hd__clkinvlp_2 _20225_ (.A(_10010_),
    .Y(_10011_));
 sky130_fd_sc_hd__nand2_1 _20226_ (.A(_09742_),
    .B(_09805_),
    .Y(_10012_));
 sky130_fd_sc_hd__nand2_1 _20227_ (.A(_09806_),
    .B(_09803_),
    .Y(_10013_));
 sky130_fd_sc_hd__xnor2_1 _20228_ (.A(_09798_),
    .B(_10013_),
    .Y(_10014_));
 sky130_fd_sc_hd__nand3_1 _20229_ (.A(_09740_),
    .B(_09741_),
    .C(_10014_),
    .Y(_10015_));
 sky130_fd_sc_hd__nand2_1 _20230_ (.A(_10012_),
    .B(_10015_),
    .Y(_10016_));
 sky130_fd_sc_hd__nand2_1 _20231_ (.A(_10016_),
    .B(_07102_),
    .Y(_10017_));
 sky130_fd_sc_hd__nand3_1 _20232_ (.A(_10012_),
    .B(_06046_),
    .C(_10015_),
    .Y(_10018_));
 sky130_fd_sc_hd__nand2_1 _20233_ (.A(_10017_),
    .B(_10018_),
    .Y(_10019_));
 sky130_fd_sc_hd__inv_2 _20234_ (.A(_10019_),
    .Y(_10021_));
 sky130_fd_sc_hd__nand2_1 _20235_ (.A(_10011_),
    .B(_10021_),
    .Y(_10022_));
 sky130_fd_sc_hd__nor2_1 _20236_ (.A(_09999_),
    .B(_10022_),
    .Y(_10023_));
 sky130_fd_sc_hd__nand2_1 _20237_ (.A(_09974_),
    .B(_10023_),
    .Y(_10024_));
 sky130_fd_sc_hd__inv_2 _20238_ (.A(_10008_),
    .Y(_10025_));
 sky130_fd_sc_hd__o21ai_2 _20239_ (.A1(_10017_),
    .A2(_10025_),
    .B1(_10007_),
    .Y(_10026_));
 sky130_fd_sc_hd__nor2_1 _20240_ (.A(_09986_),
    .B(_09996_),
    .Y(_10027_));
 sky130_fd_sc_hd__clkinvlp_2 _20241_ (.A(_09985_),
    .Y(_10028_));
 sky130_fd_sc_hd__o21ai_1 _20242_ (.A1(_09995_),
    .A2(_10028_),
    .B1(_09984_),
    .Y(_10029_));
 sky130_fd_sc_hd__a21oi_1 _20243_ (.A1(_10026_),
    .A2(_10027_),
    .B1(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__nand2_2 _20244_ (.A(_10024_),
    .B(_10030_),
    .Y(_10032_));
 sky130_fd_sc_hd__nand2_1 _20245_ (.A(_09852_),
    .B(_09858_),
    .Y(_10033_));
 sky130_fd_sc_hd__or2_1 _20246_ (.A(_09858_),
    .B(_09852_),
    .X(_10034_));
 sky130_fd_sc_hd__nand3_1 _20247_ (.A(_09904_),
    .B(_10033_),
    .C(_10034_),
    .Y(_10035_));
 sky130_fd_sc_hd__nand2_1 _20248_ (.A(_09742_),
    .B(_09774_),
    .Y(_10036_));
 sky130_fd_sc_hd__nand2_1 _20249_ (.A(_10035_),
    .B(_10036_),
    .Y(_10037_));
 sky130_fd_sc_hd__nand2_1 _20250_ (.A(_10037_),
    .B(_06695_),
    .Y(_10038_));
 sky130_fd_sc_hd__nand3_1 _20251_ (.A(_10035_),
    .B(_06697_),
    .C(_10036_),
    .Y(_10039_));
 sky130_fd_sc_hd__nand2_1 _20252_ (.A(_10038_),
    .B(_10039_),
    .Y(_10040_));
 sky130_fd_sc_hd__inv_2 _20253_ (.A(_10040_),
    .Y(_10041_));
 sky130_fd_sc_hd__nand2_1 _20254_ (.A(_09838_),
    .B(_09846_),
    .Y(_10043_));
 sky130_fd_sc_hd__nand2_1 _20255_ (.A(_09978_),
    .B(_09842_),
    .Y(_10044_));
 sky130_fd_sc_hd__xor2_1 _20256_ (.A(_10043_),
    .B(_10044_),
    .X(_10045_));
 sky130_fd_sc_hd__nand2_1 _20257_ (.A(_10045_),
    .B(_09904_),
    .Y(_10046_));
 sky130_fd_sc_hd__nand2_1 _20258_ (.A(_09743_),
    .B(_09837_),
    .Y(_10047_));
 sky130_fd_sc_hd__nand2_1 _20259_ (.A(_10046_),
    .B(_10047_),
    .Y(_10048_));
 sky130_fd_sc_hd__nand2_1 _20260_ (.A(_10048_),
    .B(_09410_),
    .Y(_10049_));
 sky130_fd_sc_hd__nand3_1 _20261_ (.A(_10046_),
    .B(_08951_),
    .C(_10047_),
    .Y(_10050_));
 sky130_fd_sc_hd__nand2_1 _20262_ (.A(_10049_),
    .B(_10050_),
    .Y(_10051_));
 sky130_fd_sc_hd__inv_2 _20263_ (.A(_10051_),
    .Y(_10052_));
 sky130_fd_sc_hd__nand2_1 _20264_ (.A(_10041_),
    .B(_10052_),
    .Y(_10054_));
 sky130_fd_sc_hd__nand2_1 _20265_ (.A(_10033_),
    .B(_09775_),
    .Y(_10055_));
 sky130_fd_sc_hd__nand2_1 _20266_ (.A(_10055_),
    .B(_09854_),
    .Y(_10056_));
 sky130_fd_sc_hd__nand3_1 _20267_ (.A(_10033_),
    .B(_09853_),
    .C(_09775_),
    .Y(_10057_));
 sky130_fd_sc_hd__nand2_1 _20268_ (.A(_10056_),
    .B(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__nand2_1 _20269_ (.A(_10058_),
    .B(_09904_),
    .Y(_10059_));
 sky130_fd_sc_hd__nand2_1 _20270_ (.A(_09743_),
    .B(_09770_),
    .Y(_10060_));
 sky130_fd_sc_hd__nand2_1 _20271_ (.A(_10059_),
    .B(_10060_),
    .Y(_10061_));
 sky130_fd_sc_hd__nand2_1 _20272_ (.A(_10061_),
    .B(_06721_),
    .Y(_10062_));
 sky130_fd_sc_hd__nand3_2 _20273_ (.A(_10059_),
    .B(_06723_),
    .C(_10060_),
    .Y(_10063_));
 sky130_fd_sc_hd__nand2_1 _20274_ (.A(_10062_),
    .B(_10063_),
    .Y(_10065_));
 sky130_fd_sc_hd__or2_1 _20275_ (.A(_09782_),
    .B(_09904_),
    .X(_10066_));
 sky130_fd_sc_hd__nand3_1 _20276_ (.A(_09926_),
    .B(_09784_),
    .C(_09781_),
    .Y(_10067_));
 sky130_fd_sc_hd__nand3_1 _20277_ (.A(_09928_),
    .B(_09904_),
    .C(_10067_),
    .Y(_10068_));
 sky130_fd_sc_hd__nand2_1 _20278_ (.A(_10066_),
    .B(_10068_),
    .Y(_10069_));
 sky130_fd_sc_hd__nand2_1 _20279_ (.A(_10069_),
    .B(_06731_),
    .Y(_10070_));
 sky130_fd_sc_hd__nand3_1 _20280_ (.A(_10066_),
    .B(_10068_),
    .C(_06733_),
    .Y(_10071_));
 sky130_fd_sc_hd__nand2_2 _20281_ (.A(_10070_),
    .B(_10071_),
    .Y(_10072_));
 sky130_fd_sc_hd__nor2_1 _20282_ (.A(_10065_),
    .B(_10072_),
    .Y(_10073_));
 sky130_fd_sc_hd__nor2b_1 _20283_ (.A(_10073_),
    .B_N(_10054_),
    .Y(_10074_));
 sky130_fd_sc_hd__nand2_1 _20284_ (.A(_10032_),
    .B(_10074_),
    .Y(_10076_));
 sky130_fd_sc_hd__inv_2 _20285_ (.A(_10039_),
    .Y(_10077_));
 sky130_fd_sc_hd__o21ai_2 _20286_ (.A1(_10050_),
    .A2(_10077_),
    .B1(_10038_),
    .Y(_10078_));
 sky130_fd_sc_hd__inv_2 _20287_ (.A(_10071_),
    .Y(_10079_));
 sky130_fd_sc_hd__o21ai_1 _20288_ (.A1(_10063_),
    .A2(_10079_),
    .B1(_10070_),
    .Y(_10080_));
 sky130_fd_sc_hd__a21oi_1 _20289_ (.A1(_10073_),
    .A2(_10078_),
    .B1(_10080_),
    .Y(_10081_));
 sky130_fd_sc_hd__nand2_2 _20290_ (.A(_10076_),
    .B(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__nand2_1 _20291_ (.A(_09935_),
    .B(_09936_),
    .Y(_10083_));
 sky130_fd_sc_hd__nand2_1 _20292_ (.A(_10083_),
    .B(_06159_),
    .Y(_10084_));
 sky130_fd_sc_hd__nand2_1 _20293_ (.A(_10084_),
    .B(_09937_),
    .Y(_10085_));
 sky130_fd_sc_hd__nand2_1 _20294_ (.A(_09945_),
    .B(_09941_),
    .Y(_10087_));
 sky130_fd_sc_hd__nor2_1 _20295_ (.A(_10085_),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__nand3_1 _20296_ (.A(_10082_),
    .B(_09925_),
    .C(_10088_),
    .Y(_10089_));
 sky130_fd_sc_hd__nand2_2 _20297_ (.A(_09949_),
    .B(_10089_),
    .Y(_10090_));
 sky130_fd_sc_hd__nand2_1 _20298_ (.A(_09619_),
    .B(_09620_),
    .Y(_10091_));
 sky130_fd_sc_hd__inv_4 _20299_ (.A(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__or2_1 _20300_ (.A(_10092_),
    .B(_09533_),
    .X(_10093_));
 sky130_fd_sc_hd__nand2_1 _20301_ (.A(_09533_),
    .B(_10092_),
    .Y(_10094_));
 sky130_fd_sc_hd__nand2_1 _20302_ (.A(_10093_),
    .B(_10094_),
    .Y(_10095_));
 sky130_fd_sc_hd__inv_2 _20303_ (.A(_10095_),
    .Y(_10096_));
 sky130_fd_sc_hd__nand2_1 _20304_ (.A(_10096_),
    .B(_06207_),
    .Y(_10098_));
 sky130_fd_sc_hd__nand2_1 _20305_ (.A(_10095_),
    .B(_08465_),
    .Y(_10099_));
 sky130_fd_sc_hd__nand2_1 _20306_ (.A(_10098_),
    .B(_10099_),
    .Y(_10100_));
 sky130_fd_sc_hd__inv_2 _20307_ (.A(_10100_),
    .Y(_10101_));
 sky130_fd_sc_hd__nand2_1 _20308_ (.A(_09894_),
    .B(_09505_),
    .Y(_10102_));
 sky130_fd_sc_hd__inv_2 _20309_ (.A(_09494_),
    .Y(_10103_));
 sky130_fd_sc_hd__nand2_1 _20310_ (.A(_10102_),
    .B(_10103_),
    .Y(_10104_));
 sky130_fd_sc_hd__nand3_1 _20311_ (.A(_09894_),
    .B(_09505_),
    .C(_09494_),
    .Y(_10105_));
 sky130_fd_sc_hd__nand2_1 _20312_ (.A(_10104_),
    .B(_10105_),
    .Y(_10106_));
 sky130_fd_sc_hd__nand2_1 _20313_ (.A(_10106_),
    .B(_07905_),
    .Y(_10107_));
 sky130_fd_sc_hd__nand3_1 _20314_ (.A(_10104_),
    .B(_06772_),
    .C(_10105_),
    .Y(_10109_));
 sky130_fd_sc_hd__nand3_1 _20315_ (.A(_09902_),
    .B(_10107_),
    .C(_10109_),
    .Y(_10110_));
 sky130_fd_sc_hd__inv_2 _20316_ (.A(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__nand3_1 _20317_ (.A(_09862_),
    .B(_09884_),
    .C(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__inv_2 _20318_ (.A(_10107_),
    .Y(_10113_));
 sky130_fd_sc_hd__o21ai_1 _20319_ (.A1(_09898_),
    .A2(_10113_),
    .B1(_10109_),
    .Y(_10114_));
 sky130_fd_sc_hd__nor2_1 _20320_ (.A(_09887_),
    .B(_10110_),
    .Y(_10115_));
 sky130_fd_sc_hd__nor2_1 _20321_ (.A(_10114_),
    .B(_10115_),
    .Y(_10116_));
 sky130_fd_sc_hd__nand2_2 _20322_ (.A(_10112_),
    .B(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__or2_1 _20323_ (.A(_10101_),
    .B(_10117_),
    .X(_10118_));
 sky130_fd_sc_hd__buf_6 _20324_ (.A(_09904_),
    .X(_10120_));
 sky130_fd_sc_hd__nand2_1 _20325_ (.A(_10117_),
    .B(_10101_),
    .Y(_10121_));
 sky130_fd_sc_hd__nand3_1 _20326_ (.A(_10118_),
    .B(_10120_),
    .C(_10121_),
    .Y(_10122_));
 sky130_fd_sc_hd__nand2_1 _20327_ (.A(\div1i.quot[12] ),
    .B(_10096_),
    .Y(_10123_));
 sky130_fd_sc_hd__nand2_1 _20328_ (.A(_10122_),
    .B(_10123_),
    .Y(_10124_));
 sky130_fd_sc_hd__xor2_2 _20329_ (.A(_06754_),
    .B(_10124_),
    .X(_10125_));
 sky130_fd_sc_hd__nand2_1 _20330_ (.A(_10107_),
    .B(_10109_),
    .Y(_10126_));
 sky130_fd_sc_hd__nand2_1 _20331_ (.A(_09903_),
    .B(_09898_),
    .Y(_10127_));
 sky130_fd_sc_hd__xor2_1 _20332_ (.A(_10126_),
    .B(_10127_),
    .X(_10128_));
 sky130_fd_sc_hd__nand2_1 _20333_ (.A(_10128_),
    .B(_10120_),
    .Y(_10129_));
 sky130_fd_sc_hd__nand2_1 _20334_ (.A(\div1i.quot[12] ),
    .B(_10106_),
    .Y(_10131_));
 sky130_fd_sc_hd__nand2_1 _20335_ (.A(_10129_),
    .B(_10131_),
    .Y(_10132_));
 sky130_fd_sc_hd__nand2_1 _20336_ (.A(_10132_),
    .B(_06797_),
    .Y(_10133_));
 sky130_fd_sc_hd__nand3_1 _20337_ (.A(_10129_),
    .B(_06799_),
    .C(_10131_),
    .Y(_10134_));
 sky130_fd_sc_hd__nand2_1 _20338_ (.A(_10133_),
    .B(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__nor2_1 _20339_ (.A(_10125_),
    .B(_10135_),
    .Y(_10136_));
 sky130_fd_sc_hd__nand2_1 _20340_ (.A(_10090_),
    .B(_10136_),
    .Y(_10137_));
 sky130_fd_sc_hd__buf_6 _20341_ (.A(_06805_),
    .X(_10138_));
 sky130_fd_sc_hd__nand2_1 _20342_ (.A(_10124_),
    .B(_10138_),
    .Y(_10139_));
 sky130_fd_sc_hd__o21a_1 _20343_ (.A1(_10134_),
    .A2(_10125_),
    .B1(_10139_),
    .X(_10140_));
 sky130_fd_sc_hd__nand2_1 _20344_ (.A(_10137_),
    .B(_10140_),
    .Y(_10142_));
 sky130_fd_sc_hd__nand2_1 _20345_ (.A(_09533_),
    .B(_09622_),
    .Y(_10143_));
 sky130_fd_sc_hd__inv_2 _20346_ (.A(_09626_),
    .Y(_10144_));
 sky130_fd_sc_hd__a21o_1 _20347_ (.A1(_10143_),
    .A2(_10144_),
    .B1(_09604_),
    .X(_10145_));
 sky130_fd_sc_hd__nand3_1 _20348_ (.A(_10143_),
    .B(_09604_),
    .C(_10144_),
    .Y(_10146_));
 sky130_fd_sc_hd__nand2_1 _20349_ (.A(_10145_),
    .B(_10146_),
    .Y(_10147_));
 sky130_fd_sc_hd__inv_2 _20350_ (.A(_10147_),
    .Y(_10148_));
 sky130_fd_sc_hd__nand2_1 _20351_ (.A(_10148_),
    .B(_06819_),
    .Y(_10149_));
 sky130_fd_sc_hd__nand2_1 _20352_ (.A(_10147_),
    .B(_07948_),
    .Y(_10150_));
 sky130_fd_sc_hd__nand2_1 _20353_ (.A(_10149_),
    .B(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__inv_4 _20354_ (.A(_10151_),
    .Y(_10153_));
 sky130_fd_sc_hd__nand2_1 _20355_ (.A(_10094_),
    .B(_09620_),
    .Y(_10154_));
 sky130_fd_sc_hd__xor2_2 _20356_ (.A(_09612_),
    .B(_10154_),
    .X(_10155_));
 sky130_fd_sc_hd__inv_2 _20357_ (.A(_10155_),
    .Y(_10156_));
 sky130_fd_sc_hd__nand2_1 _20358_ (.A(_10156_),
    .B(_06827_),
    .Y(_10157_));
 sky130_fd_sc_hd__nand2_1 _20359_ (.A(_10155_),
    .B(_07957_),
    .Y(_10158_));
 sky130_fd_sc_hd__nand2_1 _20360_ (.A(_10157_),
    .B(_10158_),
    .Y(_10159_));
 sky130_fd_sc_hd__or2_1 _20361_ (.A(_10100_),
    .B(_10159_),
    .X(_10160_));
 sky130_fd_sc_hd__inv_4 _20362_ (.A(_10160_),
    .Y(_10161_));
 sky130_fd_sc_hd__nand2_1 _20363_ (.A(_10117_),
    .B(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__inv_2 _20364_ (.A(_10098_),
    .Y(_10164_));
 sky130_fd_sc_hd__a21boi_1 _20365_ (.A1(_10164_),
    .A2(_10158_),
    .B1_N(_10157_),
    .Y(_10165_));
 sky130_fd_sc_hd__nand2_1 _20366_ (.A(_10162_),
    .B(_10165_),
    .Y(_10166_));
 sky130_fd_sc_hd__or2_1 _20367_ (.A(_10153_),
    .B(_10166_),
    .X(_10167_));
 sky130_fd_sc_hd__nand2_1 _20368_ (.A(_10166_),
    .B(_10153_),
    .Y(_10168_));
 sky130_fd_sc_hd__nand3_1 _20369_ (.A(_10167_),
    .B(_10120_),
    .C(_10168_),
    .Y(_10169_));
 sky130_fd_sc_hd__nand2_1 _20370_ (.A(\div1i.quot[12] ),
    .B(_10148_),
    .Y(_10170_));
 sky130_fd_sc_hd__nand2_1 _20371_ (.A(_10169_),
    .B(_10170_),
    .Y(_10171_));
 sky130_fd_sc_hd__xor2_2 _20372_ (.A(_06809_),
    .B(_10171_),
    .X(_10172_));
 sky130_fd_sc_hd__buf_6 _20373_ (.A(_06844_),
    .X(_10173_));
 sky130_fd_sc_hd__nand2_1 _20374_ (.A(_10121_),
    .B(_10098_),
    .Y(_10175_));
 sky130_fd_sc_hd__xor2_1 _20375_ (.A(_10159_),
    .B(_10175_),
    .X(_10176_));
 sky130_fd_sc_hd__nand2_1 _20376_ (.A(_10176_),
    .B(_10120_),
    .Y(_10177_));
 sky130_fd_sc_hd__nand2_1 _20377_ (.A(\div1i.quot[12] ),
    .B(_10155_),
    .Y(_10178_));
 sky130_fd_sc_hd__nand2_1 _20378_ (.A(_10177_),
    .B(_10178_),
    .Y(_10179_));
 sky130_fd_sc_hd__or2_1 _20379_ (.A(_10173_),
    .B(_10179_),
    .X(_10180_));
 sky130_fd_sc_hd__nand2_1 _20380_ (.A(_10179_),
    .B(_10173_),
    .Y(_10181_));
 sky130_fd_sc_hd__nand2_1 _20381_ (.A(_10180_),
    .B(_10181_),
    .Y(_10182_));
 sky130_fd_sc_hd__nor2_1 _20382_ (.A(_10172_),
    .B(_10182_),
    .Y(_10183_));
 sky130_fd_sc_hd__nand2_1 _20383_ (.A(_10142_),
    .B(_10183_),
    .Y(_10184_));
 sky130_fd_sc_hd__nand2_1 _20384_ (.A(_10171_),
    .B(_06856_),
    .Y(_10186_));
 sky130_fd_sc_hd__o21a_1 _20385_ (.A1(_10180_),
    .A2(_10172_),
    .B1(_10186_),
    .X(_10187_));
 sky130_fd_sc_hd__nand2_2 _20386_ (.A(_10184_),
    .B(_10187_),
    .Y(_10188_));
 sky130_fd_sc_hd__nand2_1 _20387_ (.A(_09675_),
    .B(_09676_),
    .Y(_10189_));
 sky130_fd_sc_hd__nand2b_1 _20388_ (.A_N(_09629_),
    .B(_10189_),
    .Y(_10190_));
 sky130_fd_sc_hd__nand2b_1 _20389_ (.A_N(_10189_),
    .B(_09629_),
    .Y(_10191_));
 sky130_fd_sc_hd__nand2_1 _20390_ (.A(_10190_),
    .B(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__or2_1 _20391_ (.A(_07450_),
    .B(_10192_),
    .X(_10193_));
 sky130_fd_sc_hd__nand2_1 _20392_ (.A(_10192_),
    .B(_07450_),
    .Y(_10194_));
 sky130_fd_sc_hd__nand2_1 _20393_ (.A(_10193_),
    .B(_10194_),
    .Y(_10195_));
 sky130_fd_sc_hd__inv_4 _20394_ (.A(_10195_),
    .Y(_10197_));
 sky130_fd_sc_hd__nand2_1 _20395_ (.A(_10145_),
    .B(_09602_),
    .Y(_10198_));
 sky130_fd_sc_hd__inv_2 _20396_ (.A(_09594_),
    .Y(_10199_));
 sky130_fd_sc_hd__nand2_1 _20397_ (.A(_10198_),
    .B(_10199_),
    .Y(_10200_));
 sky130_fd_sc_hd__nand3_1 _20398_ (.A(_10145_),
    .B(_09594_),
    .C(_09602_),
    .Y(_10201_));
 sky130_fd_sc_hd__nand2_1 _20399_ (.A(_10200_),
    .B(_10201_),
    .Y(_10202_));
 sky130_fd_sc_hd__nand2_1 _20400_ (.A(_10202_),
    .B(_08001_),
    .Y(_10203_));
 sky130_fd_sc_hd__nand3_1 _20401_ (.A(_10200_),
    .B(_06874_),
    .C(_10201_),
    .Y(_10204_));
 sky130_fd_sc_hd__nand3_1 _20402_ (.A(_10153_),
    .B(_10203_),
    .C(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__inv_2 _20403_ (.A(_10205_),
    .Y(_10206_));
 sky130_fd_sc_hd__nand3_1 _20404_ (.A(_10117_),
    .B(_10161_),
    .C(_10206_),
    .Y(_10208_));
 sky130_fd_sc_hd__inv_2 _20405_ (.A(_10149_),
    .Y(_10209_));
 sky130_fd_sc_hd__inv_2 _20406_ (.A(_10204_),
    .Y(_10210_));
 sky130_fd_sc_hd__a21o_1 _20407_ (.A1(_10203_),
    .A2(_10209_),
    .B1(_10210_),
    .X(_10211_));
 sky130_fd_sc_hd__nor2_1 _20408_ (.A(_10165_),
    .B(_10205_),
    .Y(_10212_));
 sky130_fd_sc_hd__nor2_1 _20409_ (.A(_10211_),
    .B(_10212_),
    .Y(_10213_));
 sky130_fd_sc_hd__nand2_1 _20410_ (.A(_10208_),
    .B(_10213_),
    .Y(_10214_));
 sky130_fd_sc_hd__or2_1 _20411_ (.A(_10197_),
    .B(_10214_),
    .X(_10215_));
 sky130_fd_sc_hd__nand2_1 _20412_ (.A(_10214_),
    .B(_10197_),
    .Y(_10216_));
 sky130_fd_sc_hd__nand2_1 _20413_ (.A(_10215_),
    .B(_10216_),
    .Y(_10217_));
 sky130_fd_sc_hd__nand2_1 _20414_ (.A(_10217_),
    .B(_10120_),
    .Y(_10219_));
 sky130_fd_sc_hd__nand2_1 _20415_ (.A(\div1i.quot[12] ),
    .B(_10192_),
    .Y(_10220_));
 sky130_fd_sc_hd__nand2_1 _20416_ (.A(_10219_),
    .B(_10220_),
    .Y(_10221_));
 sky130_fd_sc_hd__nand2_1 _20417_ (.A(_10221_),
    .B(_08020_),
    .Y(_10222_));
 sky130_fd_sc_hd__nand3_1 _20418_ (.A(_10219_),
    .B(_09664_),
    .C(_10220_),
    .Y(_10223_));
 sky130_fd_sc_hd__nand2_2 _20419_ (.A(_10222_),
    .B(_10223_),
    .Y(_10224_));
 sky130_fd_sc_hd__inv_2 _20420_ (.A(_10224_),
    .Y(_10225_));
 sky130_fd_sc_hd__nand2_1 _20421_ (.A(_10203_),
    .B(_10204_),
    .Y(_10226_));
 sky130_fd_sc_hd__nand2_1 _20422_ (.A(_10168_),
    .B(_10149_),
    .Y(_10227_));
 sky130_fd_sc_hd__xor2_1 _20423_ (.A(_10226_),
    .B(_10227_),
    .X(_10228_));
 sky130_fd_sc_hd__nand2_1 _20424_ (.A(_10228_),
    .B(_10120_),
    .Y(_10230_));
 sky130_fd_sc_hd__nand2_1 _20425_ (.A(_10202_),
    .B(\div1i.quot[12] ),
    .Y(_10231_));
 sky130_fd_sc_hd__nand2_1 _20426_ (.A(_10230_),
    .B(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__nand2_1 _20427_ (.A(_10232_),
    .B(_06903_),
    .Y(_10233_));
 sky130_fd_sc_hd__nand3_2 _20428_ (.A(_10230_),
    .B(_06898_),
    .C(_10231_),
    .Y(_10234_));
 sky130_fd_sc_hd__nand3_1 _20429_ (.A(_10225_),
    .B(_10233_),
    .C(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__nand2_1 _20430_ (.A(_10216_),
    .B(_10193_),
    .Y(_10236_));
 sky130_fd_sc_hd__nand2_1 _20431_ (.A(_10191_),
    .B(_09676_),
    .Y(_10237_));
 sky130_fd_sc_hd__or2_1 _20432_ (.A(_09667_),
    .B(_10237_),
    .X(_10238_));
 sky130_fd_sc_hd__nand2_1 _20433_ (.A(_10237_),
    .B(_09667_),
    .Y(_10239_));
 sky130_fd_sc_hd__nand2_1 _20434_ (.A(_10238_),
    .B(_10239_),
    .Y(_10241_));
 sky130_fd_sc_hd__nand2_1 _20435_ (.A(_10241_),
    .B(_08041_),
    .Y(_10242_));
 sky130_fd_sc_hd__nand3_1 _20436_ (.A(_10238_),
    .B(_07461_),
    .C(_10239_),
    .Y(_10243_));
 sky130_fd_sc_hd__nand2_1 _20437_ (.A(_10242_),
    .B(_10243_),
    .Y(_10244_));
 sky130_fd_sc_hd__inv_2 _20438_ (.A(_10244_),
    .Y(_10245_));
 sky130_fd_sc_hd__nand2_1 _20439_ (.A(_10236_),
    .B(_10245_),
    .Y(_10246_));
 sky130_fd_sc_hd__nand3_1 _20440_ (.A(_10216_),
    .B(_10244_),
    .C(_10193_),
    .Y(_10247_));
 sky130_fd_sc_hd__nand2_1 _20441_ (.A(_10246_),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__nand2_1 _20442_ (.A(_10248_),
    .B(_10120_),
    .Y(_10249_));
 sky130_fd_sc_hd__nand2_1 _20443_ (.A(_10241_),
    .B(\div1i.quot[12] ),
    .Y(_10250_));
 sky130_fd_sc_hd__nand2_1 _20444_ (.A(_10249_),
    .B(_10250_),
    .Y(_10252_));
 sky130_fd_sc_hd__nand2_1 _20445_ (.A(_10252_),
    .B(_07474_),
    .Y(_10253_));
 sky130_fd_sc_hd__nand3_1 _20446_ (.A(_10249_),
    .B(_06366_),
    .C(_10250_),
    .Y(_10254_));
 sky130_fd_sc_hd__nand2_1 _20447_ (.A(_10253_),
    .B(_10254_),
    .Y(_10255_));
 sky130_fd_sc_hd__inv_2 _20448_ (.A(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__nand2_1 _20449_ (.A(_10245_),
    .B(_10197_),
    .Y(_10257_));
 sky130_fd_sc_hd__inv_2 _20450_ (.A(_10257_),
    .Y(_10258_));
 sky130_fd_sc_hd__nand2_1 _20451_ (.A(_10214_),
    .B(_10258_),
    .Y(_10259_));
 sky130_fd_sc_hd__o21a_1 _20452_ (.A1(_10193_),
    .A2(_10244_),
    .B1(_10243_),
    .X(_10260_));
 sky130_fd_sc_hd__nand2_1 _20453_ (.A(_10259_),
    .B(_10260_),
    .Y(_10261_));
 sky130_fd_sc_hd__a41o_1 _20454_ (.A1(_09629_),
    .A2(_09667_),
    .A3(_09676_),
    .A4(_09675_),
    .B1(_09728_),
    .X(_10263_));
 sky130_fd_sc_hd__or2_1 _20455_ (.A(_09697_),
    .B(_10263_),
    .X(_10264_));
 sky130_fd_sc_hd__nand2_1 _20456_ (.A(_10263_),
    .B(_09697_),
    .Y(_10265_));
 sky130_fd_sc_hd__nand2_1 _20457_ (.A(_10264_),
    .B(_10265_),
    .Y(_10266_));
 sky130_fd_sc_hd__inv_2 _20458_ (.A(_10266_),
    .Y(_10267_));
 sky130_fd_sc_hd__nand2_1 _20459_ (.A(_10267_),
    .B(_06936_),
    .Y(_10268_));
 sky130_fd_sc_hd__nand2_1 _20460_ (.A(_10266_),
    .B(_08611_),
    .Y(_10269_));
 sky130_fd_sc_hd__nand2_1 _20461_ (.A(_10268_),
    .B(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__inv_2 _20462_ (.A(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__nand2_1 _20463_ (.A(_10261_),
    .B(_10271_),
    .Y(_10272_));
 sky130_fd_sc_hd__nand3_1 _20464_ (.A(_10259_),
    .B(_10270_),
    .C(_10260_),
    .Y(_10274_));
 sky130_fd_sc_hd__nand3_1 _20465_ (.A(_10272_),
    .B(_10274_),
    .C(_10120_),
    .Y(_10275_));
 sky130_fd_sc_hd__nand2_1 _20466_ (.A(_10267_),
    .B(\div1i.quot[12] ),
    .Y(_10276_));
 sky130_fd_sc_hd__nand2_1 _20467_ (.A(_10275_),
    .B(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__nand2_1 _20468_ (.A(_10277_),
    .B(_06947_),
    .Y(_10278_));
 sky130_fd_sc_hd__nand3_1 _20469_ (.A(_10275_),
    .B(_06949_),
    .C(_10276_),
    .Y(_10279_));
 sky130_fd_sc_hd__nand2_4 _20470_ (.A(_10279_),
    .B(_10278_),
    .Y(_10280_));
 sky130_fd_sc_hd__inv_2 _20471_ (.A(_10280_),
    .Y(_10281_));
 sky130_fd_sc_hd__nand2_1 _20472_ (.A(_10256_),
    .B(_10281_),
    .Y(_10282_));
 sky130_fd_sc_hd__nor2_2 _20473_ (.A(_10235_),
    .B(_10282_),
    .Y(_10283_));
 sky130_fd_sc_hd__nand2_4 _20474_ (.A(_10188_),
    .B(_10283_),
    .Y(_10285_));
 sky130_fd_sc_hd__o21ai_1 _20475_ (.A1(_10234_),
    .A2(_10224_),
    .B1(_10223_),
    .Y(_10286_));
 sky130_fd_sc_hd__nor2_1 _20476_ (.A(_10280_),
    .B(_10255_),
    .Y(_10287_));
 sky130_fd_sc_hd__o21ai_1 _20477_ (.A1(_10254_),
    .A2(_10280_),
    .B1(_10278_),
    .Y(_10288_));
 sky130_fd_sc_hd__a21oi_2 _20478_ (.A1(_10286_),
    .A2(_10287_),
    .B1(_10288_),
    .Y(_10289_));
 sky130_fd_sc_hd__nand2_2 _20479_ (.A(_10285_),
    .B(_10289_),
    .Y(_10290_));
 sky130_fd_sc_hd__nand2_2 _20480_ (.A(_10265_),
    .B(_09695_),
    .Y(_10291_));
 sky130_fd_sc_hd__xor2_4 _20481_ (.A(_09722_),
    .B(_10291_),
    .X(_10292_));
 sky130_fd_sc_hd__nand3_2 _20482_ (.A(_10272_),
    .B(_10120_),
    .C(_10268_),
    .Y(_10293_));
 sky130_fd_sc_hd__xnor2_4 _20483_ (.A(_10292_),
    .B(_10293_),
    .Y(_10294_));
 sky130_fd_sc_hd__nand2_8 _20484_ (.A(_10290_),
    .B(_10294_),
    .Y(_10296_));
 sky130_fd_sc_hd__clkinvlp_2 _20485_ (.A(_10294_),
    .Y(_10297_));
 sky130_fd_sc_hd__nand3_4 _20486_ (.A(_10285_),
    .B(_10289_),
    .C(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__nand2_8 _20487_ (.A(_10296_),
    .B(_10298_),
    .Y(_10299_));
 sky130_fd_sc_hd__buf_8 _20488_ (.A(_10299_),
    .X(_10300_));
 sky130_fd_sc_hd__buf_8 _20489_ (.A(net225),
    .X(\div1i.quot[11] ));
 sky130_fd_sc_hd__nand2_1 _20490_ (.A(_09966_),
    .B(_09969_),
    .Y(_10301_));
 sky130_fd_sc_hd__nand2_1 _20491_ (.A(_10301_),
    .B(_09970_),
    .Y(_10302_));
 sky130_fd_sc_hd__nand2_1 _20492_ (.A(_10302_),
    .B(_09972_),
    .Y(_10303_));
 sky130_fd_sc_hd__inv_2 _20493_ (.A(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__nand2_1 _20494_ (.A(_10300_),
    .B(_10304_),
    .Y(_10306_));
 sky130_fd_sc_hd__o21ai_1 _20495_ (.A1(_09215_),
    .A2(\div1i.quot[12] ),
    .B1(_09228_),
    .Y(_10307_));
 sky130_fd_sc_hd__nand2_1 _20496_ (.A(_10303_),
    .B(_06982_),
    .Y(_10308_));
 sky130_fd_sc_hd__nand3_1 _20497_ (.A(_10302_),
    .B(_06984_),
    .C(_09972_),
    .Y(_10309_));
 sky130_fd_sc_hd__nand2_1 _20498_ (.A(_10308_),
    .B(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__xor2_1 _20499_ (.A(_10307_),
    .B(_10310_),
    .X(_10311_));
 sky130_fd_sc_hd__nand3b_1 _20500_ (.A_N(_10311_),
    .B(_10296_),
    .C(_10298_),
    .Y(_10312_));
 sky130_fd_sc_hd__nand2_1 _20501_ (.A(_10306_),
    .B(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__nand2_1 _20502_ (.A(_10313_),
    .B(_08857_),
    .Y(_10314_));
 sky130_fd_sc_hd__nor2_1 _20503_ (.A(_09215_),
    .B(_10120_),
    .Y(_10315_));
 sky130_fd_sc_hd__or2_1 _20504_ (.A(_06607_),
    .B(_10315_),
    .X(_10317_));
 sky130_fd_sc_hd__nand2_1 _20505_ (.A(_10317_),
    .B(_09970_),
    .Y(_10318_));
 sky130_fd_sc_hd__inv_2 _20506_ (.A(_10318_),
    .Y(_10319_));
 sky130_fd_sc_hd__nand2_2 _20507_ (.A(_10300_),
    .B(_10319_),
    .Y(_10320_));
 sky130_fd_sc_hd__nand3_1 _20508_ (.A(_10296_),
    .B(_10298_),
    .C(_10315_),
    .Y(_10321_));
 sky130_fd_sc_hd__nand2_2 _20509_ (.A(_10320_),
    .B(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__nand2_4 _20510_ (.A(_10322_),
    .B(_06615_),
    .Y(_10323_));
 sky130_fd_sc_hd__nand2_2 _20511_ (.A(_10314_),
    .B(_10323_),
    .Y(_10324_));
 sky130_fd_sc_hd__inv_2 _20512_ (.A(_10324_),
    .Y(_10325_));
 sky130_fd_sc_hd__nand3_2 _20513_ (.A(_10320_),
    .B(_06620_),
    .C(_10321_),
    .Y(_10326_));
 sky130_fd_sc_hd__nand3_2 _20514_ (.A(_10300_),
    .B(_09228_),
    .C(_07004_),
    .Y(_10328_));
 sky130_fd_sc_hd__inv_2 _20515_ (.A(_10328_),
    .Y(_10329_));
 sky130_fd_sc_hd__nand3_4 _20516_ (.A(_10323_),
    .B(_10326_),
    .C(_10329_),
    .Y(_10330_));
 sky130_fd_sc_hd__or2_4 _20517_ (.A(_08857_),
    .B(_10313_),
    .X(_10331_));
 sky130_fd_sc_hd__inv_2 _20518_ (.A(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__a21oi_2 _20519_ (.A1(_10325_),
    .A2(_10330_),
    .B1(_10332_),
    .Y(_10333_));
 sky130_fd_sc_hd__nand2_1 _20520_ (.A(_09968_),
    .B(_09972_),
    .Y(_10334_));
 sky130_fd_sc_hd__nand2_1 _20521_ (.A(_10334_),
    .B(_09973_),
    .Y(_10335_));
 sky130_fd_sc_hd__inv_2 _20522_ (.A(_10026_),
    .Y(_10336_));
 sky130_fd_sc_hd__o21ai_1 _20523_ (.A1(_10022_),
    .A2(_10335_),
    .B1(_10336_),
    .Y(_10337_));
 sky130_fd_sc_hd__or2_1 _20524_ (.A(_09997_),
    .B(_10337_),
    .X(_10339_));
 sky130_fd_sc_hd__nand2_1 _20525_ (.A(_10337_),
    .B(_09997_),
    .Y(_10340_));
 sky130_fd_sc_hd__nand2_1 _20526_ (.A(_10339_),
    .B(_10340_),
    .Y(_10341_));
 sky130_fd_sc_hd__inv_2 _20527_ (.A(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__nand2_1 _20528_ (.A(_10299_),
    .B(_10342_),
    .Y(_10343_));
 sky130_fd_sc_hd__nand2_1 _20529_ (.A(_10342_),
    .B(_07021_),
    .Y(_10344_));
 sky130_fd_sc_hd__nand2_1 _20530_ (.A(_10341_),
    .B(_07024_),
    .Y(_10345_));
 sky130_fd_sc_hd__nand2_1 _20531_ (.A(_10344_),
    .B(_10345_),
    .Y(_10346_));
 sky130_fd_sc_hd__inv_2 _20532_ (.A(_10346_),
    .Y(_10347_));
 sky130_fd_sc_hd__nand2_1 _20533_ (.A(_09974_),
    .B(_10021_),
    .Y(_10348_));
 sky130_fd_sc_hd__nand2_1 _20534_ (.A(_10335_),
    .B(_10019_),
    .Y(_10350_));
 sky130_fd_sc_hd__nand2_1 _20535_ (.A(_10348_),
    .B(_10350_),
    .Y(_10351_));
 sky130_fd_sc_hd__nand2_1 _20536_ (.A(_10351_),
    .B(_07031_),
    .Y(_10352_));
 sky130_fd_sc_hd__nand3_1 _20537_ (.A(_10348_),
    .B(_07034_),
    .C(_10350_),
    .Y(_10353_));
 sky130_fd_sc_hd__nand2_1 _20538_ (.A(_10352_),
    .B(_10353_),
    .Y(_10354_));
 sky130_fd_sc_hd__inv_2 _20539_ (.A(_10354_),
    .Y(_10355_));
 sky130_fd_sc_hd__inv_2 _20540_ (.A(_10309_),
    .Y(_10356_));
 sky130_fd_sc_hd__a21o_1 _20541_ (.A1(_10308_),
    .A2(_10307_),
    .B1(_10356_),
    .X(_10357_));
 sky130_fd_sc_hd__nand2_1 _20542_ (.A(_09973_),
    .B(_09957_),
    .Y(_10358_));
 sky130_fd_sc_hd__nand2_1 _20543_ (.A(_09972_),
    .B(_09966_),
    .Y(_10359_));
 sky130_fd_sc_hd__xor2_1 _20544_ (.A(_10358_),
    .B(_10359_),
    .X(_10361_));
 sky130_fd_sc_hd__nand2_1 _20545_ (.A(_10361_),
    .B(_07043_),
    .Y(_10362_));
 sky130_fd_sc_hd__nand2_1 _20546_ (.A(_10357_),
    .B(_10362_),
    .Y(_10363_));
 sky130_fd_sc_hd__inv_2 _20547_ (.A(_10361_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand2_1 _20548_ (.A(_10364_),
    .B(_07048_),
    .Y(_10365_));
 sky130_fd_sc_hd__nand2_1 _20549_ (.A(_10363_),
    .B(_10365_),
    .Y(_10366_));
 sky130_fd_sc_hd__nand2_1 _20550_ (.A(_10355_),
    .B(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__nand2_1 _20551_ (.A(_10367_),
    .B(_10353_),
    .Y(_10368_));
 sky130_fd_sc_hd__nand2_1 _20552_ (.A(_10348_),
    .B(_10017_),
    .Y(_10369_));
 sky130_fd_sc_hd__xor2_1 _20553_ (.A(_10010_),
    .B(_10369_),
    .X(_10370_));
 sky130_fd_sc_hd__nand2_1 _20554_ (.A(_10370_),
    .B(_09823_),
    .Y(_10372_));
 sky130_fd_sc_hd__nand2_1 _20555_ (.A(_10368_),
    .B(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__inv_2 _20556_ (.A(_10370_),
    .Y(_10374_));
 sky130_fd_sc_hd__nand2_1 _20557_ (.A(_10374_),
    .B(_08176_),
    .Y(_10375_));
 sky130_fd_sc_hd__nand2_1 _20558_ (.A(_10373_),
    .B(_10375_),
    .Y(_10376_));
 sky130_fd_sc_hd__or2_1 _20559_ (.A(_10347_),
    .B(_10376_),
    .X(_10377_));
 sky130_fd_sc_hd__nand2_2 _20560_ (.A(_10376_),
    .B(_10347_),
    .Y(_10378_));
 sky130_fd_sc_hd__nand2_1 _20561_ (.A(_10377_),
    .B(_10378_),
    .Y(_10379_));
 sky130_fd_sc_hd__inv_2 _20562_ (.A(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__nand3_1 _20563_ (.A(_10296_),
    .B(_10298_),
    .C(_10380_),
    .Y(_10381_));
 sky130_fd_sc_hd__nand2_1 _20564_ (.A(_10343_),
    .B(_10381_),
    .Y(_10383_));
 sky130_fd_sc_hd__nand2_1 _20565_ (.A(_10383_),
    .B(_06636_),
    .Y(_10384_));
 sky130_fd_sc_hd__nand3_1 _20566_ (.A(_10343_),
    .B(_06639_),
    .C(_10381_),
    .Y(_10385_));
 sky130_fd_sc_hd__nand2_1 _20567_ (.A(_10384_),
    .B(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__inv_2 _20568_ (.A(_10386_),
    .Y(_10387_));
 sky130_fd_sc_hd__nand2_1 _20569_ (.A(_10299_),
    .B(_10374_),
    .Y(_10388_));
 sky130_fd_sc_hd__nand2_1 _20570_ (.A(_10375_),
    .B(_10372_),
    .Y(_10389_));
 sky130_fd_sc_hd__xnor2_1 _20571_ (.A(_10368_),
    .B(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__nand3_1 _20572_ (.A(_10296_),
    .B(_10298_),
    .C(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__nand2_1 _20573_ (.A(_10388_),
    .B(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__nand2_2 _20574_ (.A(_10392_),
    .B(_06651_),
    .Y(_10394_));
 sky130_fd_sc_hd__nand3_1 _20575_ (.A(_10388_),
    .B(_06648_),
    .C(_10391_),
    .Y(_10395_));
 sky130_fd_sc_hd__nand2_2 _20576_ (.A(_10394_),
    .B(_10395_),
    .Y(_10396_));
 sky130_fd_sc_hd__inv_2 _20577_ (.A(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__nand2_1 _20578_ (.A(_10387_),
    .B(_10397_),
    .Y(_10398_));
 sky130_fd_sc_hd__inv_2 _20579_ (.A(_10351_),
    .Y(_10399_));
 sky130_fd_sc_hd__nand2_1 _20580_ (.A(_10299_),
    .B(_10399_),
    .Y(_10400_));
 sky130_fd_sc_hd__or2_1 _20581_ (.A(_10366_),
    .B(_10355_),
    .X(_10401_));
 sky130_fd_sc_hd__nand2_1 _20582_ (.A(_10401_),
    .B(_10367_),
    .Y(_10402_));
 sky130_fd_sc_hd__clkinvlp_2 _20583_ (.A(_10402_),
    .Y(_10403_));
 sky130_fd_sc_hd__nand3_1 _20584_ (.A(_10296_),
    .B(_10298_),
    .C(_10403_),
    .Y(_10405_));
 sky130_fd_sc_hd__nand2_1 _20585_ (.A(_10400_),
    .B(_10405_),
    .Y(_10406_));
 sky130_fd_sc_hd__nand2_1 _20586_ (.A(_10406_),
    .B(_06033_),
    .Y(_10407_));
 sky130_fd_sc_hd__nand3_1 _20587_ (.A(_10400_),
    .B(_07092_),
    .C(_10405_),
    .Y(_10408_));
 sky130_fd_sc_hd__nand2_1 _20588_ (.A(_10407_),
    .B(_10408_),
    .Y(_10409_));
 sky130_fd_sc_hd__inv_2 _20589_ (.A(_10409_),
    .Y(_10410_));
 sky130_fd_sc_hd__nand2_1 _20590_ (.A(_10299_),
    .B(_10364_),
    .Y(_10411_));
 sky130_fd_sc_hd__nand2_1 _20591_ (.A(_10365_),
    .B(_10362_),
    .Y(_10412_));
 sky130_fd_sc_hd__xnor2_1 _20592_ (.A(_10357_),
    .B(_10412_),
    .Y(_10413_));
 sky130_fd_sc_hd__nand3_1 _20593_ (.A(_10296_),
    .B(_10298_),
    .C(_10413_),
    .Y(_10414_));
 sky130_fd_sc_hd__nand2_1 _20594_ (.A(_10411_),
    .B(_10414_),
    .Y(_10416_));
 sky130_fd_sc_hd__nand2_1 _20595_ (.A(_10416_),
    .B(_07102_),
    .Y(_10417_));
 sky130_fd_sc_hd__nand3_1 _20596_ (.A(_10411_),
    .B(_06046_),
    .C(_10414_),
    .Y(_10418_));
 sky130_fd_sc_hd__nand2_2 _20597_ (.A(_10417_),
    .B(_10418_),
    .Y(_10419_));
 sky130_fd_sc_hd__inv_2 _20598_ (.A(_10419_),
    .Y(_10420_));
 sky130_fd_sc_hd__nand2_1 _20599_ (.A(_10410_),
    .B(_10420_),
    .Y(_10421_));
 sky130_fd_sc_hd__nor2_1 _20600_ (.A(_10398_),
    .B(_10421_),
    .Y(_10422_));
 sky130_fd_sc_hd__nand2_1 _20601_ (.A(_10333_),
    .B(_10422_),
    .Y(_10423_));
 sky130_fd_sc_hd__inv_2 _20602_ (.A(_10408_),
    .Y(_10424_));
 sky130_fd_sc_hd__o21ai_2 _20603_ (.A1(_10417_),
    .A2(_10424_),
    .B1(_10407_),
    .Y(_10425_));
 sky130_fd_sc_hd__nor2_1 _20604_ (.A(_10386_),
    .B(_10396_),
    .Y(_10427_));
 sky130_fd_sc_hd__inv_2 _20605_ (.A(_10385_),
    .Y(_10428_));
 sky130_fd_sc_hd__o21ai_1 _20606_ (.A1(_10394_),
    .A2(_10428_),
    .B1(_10384_),
    .Y(_10429_));
 sky130_fd_sc_hd__a21oi_1 _20607_ (.A1(_10425_),
    .A2(_10427_),
    .B1(_10429_),
    .Y(_10430_));
 sky130_fd_sc_hd__nand2_2 _20608_ (.A(_10423_),
    .B(_10430_),
    .Y(_10431_));
 sky130_fd_sc_hd__inv_2 _20609_ (.A(_10054_),
    .Y(_10432_));
 sky130_fd_sc_hd__nand2_1 _20610_ (.A(_10032_),
    .B(_10432_),
    .Y(_10433_));
 sky130_fd_sc_hd__inv_2 _20611_ (.A(_10078_),
    .Y(_10434_));
 sky130_fd_sc_hd__nand2_1 _20612_ (.A(_10433_),
    .B(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__inv_2 _20613_ (.A(_10065_),
    .Y(_10436_));
 sky130_fd_sc_hd__nand2_1 _20614_ (.A(_10435_),
    .B(_10436_),
    .Y(_10438_));
 sky130_fd_sc_hd__nand3_1 _20615_ (.A(_10433_),
    .B(_10065_),
    .C(_10434_),
    .Y(_10439_));
 sky130_fd_sc_hd__nand2_1 _20616_ (.A(_10438_),
    .B(_10439_),
    .Y(_10440_));
 sky130_fd_sc_hd__inv_2 _20617_ (.A(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__nand2_1 _20618_ (.A(_10441_),
    .B(_07128_),
    .Y(_10442_));
 sky130_fd_sc_hd__nand2_1 _20619_ (.A(_10440_),
    .B(_07130_),
    .Y(_10443_));
 sky130_fd_sc_hd__nand2_1 _20620_ (.A(_10442_),
    .B(_10443_),
    .Y(_10444_));
 sky130_fd_sc_hd__inv_2 _20621_ (.A(_10444_),
    .Y(_10445_));
 sky130_fd_sc_hd__nand2_1 _20622_ (.A(_10340_),
    .B(_09995_),
    .Y(_10446_));
 sky130_fd_sc_hd__or2_1 _20623_ (.A(_09988_),
    .B(_10446_),
    .X(_10447_));
 sky130_fd_sc_hd__nand2_1 _20624_ (.A(_10446_),
    .B(_09988_),
    .Y(_10449_));
 sky130_fd_sc_hd__nand3_1 _20625_ (.A(_10447_),
    .B(_05896_),
    .C(_10449_),
    .Y(_10450_));
 sky130_fd_sc_hd__nand2_1 _20626_ (.A(_10450_),
    .B(_10344_),
    .Y(_10451_));
 sky130_fd_sc_hd__inv_2 _20627_ (.A(_10451_),
    .Y(_10452_));
 sky130_fd_sc_hd__nand2_2 _20628_ (.A(_10378_),
    .B(_10452_),
    .Y(_10453_));
 sky130_fd_sc_hd__nand2_2 _20629_ (.A(_10032_),
    .B(_10052_),
    .Y(_10454_));
 sky130_fd_sc_hd__nand2_2 _20630_ (.A(_10454_),
    .B(_10050_),
    .Y(_10455_));
 sky130_fd_sc_hd__xor2_1 _20631_ (.A(_10040_),
    .B(_10455_),
    .X(_10456_));
 sky130_fd_sc_hd__nand2_1 _20632_ (.A(_10456_),
    .B(_07146_),
    .Y(_10457_));
 sky130_fd_sc_hd__or2_1 _20633_ (.A(_10041_),
    .B(_10455_),
    .X(_10458_));
 sky130_fd_sc_hd__nand2_1 _20634_ (.A(_10455_),
    .B(_10041_),
    .Y(_10460_));
 sky130_fd_sc_hd__nand3_2 _20635_ (.A(_10458_),
    .B(_07149_),
    .C(_10460_),
    .Y(_10461_));
 sky130_fd_sc_hd__or2_1 _20636_ (.A(_10052_),
    .B(_10032_),
    .X(_10462_));
 sky130_fd_sc_hd__nand2_1 _20637_ (.A(_10462_),
    .B(_10454_),
    .Y(_10463_));
 sky130_fd_sc_hd__nand2_1 _20638_ (.A(_10463_),
    .B(_07155_),
    .Y(_10464_));
 sky130_fd_sc_hd__nand3_2 _20639_ (.A(_10462_),
    .B(_07157_),
    .C(_10454_),
    .Y(_10465_));
 sky130_fd_sc_hd__nand2_1 _20640_ (.A(_10464_),
    .B(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__inv_2 _20641_ (.A(_10466_),
    .Y(_10467_));
 sky130_fd_sc_hd__nand3_1 _20642_ (.A(_10457_),
    .B(_10461_),
    .C(_10467_),
    .Y(_10468_));
 sky130_fd_sc_hd__inv_2 _20643_ (.A(_10468_),
    .Y(_10469_));
 sky130_fd_sc_hd__nand2_1 _20644_ (.A(_10447_),
    .B(_10449_),
    .Y(_10471_));
 sky130_fd_sc_hd__nand2_1 _20645_ (.A(_10471_),
    .B(_08738_),
    .Y(_10472_));
 sky130_fd_sc_hd__nand3_2 _20646_ (.A(_10453_),
    .B(_10469_),
    .C(_10472_),
    .Y(_10473_));
 sky130_fd_sc_hd__inv_2 _20647_ (.A(_10465_),
    .Y(_10474_));
 sky130_fd_sc_hd__a21boi_1 _20648_ (.A1(_10457_),
    .A2(_10474_),
    .B1_N(_10461_),
    .Y(_10475_));
 sky130_fd_sc_hd__nand2_1 _20649_ (.A(_10473_),
    .B(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__or2_1 _20650_ (.A(_10445_),
    .B(_10476_),
    .X(_10477_));
 sky130_fd_sc_hd__inv_6 _20651_ (.A(_10299_),
    .Y(_10478_));
 sky130_fd_sc_hd__nand2_1 _20652_ (.A(_10476_),
    .B(_10445_),
    .Y(_10479_));
 sky130_fd_sc_hd__nand3_1 _20653_ (.A(_10477_),
    .B(_10478_),
    .C(_10479_),
    .Y(_10480_));
 sky130_fd_sc_hd__nand2_1 _20654_ (.A(net225),
    .B(_10441_),
    .Y(_10482_));
 sky130_fd_sc_hd__nand2_1 _20655_ (.A(_10480_),
    .B(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__nand2_1 _20656_ (.A(_10483_),
    .B(_06731_),
    .Y(_10484_));
 sky130_fd_sc_hd__nand3_1 _20657_ (.A(_10480_),
    .B(_06733_),
    .C(_10482_),
    .Y(_10485_));
 sky130_fd_sc_hd__nand2_2 _20658_ (.A(_10484_),
    .B(_10485_),
    .Y(_10486_));
 sky130_fd_sc_hd__nand3_1 _20659_ (.A(_10453_),
    .B(_10472_),
    .C(_10467_),
    .Y(_10487_));
 sky130_fd_sc_hd__nand2_1 _20660_ (.A(_10487_),
    .B(_10465_),
    .Y(_10488_));
 sky130_fd_sc_hd__nand3_1 _20661_ (.A(_10488_),
    .B(_10461_),
    .C(_10457_),
    .Y(_10489_));
 sky130_fd_sc_hd__nand2_1 _20662_ (.A(_10457_),
    .B(_10461_),
    .Y(_10490_));
 sky130_fd_sc_hd__nand3_1 _20663_ (.A(_10487_),
    .B(_10490_),
    .C(_10465_),
    .Y(_10491_));
 sky130_fd_sc_hd__a21o_1 _20664_ (.A1(_10489_),
    .A2(_10491_),
    .B1(_10300_),
    .X(_10493_));
 sky130_fd_sc_hd__nand2_2 _20665_ (.A(net225),
    .B(_10456_),
    .Y(_10494_));
 sky130_fd_sc_hd__nand2_1 _20666_ (.A(_10493_),
    .B(_10494_),
    .Y(_10495_));
 sky130_fd_sc_hd__nand2_1 _20667_ (.A(_10495_),
    .B(_06721_),
    .Y(_10496_));
 sky130_fd_sc_hd__nand3_4 _20668_ (.A(_10493_),
    .B(_06723_),
    .C(_10494_),
    .Y(_10497_));
 sky130_fd_sc_hd__nand2_2 _20669_ (.A(_10497_),
    .B(_10496_),
    .Y(_10498_));
 sky130_fd_sc_hd__nor2_2 _20670_ (.A(_10486_),
    .B(_10498_),
    .Y(_10499_));
 sky130_fd_sc_hd__a21o_1 _20671_ (.A1(_10453_),
    .A2(_10472_),
    .B1(_10467_),
    .X(_10500_));
 sky130_fd_sc_hd__nand3_1 _20672_ (.A(_10478_),
    .B(_10487_),
    .C(_10500_),
    .Y(_10501_));
 sky130_fd_sc_hd__a21o_1 _20673_ (.A1(_10296_),
    .A2(_10298_),
    .B1(_10463_),
    .X(_10502_));
 sky130_fd_sc_hd__nand2_1 _20674_ (.A(_10501_),
    .B(_10502_),
    .Y(_10504_));
 sky130_fd_sc_hd__nand2_1 _20675_ (.A(_10504_),
    .B(_06695_),
    .Y(_10505_));
 sky130_fd_sc_hd__nand3_1 _20676_ (.A(_10501_),
    .B(_06697_),
    .C(_10502_),
    .Y(_10506_));
 sky130_fd_sc_hd__nand2_1 _20677_ (.A(_10505_),
    .B(_10506_),
    .Y(_10507_));
 sky130_fd_sc_hd__nand2_1 _20678_ (.A(_10472_),
    .B(_10450_),
    .Y(_10508_));
 sky130_fd_sc_hd__nand2_1 _20679_ (.A(_10378_),
    .B(_10344_),
    .Y(_10509_));
 sky130_fd_sc_hd__xor2_1 _20680_ (.A(_10508_),
    .B(_10509_),
    .X(_10510_));
 sky130_fd_sc_hd__nand2_1 _20681_ (.A(_10478_),
    .B(_10510_),
    .Y(_10511_));
 sky130_fd_sc_hd__nand2_1 _20682_ (.A(_10300_),
    .B(_10471_),
    .Y(_10512_));
 sky130_fd_sc_hd__nand2_1 _20683_ (.A(_10511_),
    .B(_10512_),
    .Y(_10513_));
 sky130_fd_sc_hd__or2_4 _20684_ (.A(_09410_),
    .B(_10513_),
    .X(_10515_));
 sky130_fd_sc_hd__nand2_1 _20685_ (.A(_10513_),
    .B(_09410_),
    .Y(_10516_));
 sky130_fd_sc_hd__nand2_1 _20686_ (.A(_10515_),
    .B(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__nor2_1 _20687_ (.A(_10507_),
    .B(_10517_),
    .Y(_10518_));
 sky130_fd_sc_hd__nand2_1 _20688_ (.A(_10499_),
    .B(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__inv_2 _20689_ (.A(_10519_),
    .Y(_10520_));
 sky130_fd_sc_hd__nand2_1 _20690_ (.A(_10431_),
    .B(_10520_),
    .Y(_10521_));
 sky130_fd_sc_hd__o21ai_2 _20691_ (.A1(_10515_),
    .A2(_10507_),
    .B1(_10505_),
    .Y(_10522_));
 sky130_fd_sc_hd__o21ai_1 _20692_ (.A1(_10497_),
    .A2(_10486_),
    .B1(_10484_),
    .Y(_10523_));
 sky130_fd_sc_hd__a21oi_1 _20693_ (.A1(_10522_),
    .A2(_10499_),
    .B1(_10523_),
    .Y(_10524_));
 sky130_fd_sc_hd__nand2_2 _20694_ (.A(_10521_),
    .B(_10524_),
    .Y(_10526_));
 sky130_fd_sc_hd__inv_2 _20695_ (.A(_10473_),
    .Y(_10527_));
 sky130_fd_sc_hd__nand2_1 _20696_ (.A(_10438_),
    .B(_10063_),
    .Y(_10528_));
 sky130_fd_sc_hd__inv_2 _20697_ (.A(_10072_),
    .Y(_10529_));
 sky130_fd_sc_hd__nand2_1 _20698_ (.A(_10528_),
    .B(_10529_),
    .Y(_10530_));
 sky130_fd_sc_hd__nand3_1 _20699_ (.A(_10438_),
    .B(_10072_),
    .C(_10063_),
    .Y(_10531_));
 sky130_fd_sc_hd__nand2_1 _20700_ (.A(_10530_),
    .B(_10531_),
    .Y(_10532_));
 sky130_fd_sc_hd__nand2_1 _20701_ (.A(_10532_),
    .B(_07226_),
    .Y(_10533_));
 sky130_fd_sc_hd__nand3_1 _20702_ (.A(_10530_),
    .B(_07228_),
    .C(_10531_),
    .Y(_10534_));
 sky130_fd_sc_hd__nand3_1 _20703_ (.A(_10445_),
    .B(_10533_),
    .C(_10534_),
    .Y(_10535_));
 sky130_fd_sc_hd__inv_2 _20704_ (.A(_10535_),
    .Y(_10537_));
 sky130_fd_sc_hd__nand2_1 _20705_ (.A(_10527_),
    .B(_10537_),
    .Y(_10538_));
 sky130_fd_sc_hd__nor2_1 _20706_ (.A(_10475_),
    .B(_10535_),
    .Y(_10539_));
 sky130_fd_sc_hd__nand2_1 _20707_ (.A(_10533_),
    .B(_10534_),
    .Y(_10540_));
 sky130_fd_sc_hd__o21ai_1 _20708_ (.A1(_10442_),
    .A2(_10540_),
    .B1(_10534_),
    .Y(_10541_));
 sky130_fd_sc_hd__nor2_1 _20709_ (.A(_10539_),
    .B(_10541_),
    .Y(_10542_));
 sky130_fd_sc_hd__nand2_1 _20710_ (.A(_10538_),
    .B(_10542_),
    .Y(_10543_));
 sky130_fd_sc_hd__inv_2 _20711_ (.A(_10087_),
    .Y(_10544_));
 sky130_fd_sc_hd__inv_2 _20712_ (.A(_10085_),
    .Y(_10545_));
 sky130_fd_sc_hd__nand2_1 _20713_ (.A(_10082_),
    .B(_10545_),
    .Y(_10546_));
 sky130_fd_sc_hd__nand2_1 _20714_ (.A(_10546_),
    .B(_09937_),
    .Y(_10548_));
 sky130_fd_sc_hd__or2_1 _20715_ (.A(_10544_),
    .B(_10548_),
    .X(_10549_));
 sky130_fd_sc_hd__nand2_1 _20716_ (.A(_10548_),
    .B(_10544_),
    .Y(_10550_));
 sky130_fd_sc_hd__nand2_1 _20717_ (.A(_10549_),
    .B(_10550_),
    .Y(_10551_));
 sky130_fd_sc_hd__nand2_1 _20718_ (.A(_10551_),
    .B(_07247_),
    .Y(_10552_));
 sky130_fd_sc_hd__nand3_1 _20719_ (.A(_10549_),
    .B(_07249_),
    .C(_10550_),
    .Y(_10553_));
 sky130_fd_sc_hd__nand2_1 _20720_ (.A(_10552_),
    .B(_10553_),
    .Y(_10554_));
 sky130_fd_sc_hd__inv_2 _20721_ (.A(_10554_),
    .Y(_10555_));
 sky130_fd_sc_hd__or2_1 _20722_ (.A(_10545_),
    .B(_10082_),
    .X(_10556_));
 sky130_fd_sc_hd__nand2_1 _20723_ (.A(_10556_),
    .B(_10546_),
    .Y(_10557_));
 sky130_fd_sc_hd__inv_2 _20724_ (.A(_10557_),
    .Y(_10559_));
 sky130_fd_sc_hd__nand2_1 _20725_ (.A(_10559_),
    .B(_06521_),
    .Y(_10560_));
 sky130_fd_sc_hd__nand2_1 _20726_ (.A(_10557_),
    .B(_07677_),
    .Y(_10561_));
 sky130_fd_sc_hd__nand2_2 _20727_ (.A(_10560_),
    .B(_10561_),
    .Y(_10562_));
 sky130_fd_sc_hd__inv_4 _20728_ (.A(_10562_),
    .Y(_10563_));
 sky130_fd_sc_hd__nand2_1 _20729_ (.A(_10555_),
    .B(_10563_),
    .Y(_10564_));
 sky130_fd_sc_hd__inv_2 _20730_ (.A(_10564_),
    .Y(_10565_));
 sky130_fd_sc_hd__nand2_1 _20731_ (.A(_10543_),
    .B(_10565_),
    .Y(_10566_));
 sky130_fd_sc_hd__inv_2 _20732_ (.A(_10560_),
    .Y(_10567_));
 sky130_fd_sc_hd__a21boi_2 _20733_ (.A1(_10552_),
    .A2(_10567_),
    .B1_N(_10553_),
    .Y(_10568_));
 sky130_fd_sc_hd__nand2_1 _20734_ (.A(_10566_),
    .B(_10568_),
    .Y(_10570_));
 sky130_fd_sc_hd__nand2_1 _20735_ (.A(_10082_),
    .B(_10088_),
    .Y(_10571_));
 sky130_fd_sc_hd__inv_2 _20736_ (.A(_09946_),
    .Y(_10572_));
 sky130_fd_sc_hd__nand2_1 _20737_ (.A(_10571_),
    .B(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__inv_2 _20738_ (.A(_09924_),
    .Y(_10574_));
 sky130_fd_sc_hd__nand2_1 _20739_ (.A(_10573_),
    .B(_10574_),
    .Y(_10575_));
 sky130_fd_sc_hd__nand3_1 _20740_ (.A(_10571_),
    .B(_10572_),
    .C(_09924_),
    .Y(_10576_));
 sky130_fd_sc_hd__nand2_1 _20741_ (.A(_10575_),
    .B(_10576_),
    .Y(_10577_));
 sky130_fd_sc_hd__nand2_1 _20742_ (.A(_10577_),
    .B(_07276_),
    .Y(_10578_));
 sky130_fd_sc_hd__nand3_1 _20743_ (.A(_10575_),
    .B(_10576_),
    .C(_07278_),
    .Y(_10579_));
 sky130_fd_sc_hd__nand2_1 _20744_ (.A(_10578_),
    .B(_10579_),
    .Y(_10581_));
 sky130_fd_sc_hd__inv_2 _20745_ (.A(_10581_),
    .Y(_10582_));
 sky130_fd_sc_hd__nand2_1 _20746_ (.A(_10570_),
    .B(_10582_),
    .Y(_10583_));
 sky130_fd_sc_hd__nand3_1 _20747_ (.A(_10566_),
    .B(_10581_),
    .C(_10568_),
    .Y(_10584_));
 sky130_fd_sc_hd__nand3_1 _20748_ (.A(_10583_),
    .B(_10478_),
    .C(_10584_),
    .Y(_10585_));
 sky130_fd_sc_hd__or2_1 _20749_ (.A(_10577_),
    .B(_10478_),
    .X(_10586_));
 sky130_fd_sc_hd__nand2_1 _20750_ (.A(_10585_),
    .B(_10586_),
    .Y(_10587_));
 sky130_fd_sc_hd__nand2_1 _20751_ (.A(_10587_),
    .B(_06554_),
    .Y(_10588_));
 sky130_fd_sc_hd__nand3_1 _20752_ (.A(_10585_),
    .B(_06556_),
    .C(_10586_),
    .Y(_10589_));
 sky130_fd_sc_hd__nand2_1 _20753_ (.A(_10588_),
    .B(_10589_),
    .Y(_10590_));
 sky130_fd_sc_hd__nand2_1 _20754_ (.A(_10543_),
    .B(_10563_),
    .Y(_10592_));
 sky130_fd_sc_hd__nand2_1 _20755_ (.A(_10592_),
    .B(_10560_),
    .Y(_10593_));
 sky130_fd_sc_hd__nand2_1 _20756_ (.A(_10593_),
    .B(_10555_),
    .Y(_10594_));
 sky130_fd_sc_hd__nand3_1 _20757_ (.A(_10592_),
    .B(_10554_),
    .C(_10560_),
    .Y(_10595_));
 sky130_fd_sc_hd__nand2_1 _20758_ (.A(_10594_),
    .B(_10595_),
    .Y(_10596_));
 sky130_fd_sc_hd__nand2_1 _20759_ (.A(_10596_),
    .B(_10478_),
    .Y(_10597_));
 sky130_fd_sc_hd__nand2_1 _20760_ (.A(\div1i.quot[11] ),
    .B(_10551_),
    .Y(_10598_));
 sky130_fd_sc_hd__nand2_1 _20761_ (.A(_10597_),
    .B(_10598_),
    .Y(_10599_));
 sky130_fd_sc_hd__nand2_1 _20762_ (.A(_10599_),
    .B(_06568_),
    .Y(_10600_));
 sky130_fd_sc_hd__nand3_2 _20763_ (.A(_10597_),
    .B(_06570_),
    .C(_10598_),
    .Y(_10601_));
 sky130_fd_sc_hd__nand2_2 _20764_ (.A(_10600_),
    .B(_10601_),
    .Y(_10603_));
 sky130_fd_sc_hd__nor2_2 _20765_ (.A(_10590_),
    .B(_10603_),
    .Y(_10604_));
 sky130_fd_sc_hd__or2_1 _20766_ (.A(_10563_),
    .B(_10543_),
    .X(_10605_));
 sky130_fd_sc_hd__nand3_1 _20767_ (.A(_10605_),
    .B(_10478_),
    .C(_10592_),
    .Y(_10606_));
 sky130_fd_sc_hd__nand2_1 _20768_ (.A(net225),
    .B(_10559_),
    .Y(_10607_));
 sky130_fd_sc_hd__nand2_1 _20769_ (.A(_10606_),
    .B(_10607_),
    .Y(_10608_));
 sky130_fd_sc_hd__nand2_1 _20770_ (.A(_10608_),
    .B(_06149_),
    .Y(_10609_));
 sky130_fd_sc_hd__nand3_1 _20771_ (.A(_10606_),
    .B(_09944_),
    .C(_10607_),
    .Y(_10610_));
 sky130_fd_sc_hd__nand2_1 _20772_ (.A(_10609_),
    .B(_10610_),
    .Y(_10611_));
 sky130_fd_sc_hd__nand2_1 _20773_ (.A(_10479_),
    .B(_10442_),
    .Y(_10612_));
 sky130_fd_sc_hd__xor2_1 _20774_ (.A(_10540_),
    .B(_10612_),
    .X(_10614_));
 sky130_fd_sc_hd__nand2_1 _20775_ (.A(_10614_),
    .B(_10478_),
    .Y(_10615_));
 sky130_fd_sc_hd__nand2_1 _20776_ (.A(\div1i.quot[11] ),
    .B(_10532_),
    .Y(_10616_));
 sky130_fd_sc_hd__nand2_1 _20777_ (.A(_10615_),
    .B(_10616_),
    .Y(_10617_));
 sky130_fd_sc_hd__nand2_1 _20778_ (.A(_10617_),
    .B(_06159_),
    .Y(_10618_));
 sky130_fd_sc_hd__nand3_2 _20779_ (.A(_10615_),
    .B(_07318_),
    .C(_10616_),
    .Y(_10619_));
 sky130_fd_sc_hd__nand2_2 _20780_ (.A(_10618_),
    .B(_10619_),
    .Y(_10620_));
 sky130_fd_sc_hd__nor2_2 _20781_ (.A(_10620_),
    .B(_10611_),
    .Y(_10621_));
 sky130_fd_sc_hd__nand2_1 _20782_ (.A(_10604_),
    .B(_10621_),
    .Y(_10622_));
 sky130_fd_sc_hd__inv_2 _20783_ (.A(_10622_),
    .Y(_10623_));
 sky130_fd_sc_hd__nand2_2 _20784_ (.A(_10526_),
    .B(_10623_),
    .Y(_10625_));
 sky130_fd_sc_hd__o21ai_2 _20785_ (.A1(_10619_),
    .A2(_10611_),
    .B1(_10609_),
    .Y(_10626_));
 sky130_fd_sc_hd__o21ai_1 _20786_ (.A1(_10601_),
    .A2(_10590_),
    .B1(_10588_),
    .Y(_10627_));
 sky130_fd_sc_hd__a21oi_2 _20787_ (.A1(_10604_),
    .A2(_10626_),
    .B1(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__nand2_4 _20788_ (.A(_10625_),
    .B(_10628_),
    .Y(_10629_));
 sky130_fd_sc_hd__nand2_1 _20789_ (.A(_10575_),
    .B(_09923_),
    .Y(_10630_));
 sky130_fd_sc_hd__inv_2 _20790_ (.A(_09912_),
    .Y(_10631_));
 sky130_fd_sc_hd__nand2_1 _20791_ (.A(_10630_),
    .B(_10631_),
    .Y(_10632_));
 sky130_fd_sc_hd__nand3_1 _20792_ (.A(_10575_),
    .B(_09912_),
    .C(_09923_),
    .Y(_10633_));
 sky130_fd_sc_hd__nand2_1 _20793_ (.A(_10632_),
    .B(_10633_),
    .Y(_10634_));
 sky130_fd_sc_hd__nand2_1 _20794_ (.A(_10634_),
    .B(_07905_),
    .Y(_10636_));
 sky130_fd_sc_hd__nand3_1 _20795_ (.A(_10632_),
    .B(_06772_),
    .C(_10633_),
    .Y(_10637_));
 sky130_fd_sc_hd__nand3_1 _20796_ (.A(_10636_),
    .B(_10637_),
    .C(_10582_),
    .Y(_10638_));
 sky130_fd_sc_hd__nor2_1 _20797_ (.A(_10638_),
    .B(_10564_),
    .Y(_10639_));
 sky130_fd_sc_hd__nand2_2 _20798_ (.A(_10543_),
    .B(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__nor2_1 _20799_ (.A(_10638_),
    .B(_10568_),
    .Y(_10641_));
 sky130_fd_sc_hd__nand2_1 _20800_ (.A(_10636_),
    .B(_10637_),
    .Y(_10642_));
 sky130_fd_sc_hd__o21ai_1 _20801_ (.A1(_10579_),
    .A2(_10642_),
    .B1(_10637_),
    .Y(_10643_));
 sky130_fd_sc_hd__nor2_1 _20802_ (.A(_10641_),
    .B(_10643_),
    .Y(_10644_));
 sky130_fd_sc_hd__nand2_2 _20803_ (.A(_10640_),
    .B(_10644_),
    .Y(_10645_));
 sky130_fd_sc_hd__clkinvlp_2 _20804_ (.A(_10125_),
    .Y(_10647_));
 sky130_fd_sc_hd__inv_2 _20805_ (.A(_10135_),
    .Y(_10648_));
 sky130_fd_sc_hd__nand2_1 _20806_ (.A(_10090_),
    .B(_10648_),
    .Y(_10649_));
 sky130_fd_sc_hd__nand2_1 _20807_ (.A(_10649_),
    .B(_10134_),
    .Y(_10650_));
 sky130_fd_sc_hd__or2_1 _20808_ (.A(_10647_),
    .B(_10650_),
    .X(_10651_));
 sky130_fd_sc_hd__nand2_1 _20809_ (.A(_10650_),
    .B(_10647_),
    .Y(_10652_));
 sky130_fd_sc_hd__nand2_1 _20810_ (.A(_10651_),
    .B(_10652_),
    .Y(_10653_));
 sky130_fd_sc_hd__nand2_1 _20811_ (.A(_10653_),
    .B(_07957_),
    .Y(_10654_));
 sky130_fd_sc_hd__nand3_1 _20812_ (.A(_10651_),
    .B(_06827_),
    .C(_10652_),
    .Y(_10655_));
 sky130_fd_sc_hd__nand2_1 _20813_ (.A(_10654_),
    .B(_10655_),
    .Y(_10656_));
 sky130_fd_sc_hd__or2_1 _20814_ (.A(_10648_),
    .B(_10090_),
    .X(_10658_));
 sky130_fd_sc_hd__nand2_1 _20815_ (.A(_10658_),
    .B(_10649_),
    .Y(_10659_));
 sky130_fd_sc_hd__inv_2 _20816_ (.A(_10659_),
    .Y(_10660_));
 sky130_fd_sc_hd__nand2_1 _20817_ (.A(_10660_),
    .B(_06207_),
    .Y(_10661_));
 sky130_fd_sc_hd__nand2_1 _20818_ (.A(_10659_),
    .B(_08465_),
    .Y(_10662_));
 sky130_fd_sc_hd__nand2_1 _20819_ (.A(_10661_),
    .B(_10662_),
    .Y(_10663_));
 sky130_fd_sc_hd__inv_2 _20820_ (.A(_10663_),
    .Y(_10664_));
 sky130_fd_sc_hd__nand2b_1 _20821_ (.A_N(_10656_),
    .B(_10664_),
    .Y(_10665_));
 sky130_fd_sc_hd__inv_2 _20822_ (.A(_10665_),
    .Y(_10666_));
 sky130_fd_sc_hd__nand2_1 _20823_ (.A(_10645_),
    .B(_10666_),
    .Y(_10667_));
 sky130_fd_sc_hd__inv_2 _20824_ (.A(_10661_),
    .Y(_10669_));
 sky130_fd_sc_hd__a21boi_2 _20825_ (.A1(_10654_),
    .A2(_10669_),
    .B1_N(_10655_),
    .Y(_10670_));
 sky130_fd_sc_hd__nand2_1 _20826_ (.A(_10667_),
    .B(_10670_),
    .Y(_10671_));
 sky130_fd_sc_hd__inv_2 _20827_ (.A(_10182_),
    .Y(_10672_));
 sky130_fd_sc_hd__nand2_1 _20828_ (.A(_10142_),
    .B(_10672_),
    .Y(_10673_));
 sky130_fd_sc_hd__nand3_1 _20829_ (.A(_10137_),
    .B(_10140_),
    .C(_10182_),
    .Y(_10674_));
 sky130_fd_sc_hd__nand2_1 _20830_ (.A(_10673_),
    .B(_10674_),
    .Y(_10675_));
 sky130_fd_sc_hd__inv_2 _20831_ (.A(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__nand2_1 _20832_ (.A(_10676_),
    .B(_06819_),
    .Y(_10677_));
 sky130_fd_sc_hd__nand2_1 _20833_ (.A(_10675_),
    .B(_07948_),
    .Y(_10678_));
 sky130_fd_sc_hd__nand2_1 _20834_ (.A(_10677_),
    .B(_10678_),
    .Y(_10680_));
 sky130_fd_sc_hd__inv_2 _20835_ (.A(_10680_),
    .Y(_10681_));
 sky130_fd_sc_hd__nand2_1 _20836_ (.A(_10671_),
    .B(_10681_),
    .Y(_10682_));
 sky130_fd_sc_hd__buf_6 _20837_ (.A(_10478_),
    .X(_10683_));
 sky130_fd_sc_hd__nand3_1 _20838_ (.A(_10667_),
    .B(_10680_),
    .C(_10670_),
    .Y(_10684_));
 sky130_fd_sc_hd__nand3_1 _20839_ (.A(_10682_),
    .B(_10683_),
    .C(_10684_),
    .Y(_10685_));
 sky130_fd_sc_hd__nand2_1 _20840_ (.A(\div1i.quot[11] ),
    .B(_10676_),
    .Y(_10686_));
 sky130_fd_sc_hd__nand2_1 _20841_ (.A(_10685_),
    .B(_10686_),
    .Y(_10687_));
 sky130_fd_sc_hd__nand2_1 _20842_ (.A(_10687_),
    .B(_06856_),
    .Y(_10688_));
 sky130_fd_sc_hd__nand3_1 _20843_ (.A(_10685_),
    .B(_06809_),
    .C(_10686_),
    .Y(_10689_));
 sky130_fd_sc_hd__nand2_1 _20844_ (.A(_10688_),
    .B(_10689_),
    .Y(_10691_));
 sky130_fd_sc_hd__nand2_1 _20845_ (.A(_10645_),
    .B(_10664_),
    .Y(_10692_));
 sky130_fd_sc_hd__nand2_1 _20846_ (.A(_10692_),
    .B(_10661_),
    .Y(_10693_));
 sky130_fd_sc_hd__xor2_1 _20847_ (.A(_10656_),
    .B(_10693_),
    .X(_10694_));
 sky130_fd_sc_hd__nand2_1 _20848_ (.A(_10694_),
    .B(_10683_),
    .Y(_10695_));
 sky130_fd_sc_hd__nand2_1 _20849_ (.A(\div1i.quot[11] ),
    .B(_10653_),
    .Y(_10696_));
 sky130_fd_sc_hd__nand2_1 _20850_ (.A(_10695_),
    .B(_10696_),
    .Y(_10697_));
 sky130_fd_sc_hd__nand2_1 _20851_ (.A(_10697_),
    .B(_10173_),
    .Y(_10698_));
 sky130_fd_sc_hd__nand3_2 _20852_ (.A(_10695_),
    .B(_07400_),
    .C(_10696_),
    .Y(_10699_));
 sky130_fd_sc_hd__nand2_1 _20853_ (.A(_10698_),
    .B(_10699_),
    .Y(_10700_));
 sky130_fd_sc_hd__nor2_2 _20854_ (.A(_10691_),
    .B(_10700_),
    .Y(_10702_));
 sky130_fd_sc_hd__nand3_1 _20855_ (.A(_10640_),
    .B(_10644_),
    .C(_10663_),
    .Y(_10703_));
 sky130_fd_sc_hd__nand3_1 _20856_ (.A(_10692_),
    .B(_10478_),
    .C(_10703_),
    .Y(_10704_));
 sky130_fd_sc_hd__nand2_1 _20857_ (.A(net225),
    .B(_10660_),
    .Y(_10705_));
 sky130_fd_sc_hd__nand2_1 _20858_ (.A(_10704_),
    .B(_10705_),
    .Y(_10706_));
 sky130_fd_sc_hd__or2_1 _20859_ (.A(_10138_),
    .B(_10706_),
    .X(_10707_));
 sky130_fd_sc_hd__nand2_1 _20860_ (.A(_10706_),
    .B(_10138_),
    .Y(_10708_));
 sky130_fd_sc_hd__nand2_1 _20861_ (.A(_10707_),
    .B(_10708_),
    .Y(_10709_));
 sky130_fd_sc_hd__nand2_1 _20862_ (.A(_10583_),
    .B(_10579_),
    .Y(_10710_));
 sky130_fd_sc_hd__xor2_1 _20863_ (.A(_10642_),
    .B(_10710_),
    .X(_10711_));
 sky130_fd_sc_hd__nand2_1 _20864_ (.A(_10711_),
    .B(_10683_),
    .Y(_10713_));
 sky130_fd_sc_hd__nand2_1 _20865_ (.A(\div1i.quot[11] ),
    .B(_10634_),
    .Y(_10714_));
 sky130_fd_sc_hd__nand2_1 _20866_ (.A(_10713_),
    .B(_10714_),
    .Y(_10715_));
 sky130_fd_sc_hd__nand2_1 _20867_ (.A(_10715_),
    .B(_06797_),
    .Y(_10716_));
 sky130_fd_sc_hd__nand3_2 _20868_ (.A(_10713_),
    .B(_06799_),
    .C(_10714_),
    .Y(_10717_));
 sky130_fd_sc_hd__nand3b_1 _20869_ (.A_N(_10709_),
    .B(_10716_),
    .C(_10717_),
    .Y(_10718_));
 sky130_fd_sc_hd__inv_2 _20870_ (.A(_10718_),
    .Y(_10719_));
 sky130_fd_sc_hd__nand3_4 _20871_ (.A(_10629_),
    .B(_10702_),
    .C(_10719_),
    .Y(_10720_));
 sky130_fd_sc_hd__o21ai_1 _20872_ (.A1(_10709_),
    .A2(_10717_),
    .B1(_10708_),
    .Y(_10721_));
 sky130_fd_sc_hd__o21ai_1 _20873_ (.A1(_10691_),
    .A2(_10699_),
    .B1(_10688_),
    .Y(_10722_));
 sky130_fd_sc_hd__a21oi_2 _20874_ (.A1(_10702_),
    .A2(_10721_),
    .B1(_10722_),
    .Y(_10724_));
 sky130_fd_sc_hd__nand2_4 _20875_ (.A(_10720_),
    .B(_10724_),
    .Y(_10725_));
 sky130_fd_sc_hd__nand2_1 _20876_ (.A(_10673_),
    .B(_10180_),
    .Y(_10726_));
 sky130_fd_sc_hd__inv_2 _20877_ (.A(_10172_),
    .Y(_10727_));
 sky130_fd_sc_hd__nand2_1 _20878_ (.A(_10726_),
    .B(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__nand3_1 _20879_ (.A(_10673_),
    .B(_10172_),
    .C(_10180_),
    .Y(_10729_));
 sky130_fd_sc_hd__nand2_1 _20880_ (.A(_10728_),
    .B(_10729_),
    .Y(_10730_));
 sky130_fd_sc_hd__nand2_1 _20881_ (.A(_10730_),
    .B(_08001_),
    .Y(_10731_));
 sky130_fd_sc_hd__nand3_1 _20882_ (.A(_10728_),
    .B(_06874_),
    .C(_10729_),
    .Y(_10732_));
 sky130_fd_sc_hd__nand3_1 _20883_ (.A(_10681_),
    .B(_10731_),
    .C(_10732_),
    .Y(_10733_));
 sky130_fd_sc_hd__inv_2 _20884_ (.A(_10733_),
    .Y(_10735_));
 sky130_fd_sc_hd__nand3_2 _20885_ (.A(_10645_),
    .B(_10666_),
    .C(_10735_),
    .Y(_10736_));
 sky130_fd_sc_hd__inv_2 _20886_ (.A(_10731_),
    .Y(_10737_));
 sky130_fd_sc_hd__o21ai_1 _20887_ (.A1(_10677_),
    .A2(_10737_),
    .B1(_10732_),
    .Y(_10738_));
 sky130_fd_sc_hd__nor2_1 _20888_ (.A(_10670_),
    .B(_10733_),
    .Y(_10739_));
 sky130_fd_sc_hd__nor2_1 _20889_ (.A(_10738_),
    .B(_10739_),
    .Y(_10740_));
 sky130_fd_sc_hd__nand2_1 _20890_ (.A(_10736_),
    .B(_10740_),
    .Y(_10741_));
 sky130_fd_sc_hd__inv_2 _20891_ (.A(_10188_),
    .Y(_10742_));
 sky130_fd_sc_hd__nand2_1 _20892_ (.A(_10233_),
    .B(_10234_),
    .Y(_10743_));
 sky130_fd_sc_hd__nand2_1 _20893_ (.A(_10742_),
    .B(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__inv_2 _20894_ (.A(_10743_),
    .Y(_10746_));
 sky130_fd_sc_hd__nand2_1 _20895_ (.A(_10188_),
    .B(_10746_),
    .Y(_10747_));
 sky130_fd_sc_hd__nand2_1 _20896_ (.A(_10744_),
    .B(_10747_),
    .Y(_10748_));
 sky130_fd_sc_hd__buf_6 _20897_ (.A(_07450_),
    .X(_10749_));
 sky130_fd_sc_hd__nand2_1 _20898_ (.A(_10748_),
    .B(_10749_),
    .Y(_10750_));
 sky130_fd_sc_hd__nand3_2 _20899_ (.A(_10744_),
    .B(_08554_),
    .C(_10747_),
    .Y(_10751_));
 sky130_fd_sc_hd__nand2_1 _20900_ (.A(_10750_),
    .B(_10751_),
    .Y(_10752_));
 sky130_fd_sc_hd__inv_2 _20901_ (.A(_10752_),
    .Y(_10753_));
 sky130_fd_sc_hd__nand2_1 _20902_ (.A(_10741_),
    .B(_10753_),
    .Y(_10754_));
 sky130_fd_sc_hd__nand2_1 _20903_ (.A(_10754_),
    .B(_10751_),
    .Y(_10755_));
 sky130_fd_sc_hd__nand2_1 _20904_ (.A(_10747_),
    .B(_10234_),
    .Y(_10757_));
 sky130_fd_sc_hd__xor2_2 _20905_ (.A(_10224_),
    .B(_10757_),
    .X(_10758_));
 sky130_fd_sc_hd__inv_2 _20906_ (.A(_10758_),
    .Y(_10759_));
 sky130_fd_sc_hd__nand2_1 _20907_ (.A(_10759_),
    .B(_07461_),
    .Y(_10760_));
 sky130_fd_sc_hd__nand2_1 _20908_ (.A(_10758_),
    .B(_08041_),
    .Y(_10761_));
 sky130_fd_sc_hd__nand2_1 _20909_ (.A(_10760_),
    .B(_10761_),
    .Y(_10762_));
 sky130_fd_sc_hd__inv_2 _20910_ (.A(_10762_),
    .Y(_10763_));
 sky130_fd_sc_hd__nand2_1 _20911_ (.A(_10755_),
    .B(_10763_),
    .Y(_10764_));
 sky130_fd_sc_hd__nand3_1 _20912_ (.A(_10754_),
    .B(_10762_),
    .C(_10751_),
    .Y(_10765_));
 sky130_fd_sc_hd__nand2_1 _20913_ (.A(_10764_),
    .B(_10765_),
    .Y(_10766_));
 sky130_fd_sc_hd__nand2_1 _20914_ (.A(_10766_),
    .B(_10683_),
    .Y(_10768_));
 sky130_fd_sc_hd__nand2_1 _20915_ (.A(_10758_),
    .B(\div1i.quot[11] ),
    .Y(_10769_));
 sky130_fd_sc_hd__nand2_1 _20916_ (.A(_10768_),
    .B(_10769_),
    .Y(_10770_));
 sky130_fd_sc_hd__nand2_1 _20917_ (.A(_10770_),
    .B(_07474_),
    .Y(_10771_));
 sky130_fd_sc_hd__nand3_1 _20918_ (.A(_10768_),
    .B(_06366_),
    .C(_10769_),
    .Y(_10772_));
 sky130_fd_sc_hd__nand2_1 _20919_ (.A(_10771_),
    .B(_10772_),
    .Y(_10773_));
 sky130_fd_sc_hd__inv_2 _20920_ (.A(_10773_),
    .Y(_10774_));
 sky130_fd_sc_hd__nand3_1 _20921_ (.A(_10760_),
    .B(_10761_),
    .C(_10753_),
    .Y(_10775_));
 sky130_fd_sc_hd__inv_2 _20922_ (.A(_10775_),
    .Y(_10776_));
 sky130_fd_sc_hd__nand2_1 _20923_ (.A(_10776_),
    .B(_10741_),
    .Y(_10777_));
 sky130_fd_sc_hd__inv_2 _20924_ (.A(_10761_),
    .Y(_10779_));
 sky130_fd_sc_hd__o21a_1 _20925_ (.A1(_10751_),
    .A2(_10779_),
    .B1(_10760_),
    .X(_10780_));
 sky130_fd_sc_hd__nand2_1 _20926_ (.A(_10777_),
    .B(_10780_),
    .Y(_10781_));
 sky130_fd_sc_hd__o21bai_1 _20927_ (.A1(_10235_),
    .A2(_10742_),
    .B1_N(_10286_),
    .Y(_10782_));
 sky130_fd_sc_hd__or2_1 _20928_ (.A(_10256_),
    .B(_10782_),
    .X(_10783_));
 sky130_fd_sc_hd__nand2_1 _20929_ (.A(_10782_),
    .B(_10256_),
    .Y(_10784_));
 sky130_fd_sc_hd__nand2_1 _20930_ (.A(_10783_),
    .B(_10784_),
    .Y(_10785_));
 sky130_fd_sc_hd__inv_2 _20931_ (.A(_10785_),
    .Y(_10786_));
 sky130_fd_sc_hd__nand2_1 _20932_ (.A(_10786_),
    .B(_06936_),
    .Y(_10787_));
 sky130_fd_sc_hd__nand2_1 _20933_ (.A(_10785_),
    .B(_08611_),
    .Y(_10788_));
 sky130_fd_sc_hd__nand2_1 _20934_ (.A(_10787_),
    .B(_10788_),
    .Y(_10790_));
 sky130_fd_sc_hd__inv_2 _20935_ (.A(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__nand2_1 _20936_ (.A(_10781_),
    .B(_10791_),
    .Y(_10792_));
 sky130_fd_sc_hd__nand3_1 _20937_ (.A(_10777_),
    .B(_10780_),
    .C(_10790_),
    .Y(_10793_));
 sky130_fd_sc_hd__nand3_1 _20938_ (.A(_10792_),
    .B(_10793_),
    .C(_10683_),
    .Y(_10794_));
 sky130_fd_sc_hd__nand2_1 _20939_ (.A(_10786_),
    .B(\div1i.quot[11] ),
    .Y(_10795_));
 sky130_fd_sc_hd__nand2_1 _20940_ (.A(_10794_),
    .B(_10795_),
    .Y(_10796_));
 sky130_fd_sc_hd__nand2_1 _20941_ (.A(_10796_),
    .B(_06947_),
    .Y(_10797_));
 sky130_fd_sc_hd__nand3_1 _20942_ (.A(_10794_),
    .B(_06949_),
    .C(_10795_),
    .Y(_10798_));
 sky130_fd_sc_hd__nand2_2 _20943_ (.A(_10797_),
    .B(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__inv_2 _20944_ (.A(_10799_),
    .Y(_10801_));
 sky130_fd_sc_hd__nand2_1 _20945_ (.A(_10774_),
    .B(_10801_),
    .Y(_10802_));
 sky130_fd_sc_hd__nand3_1 _20946_ (.A(_10736_),
    .B(_10740_),
    .C(_10752_),
    .Y(_10803_));
 sky130_fd_sc_hd__nand3_1 _20947_ (.A(_10754_),
    .B(_10803_),
    .C(_10683_),
    .Y(_10804_));
 sky130_fd_sc_hd__or2_1 _20948_ (.A(_10748_),
    .B(_10683_),
    .X(_10805_));
 sky130_fd_sc_hd__nand2_1 _20949_ (.A(_10804_),
    .B(_10805_),
    .Y(_10806_));
 sky130_fd_sc_hd__or2_1 _20950_ (.A(_09664_),
    .B(_10806_),
    .X(_10807_));
 sky130_fd_sc_hd__nand2_1 _20951_ (.A(_10806_),
    .B(_09664_),
    .Y(_10808_));
 sky130_fd_sc_hd__nand2_2 _20952_ (.A(_10807_),
    .B(_10808_),
    .Y(_10809_));
 sky130_fd_sc_hd__nand2_1 _20953_ (.A(_10731_),
    .B(_10732_),
    .Y(_10810_));
 sky130_fd_sc_hd__nand2_1 _20954_ (.A(_10682_),
    .B(_10677_),
    .Y(_10812_));
 sky130_fd_sc_hd__xor2_1 _20955_ (.A(_10810_),
    .B(_10812_),
    .X(_10813_));
 sky130_fd_sc_hd__nand2_1 _20956_ (.A(_10813_),
    .B(_10683_),
    .Y(_10814_));
 sky130_fd_sc_hd__nand2_1 _20957_ (.A(\div1i.quot[11] ),
    .B(_10730_),
    .Y(_10815_));
 sky130_fd_sc_hd__nand3_2 _20958_ (.A(_10814_),
    .B(_06898_),
    .C(_10815_),
    .Y(_10816_));
 sky130_fd_sc_hd__nand2_1 _20959_ (.A(_10814_),
    .B(_10815_),
    .Y(_10817_));
 sky130_fd_sc_hd__nand2_1 _20960_ (.A(_10817_),
    .B(_06903_),
    .Y(_10818_));
 sky130_fd_sc_hd__nand3b_1 _20961_ (.A_N(_10809_),
    .B(_10816_),
    .C(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__nor2_1 _20962_ (.A(_10802_),
    .B(_10819_),
    .Y(_10820_));
 sky130_fd_sc_hd__nand2_4 _20963_ (.A(_10725_),
    .B(_10820_),
    .Y(_10821_));
 sky130_fd_sc_hd__o21ai_1 _20964_ (.A1(_10809_),
    .A2(_10816_),
    .B1(_10808_),
    .Y(_10823_));
 sky130_fd_sc_hd__nor2_1 _20965_ (.A(_10799_),
    .B(_10773_),
    .Y(_10824_));
 sky130_fd_sc_hd__inv_2 _20966_ (.A(_10798_),
    .Y(_10825_));
 sky130_fd_sc_hd__o21ai_1 _20967_ (.A1(_10772_),
    .A2(_10825_),
    .B1(_10797_),
    .Y(_10826_));
 sky130_fd_sc_hd__a21oi_2 _20968_ (.A1(_10823_),
    .A2(_10824_),
    .B1(_10826_),
    .Y(_10827_));
 sky130_fd_sc_hd__nand2_2 _20969_ (.A(_10821_),
    .B(_10827_),
    .Y(_10828_));
 sky130_fd_sc_hd__nand2_2 _20970_ (.A(_10784_),
    .B(_10254_),
    .Y(_10829_));
 sky130_fd_sc_hd__xor2_4 _20971_ (.A(_10280_),
    .B(_10829_),
    .X(_10830_));
 sky130_fd_sc_hd__nand3_2 _20972_ (.A(_10792_),
    .B(_10683_),
    .C(_10787_),
    .Y(_10831_));
 sky130_fd_sc_hd__xor2_4 _20973_ (.A(_10830_),
    .B(_10831_),
    .X(_10832_));
 sky130_fd_sc_hd__clkinvlp_2 _20974_ (.A(_10832_),
    .Y(_10834_));
 sky130_fd_sc_hd__nand2_4 _20975_ (.A(_10828_),
    .B(_10834_),
    .Y(_10835_));
 sky130_fd_sc_hd__nand3_4 _20976_ (.A(_10821_),
    .B(_10827_),
    .C(_10832_),
    .Y(_10836_));
 sky130_fd_sc_hd__nand2_8 _20977_ (.A(_10836_),
    .B(_10835_),
    .Y(_10837_));
 sky130_fd_sc_hd__buf_8 _20978_ (.A(_10837_),
    .X(_10838_));
 sky130_fd_sc_hd__buf_6 _20979_ (.A(_10838_),
    .X(\div1i.quot[10] ));
 sky130_fd_sc_hd__nand2_1 _20980_ (.A(_10431_),
    .B(_10518_),
    .Y(_10839_));
 sky130_fd_sc_hd__inv_2 _20981_ (.A(_10522_),
    .Y(_10840_));
 sky130_fd_sc_hd__nand2_1 _20982_ (.A(_10839_),
    .B(_10840_),
    .Y(_10841_));
 sky130_fd_sc_hd__inv_2 _20983_ (.A(_10498_),
    .Y(_10842_));
 sky130_fd_sc_hd__nand2_2 _20984_ (.A(_10841_),
    .B(_10842_),
    .Y(_10844_));
 sky130_fd_sc_hd__nand2_1 _20985_ (.A(_10844_),
    .B(_10497_),
    .Y(_10845_));
 sky130_fd_sc_hd__inv_2 _20986_ (.A(_10486_),
    .Y(_10846_));
 sky130_fd_sc_hd__nand2_1 _20987_ (.A(_10845_),
    .B(_10846_),
    .Y(_10847_));
 sky130_fd_sc_hd__nand3_2 _20988_ (.A(_10844_),
    .B(_10486_),
    .C(_10497_),
    .Y(_10848_));
 sky130_fd_sc_hd__nand2_1 _20989_ (.A(_10847_),
    .B(_10848_),
    .Y(_10849_));
 sky130_fd_sc_hd__nand2_2 _20990_ (.A(_10849_),
    .B(_07226_),
    .Y(_10850_));
 sky130_fd_sc_hd__nand3_1 _20991_ (.A(_10839_),
    .B(_10498_),
    .C(_10840_),
    .Y(_10851_));
 sky130_fd_sc_hd__nand3_2 _20992_ (.A(_10844_),
    .B(_07128_),
    .C(_10851_),
    .Y(_10852_));
 sky130_fd_sc_hd__inv_2 _20993_ (.A(_10852_),
    .Y(_10853_));
 sky130_fd_sc_hd__nand3_2 _20994_ (.A(_10847_),
    .B(_07228_),
    .C(_10848_),
    .Y(_10855_));
 sky130_fd_sc_hd__nand3_1 _20995_ (.A(_10850_),
    .B(_10853_),
    .C(_10855_),
    .Y(_10856_));
 sky130_fd_sc_hd__nand2_1 _20996_ (.A(_10856_),
    .B(_10855_),
    .Y(_10857_));
 sky130_fd_sc_hd__inv_2 _20997_ (.A(_10517_),
    .Y(_10858_));
 sky130_fd_sc_hd__nand2_1 _20998_ (.A(_10431_),
    .B(_10858_),
    .Y(_10859_));
 sky130_fd_sc_hd__nand2_1 _20999_ (.A(_10859_),
    .B(_10515_),
    .Y(_10860_));
 sky130_fd_sc_hd__inv_2 _21000_ (.A(_10507_),
    .Y(_10861_));
 sky130_fd_sc_hd__nand2_1 _21001_ (.A(_10860_),
    .B(_10861_),
    .Y(_10862_));
 sky130_fd_sc_hd__nand3_1 _21002_ (.A(_10859_),
    .B(_10507_),
    .C(_10515_),
    .Y(_10863_));
 sky130_fd_sc_hd__nand2_1 _21003_ (.A(_10862_),
    .B(_10863_),
    .Y(_10864_));
 sky130_fd_sc_hd__nand2_1 _21004_ (.A(_10864_),
    .B(_07146_),
    .Y(_10866_));
 sky130_fd_sc_hd__or2_1 _21005_ (.A(_10858_),
    .B(_10431_),
    .X(_10867_));
 sky130_fd_sc_hd__nand2_1 _21006_ (.A(_10867_),
    .B(_10859_),
    .Y(_10868_));
 sky130_fd_sc_hd__inv_2 _21007_ (.A(_10868_),
    .Y(_10869_));
 sky130_fd_sc_hd__nand2_1 _21008_ (.A(_10869_),
    .B(_07157_),
    .Y(_10870_));
 sky130_fd_sc_hd__inv_2 _21009_ (.A(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__inv_2 _21010_ (.A(_10864_),
    .Y(_10872_));
 sky130_fd_sc_hd__nand2_1 _21011_ (.A(_10872_),
    .B(_07149_),
    .Y(_10873_));
 sky130_fd_sc_hd__inv_2 _21012_ (.A(_10873_),
    .Y(_10874_));
 sky130_fd_sc_hd__a21oi_1 _21013_ (.A1(_10866_),
    .A2(_10871_),
    .B1(_10874_),
    .Y(_10875_));
 sky130_fd_sc_hd__nand2_1 _21014_ (.A(_10844_),
    .B(_10851_),
    .Y(_10877_));
 sky130_fd_sc_hd__nand2_1 _21015_ (.A(_10877_),
    .B(_07130_),
    .Y(_10878_));
 sky130_fd_sc_hd__nand2_1 _21016_ (.A(_10878_),
    .B(_10852_),
    .Y(_10879_));
 sky130_fd_sc_hd__inv_2 _21017_ (.A(_10879_),
    .Y(_10880_));
 sky130_fd_sc_hd__nand3_1 _21018_ (.A(_10850_),
    .B(_10880_),
    .C(_10855_),
    .Y(_10881_));
 sky130_fd_sc_hd__nor2_1 _21019_ (.A(_10875_),
    .B(_10881_),
    .Y(_10882_));
 sky130_fd_sc_hd__nor2_1 _21020_ (.A(_10857_),
    .B(_10882_),
    .Y(_10883_));
 sky130_fd_sc_hd__inv_2 _21021_ (.A(_10881_),
    .Y(_10884_));
 sky130_fd_sc_hd__nand2_1 _21022_ (.A(_10323_),
    .B(_10326_),
    .Y(_10885_));
 sky130_fd_sc_hd__nand2_1 _21023_ (.A(_10885_),
    .B(_10328_),
    .Y(_10886_));
 sky130_fd_sc_hd__nand2_1 _21024_ (.A(_10886_),
    .B(_10330_),
    .Y(_10888_));
 sky130_fd_sc_hd__nand2_1 _21025_ (.A(_10888_),
    .B(_06982_),
    .Y(_10889_));
 sky130_fd_sc_hd__o21ai_1 _21026_ (.A1(_09215_),
    .A2(\div1i.quot[11] ),
    .B1(_09228_),
    .Y(_10890_));
 sky130_fd_sc_hd__nand3_1 _21027_ (.A(_10886_),
    .B(_06984_),
    .C(_10330_),
    .Y(_10891_));
 sky130_fd_sc_hd__inv_2 _21028_ (.A(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__a21o_1 _21029_ (.A1(_10889_),
    .A2(_10890_),
    .B1(_10892_),
    .X(_10893_));
 sky130_fd_sc_hd__nand2_1 _21030_ (.A(_10331_),
    .B(_10314_),
    .Y(_10894_));
 sky130_fd_sc_hd__nand2_1 _21031_ (.A(_10330_),
    .B(_10323_),
    .Y(_10895_));
 sky130_fd_sc_hd__xor2_2 _21032_ (.A(_10894_),
    .B(_10895_),
    .X(_10896_));
 sky130_fd_sc_hd__nand2_2 _21033_ (.A(_10896_),
    .B(_07043_),
    .Y(_10897_));
 sky130_fd_sc_hd__nand2_1 _21034_ (.A(_10893_),
    .B(_10897_),
    .Y(_10899_));
 sky130_fd_sc_hd__inv_2 _21035_ (.A(_10896_),
    .Y(_10900_));
 sky130_fd_sc_hd__nand2_1 _21036_ (.A(_10900_),
    .B(_07048_),
    .Y(_10901_));
 sky130_fd_sc_hd__nand2_1 _21037_ (.A(_10899_),
    .B(_10901_),
    .Y(_10902_));
 sky130_fd_sc_hd__nand2_1 _21038_ (.A(_10325_),
    .B(_10330_),
    .Y(_10903_));
 sky130_fd_sc_hd__nand2_1 _21039_ (.A(_10903_),
    .B(_10331_),
    .Y(_10904_));
 sky130_fd_sc_hd__nand2_1 _21040_ (.A(_10904_),
    .B(_10419_),
    .Y(_10905_));
 sky130_fd_sc_hd__nand3_2 _21041_ (.A(_10903_),
    .B(_10331_),
    .C(_10420_),
    .Y(_10906_));
 sky130_fd_sc_hd__nand2_1 _21042_ (.A(_10905_),
    .B(_10906_),
    .Y(_10907_));
 sky130_fd_sc_hd__nand2_1 _21043_ (.A(_10907_),
    .B(_07031_),
    .Y(_10908_));
 sky130_fd_sc_hd__nand3_1 _21044_ (.A(_10905_),
    .B(_07034_),
    .C(_10906_),
    .Y(_10910_));
 sky130_fd_sc_hd__nand2_1 _21045_ (.A(_10908_),
    .B(_10910_),
    .Y(_10911_));
 sky130_fd_sc_hd__inv_2 _21046_ (.A(_10911_),
    .Y(_10912_));
 sky130_fd_sc_hd__nand2_1 _21047_ (.A(_10902_),
    .B(_10912_),
    .Y(_10913_));
 sky130_fd_sc_hd__nand2_1 _21048_ (.A(_10913_),
    .B(_10910_),
    .Y(_10914_));
 sky130_fd_sc_hd__nand2_1 _21049_ (.A(_10906_),
    .B(_10417_),
    .Y(_10915_));
 sky130_fd_sc_hd__xor2_1 _21050_ (.A(_10409_),
    .B(_10915_),
    .X(_10916_));
 sky130_fd_sc_hd__nand2_1 _21051_ (.A(_10916_),
    .B(_09823_),
    .Y(_10917_));
 sky130_fd_sc_hd__nand2_1 _21052_ (.A(_10914_),
    .B(_10917_),
    .Y(_10918_));
 sky130_fd_sc_hd__or2_1 _21053_ (.A(_09823_),
    .B(_10916_),
    .X(_10919_));
 sky130_fd_sc_hd__nand2_1 _21054_ (.A(_10918_),
    .B(_10919_),
    .Y(_10921_));
 sky130_fd_sc_hd__nor2_1 _21055_ (.A(_10409_),
    .B(_10419_),
    .Y(_10922_));
 sky130_fd_sc_hd__nand3_2 _21056_ (.A(_10903_),
    .B(_10922_),
    .C(_10331_),
    .Y(_10923_));
 sky130_fd_sc_hd__inv_2 _21057_ (.A(_10425_),
    .Y(_10924_));
 sky130_fd_sc_hd__nand2_1 _21058_ (.A(_10923_),
    .B(_10924_),
    .Y(_10925_));
 sky130_fd_sc_hd__nand2_1 _21059_ (.A(_10925_),
    .B(_10397_),
    .Y(_10926_));
 sky130_fd_sc_hd__nand2_1 _21060_ (.A(_10926_),
    .B(_10394_),
    .Y(_10927_));
 sky130_fd_sc_hd__nand2_1 _21061_ (.A(_10927_),
    .B(_10387_),
    .Y(_10928_));
 sky130_fd_sc_hd__nand3_1 _21062_ (.A(_10926_),
    .B(_10386_),
    .C(_10394_),
    .Y(_10929_));
 sky130_fd_sc_hd__nand2_1 _21063_ (.A(_10928_),
    .B(_10929_),
    .Y(_10930_));
 sky130_fd_sc_hd__nand2_1 _21064_ (.A(_10930_),
    .B(_08738_),
    .Y(_10932_));
 sky130_fd_sc_hd__nand3_1 _21065_ (.A(_10923_),
    .B(_10396_),
    .C(_10924_),
    .Y(_10933_));
 sky130_fd_sc_hd__nand2_1 _21066_ (.A(_10926_),
    .B(_10933_),
    .Y(_10934_));
 sky130_fd_sc_hd__nand2_1 _21067_ (.A(_10934_),
    .B(_07024_),
    .Y(_10935_));
 sky130_fd_sc_hd__nand3_2 _21068_ (.A(_10926_),
    .B(_07021_),
    .C(_10933_),
    .Y(_10936_));
 sky130_fd_sc_hd__nand2_1 _21069_ (.A(_10935_),
    .B(_10936_),
    .Y(_10937_));
 sky130_fd_sc_hd__inv_2 _21070_ (.A(_10937_),
    .Y(_10938_));
 sky130_fd_sc_hd__buf_6 _21071_ (.A(_05896_),
    .X(_10939_));
 sky130_fd_sc_hd__nand3_1 _21072_ (.A(_10928_),
    .B(_10939_),
    .C(_10929_),
    .Y(_10940_));
 sky130_fd_sc_hd__nand3_1 _21073_ (.A(_10932_),
    .B(_10938_),
    .C(_10940_),
    .Y(_10941_));
 sky130_fd_sc_hd__inv_2 _21074_ (.A(_10941_),
    .Y(_10943_));
 sky130_fd_sc_hd__nand2_1 _21075_ (.A(_10921_),
    .B(_10943_),
    .Y(_10944_));
 sky130_fd_sc_hd__inv_2 _21076_ (.A(_10936_),
    .Y(_10945_));
 sky130_fd_sc_hd__a21boi_1 _21077_ (.A1(_10932_),
    .A2(_10945_),
    .B1_N(_10940_),
    .Y(_10946_));
 sky130_fd_sc_hd__nand2_2 _21078_ (.A(_10944_),
    .B(_10946_),
    .Y(_10947_));
 sky130_fd_sc_hd__nand2_1 _21079_ (.A(_10873_),
    .B(_10866_),
    .Y(_10948_));
 sky130_fd_sc_hd__inv_2 _21080_ (.A(_10948_),
    .Y(_10949_));
 sky130_fd_sc_hd__nand2_1 _21081_ (.A(_10868_),
    .B(_07155_),
    .Y(_10950_));
 sky130_fd_sc_hd__nand2_1 _21082_ (.A(_10870_),
    .B(_10950_),
    .Y(_10951_));
 sky130_fd_sc_hd__inv_2 _21083_ (.A(_10951_),
    .Y(_10952_));
 sky130_fd_sc_hd__nand2_1 _21084_ (.A(_10949_),
    .B(_10952_),
    .Y(_10954_));
 sky130_fd_sc_hd__inv_2 _21085_ (.A(_10954_),
    .Y(_10955_));
 sky130_fd_sc_hd__nand3_2 _21086_ (.A(_10884_),
    .B(_10947_),
    .C(_10955_),
    .Y(_10956_));
 sky130_fd_sc_hd__nand2_2 _21087_ (.A(_10883_),
    .B(_10956_),
    .Y(_10957_));
 sky130_fd_sc_hd__inv_2 _21088_ (.A(_10611_),
    .Y(_10958_));
 sky130_fd_sc_hd__inv_2 _21089_ (.A(_10620_),
    .Y(_10959_));
 sky130_fd_sc_hd__nand2_1 _21090_ (.A(_10526_),
    .B(_10959_),
    .Y(_10960_));
 sky130_fd_sc_hd__nand2_1 _21091_ (.A(_10960_),
    .B(_10619_),
    .Y(_10961_));
 sky130_fd_sc_hd__or2_1 _21092_ (.A(_10958_),
    .B(_10961_),
    .X(_10962_));
 sky130_fd_sc_hd__nand2_1 _21093_ (.A(_10961_),
    .B(_10958_),
    .Y(_10963_));
 sky130_fd_sc_hd__nand2_1 _21094_ (.A(_10962_),
    .B(_10963_),
    .Y(_10965_));
 sky130_fd_sc_hd__nand2_1 _21095_ (.A(_10965_),
    .B(_07247_),
    .Y(_10966_));
 sky130_fd_sc_hd__nand3_1 _21096_ (.A(_10962_),
    .B(_07249_),
    .C(_10963_),
    .Y(_10967_));
 sky130_fd_sc_hd__nand2_1 _21097_ (.A(_10966_),
    .B(_10967_),
    .Y(_10968_));
 sky130_fd_sc_hd__inv_2 _21098_ (.A(_10968_),
    .Y(_10969_));
 sky130_fd_sc_hd__or2_1 _21099_ (.A(_10959_),
    .B(_10526_),
    .X(_10970_));
 sky130_fd_sc_hd__nand2_1 _21100_ (.A(_10970_),
    .B(_10960_),
    .Y(_10971_));
 sky130_fd_sc_hd__inv_2 _21101_ (.A(_10971_),
    .Y(_10972_));
 sky130_fd_sc_hd__nand2_1 _21102_ (.A(_10972_),
    .B(_06521_),
    .Y(_10973_));
 sky130_fd_sc_hd__nand2_1 _21103_ (.A(_10971_),
    .B(_07677_),
    .Y(_10974_));
 sky130_fd_sc_hd__nand2_1 _21104_ (.A(_10973_),
    .B(_10974_),
    .Y(_10976_));
 sky130_fd_sc_hd__inv_2 _21105_ (.A(_10976_),
    .Y(_10977_));
 sky130_fd_sc_hd__nand2_1 _21106_ (.A(_10969_),
    .B(_10977_),
    .Y(_10978_));
 sky130_fd_sc_hd__inv_4 _21107_ (.A(_10978_),
    .Y(_10979_));
 sky130_fd_sc_hd__nand2_1 _21108_ (.A(_10957_),
    .B(_10979_),
    .Y(_10980_));
 sky130_fd_sc_hd__inv_2 _21109_ (.A(_10973_),
    .Y(_10981_));
 sky130_fd_sc_hd__a21boi_1 _21110_ (.A1(_10966_),
    .A2(_10981_),
    .B1_N(_10967_),
    .Y(_10982_));
 sky130_fd_sc_hd__nand2_1 _21111_ (.A(_10980_),
    .B(_10982_),
    .Y(_10983_));
 sky130_fd_sc_hd__nand2_1 _21112_ (.A(_10526_),
    .B(_10621_),
    .Y(_10984_));
 sky130_fd_sc_hd__inv_2 _21113_ (.A(_10626_),
    .Y(_10985_));
 sky130_fd_sc_hd__nand2_1 _21114_ (.A(_10984_),
    .B(_10985_),
    .Y(_10987_));
 sky130_fd_sc_hd__inv_2 _21115_ (.A(_10603_),
    .Y(_10988_));
 sky130_fd_sc_hd__nand2_1 _21116_ (.A(_10987_),
    .B(_10988_),
    .Y(_10989_));
 sky130_fd_sc_hd__nand3_1 _21117_ (.A(_10984_),
    .B(_10603_),
    .C(_10985_),
    .Y(_10990_));
 sky130_fd_sc_hd__nand2_1 _21118_ (.A(_10989_),
    .B(_10990_),
    .Y(_10991_));
 sky130_fd_sc_hd__inv_2 _21119_ (.A(_10991_),
    .Y(_10992_));
 sky130_fd_sc_hd__nand2_1 _21120_ (.A(_10992_),
    .B(_07278_),
    .Y(_10993_));
 sky130_fd_sc_hd__nand2_1 _21121_ (.A(_10991_),
    .B(_07276_),
    .Y(_10994_));
 sky130_fd_sc_hd__nand2_1 _21122_ (.A(_10993_),
    .B(_10994_),
    .Y(_10995_));
 sky130_fd_sc_hd__inv_2 _21123_ (.A(_10995_),
    .Y(_10996_));
 sky130_fd_sc_hd__nand2_1 _21124_ (.A(_10983_),
    .B(_10996_),
    .Y(_10998_));
 sky130_fd_sc_hd__inv_4 _21125_ (.A(_10837_),
    .Y(_10999_));
 sky130_fd_sc_hd__buf_6 _21126_ (.A(_10999_),
    .X(_11000_));
 sky130_fd_sc_hd__nand3_1 _21127_ (.A(_10980_),
    .B(_10995_),
    .C(_10982_),
    .Y(_11001_));
 sky130_fd_sc_hd__nand3_1 _21128_ (.A(_10998_),
    .B(_11000_),
    .C(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__nand2_1 _21129_ (.A(_10838_),
    .B(_10992_),
    .Y(_11003_));
 sky130_fd_sc_hd__nand2_1 _21130_ (.A(_11002_),
    .B(_11003_),
    .Y(_11004_));
 sky130_fd_sc_hd__nand2_1 _21131_ (.A(_11004_),
    .B(_06554_),
    .Y(_11005_));
 sky130_fd_sc_hd__nand3_1 _21132_ (.A(_11002_),
    .B(_06556_),
    .C(_11003_),
    .Y(_11006_));
 sky130_fd_sc_hd__nand2_1 _21133_ (.A(_11005_),
    .B(_11006_),
    .Y(_11007_));
 sky130_fd_sc_hd__nand2_1 _21134_ (.A(_10957_),
    .B(_10977_),
    .Y(_11009_));
 sky130_fd_sc_hd__nand2_1 _21135_ (.A(_11009_),
    .B(_10973_),
    .Y(_11010_));
 sky130_fd_sc_hd__nand2_1 _21136_ (.A(_11010_),
    .B(_10969_),
    .Y(_11011_));
 sky130_fd_sc_hd__nand3_1 _21137_ (.A(_11009_),
    .B(_10968_),
    .C(_10973_),
    .Y(_11012_));
 sky130_fd_sc_hd__nand2_1 _21138_ (.A(_11011_),
    .B(_11012_),
    .Y(_11013_));
 sky130_fd_sc_hd__nand2_1 _21139_ (.A(_11013_),
    .B(_11000_),
    .Y(_11014_));
 sky130_fd_sc_hd__nand2_1 _21140_ (.A(_10838_),
    .B(_10965_),
    .Y(_11015_));
 sky130_fd_sc_hd__nand2_1 _21141_ (.A(_11014_),
    .B(_11015_),
    .Y(_11016_));
 sky130_fd_sc_hd__nand2_1 _21142_ (.A(_11016_),
    .B(_06568_),
    .Y(_11017_));
 sky130_fd_sc_hd__nand3_2 _21143_ (.A(_11014_),
    .B(_06570_),
    .C(_11015_),
    .Y(_11018_));
 sky130_fd_sc_hd__nand2_1 _21144_ (.A(_11017_),
    .B(_11018_),
    .Y(_11020_));
 sky130_fd_sc_hd__nor2_1 _21145_ (.A(_11007_),
    .B(_11020_),
    .Y(_11021_));
 sky130_fd_sc_hd__nand2_1 _21146_ (.A(_10955_),
    .B(_10947_),
    .Y(_11022_));
 sky130_fd_sc_hd__nand2_1 _21147_ (.A(_11022_),
    .B(_10875_),
    .Y(_11023_));
 sky130_fd_sc_hd__nand2_1 _21148_ (.A(_11023_),
    .B(_10880_),
    .Y(_11024_));
 sky130_fd_sc_hd__nand2_1 _21149_ (.A(_11024_),
    .B(_10852_),
    .Y(_11025_));
 sky130_fd_sc_hd__nand3_1 _21150_ (.A(_11025_),
    .B(_10855_),
    .C(_10850_),
    .Y(_11026_));
 sky130_fd_sc_hd__nand2_1 _21151_ (.A(_10850_),
    .B(_10855_),
    .Y(_11027_));
 sky130_fd_sc_hd__nand3_1 _21152_ (.A(_11024_),
    .B(_10852_),
    .C(_11027_),
    .Y(_11028_));
 sky130_fd_sc_hd__nand2_1 _21153_ (.A(_11026_),
    .B(_11028_),
    .Y(_11029_));
 sky130_fd_sc_hd__nand2_1 _21154_ (.A(_11029_),
    .B(_11000_),
    .Y(_11031_));
 sky130_fd_sc_hd__nand2_1 _21155_ (.A(\div1i.quot[10] ),
    .B(_10849_),
    .Y(_11032_));
 sky130_fd_sc_hd__nand3_1 _21156_ (.A(_11031_),
    .B(_07318_),
    .C(_11032_),
    .Y(_11033_));
 sky130_fd_sc_hd__or2_1 _21157_ (.A(_10977_),
    .B(_10957_),
    .X(_11034_));
 sky130_fd_sc_hd__nand3_1 _21158_ (.A(_11034_),
    .B(_11000_),
    .C(_11009_),
    .Y(_11035_));
 sky130_fd_sc_hd__nand2_1 _21159_ (.A(_10838_),
    .B(_10972_),
    .Y(_11036_));
 sky130_fd_sc_hd__nand3_1 _21160_ (.A(_11035_),
    .B(_09944_),
    .C(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__inv_2 _21161_ (.A(_11037_),
    .Y(_11038_));
 sky130_fd_sc_hd__a21o_1 _21162_ (.A1(_11035_),
    .A2(_11036_),
    .B1(_09944_),
    .X(_11039_));
 sky130_fd_sc_hd__o21ai_1 _21163_ (.A1(_11033_),
    .A2(_11038_),
    .B1(_11039_),
    .Y(_11040_));
 sky130_fd_sc_hd__inv_2 _21164_ (.A(_11006_),
    .Y(_11042_));
 sky130_fd_sc_hd__o21ai_1 _21165_ (.A1(_11018_),
    .A2(_11042_),
    .B1(_11005_),
    .Y(_11043_));
 sky130_fd_sc_hd__a21oi_1 _21166_ (.A1(_11021_),
    .A2(_11040_),
    .B1(_11043_),
    .Y(_11044_));
 sky130_fd_sc_hd__inv_2 _21167_ (.A(_10888_),
    .Y(_11045_));
 sky130_fd_sc_hd__nand2_1 _21168_ (.A(_10837_),
    .B(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__nand2_1 _21169_ (.A(_10889_),
    .B(_10891_),
    .Y(_11047_));
 sky130_fd_sc_hd__xor2_1 _21170_ (.A(_10890_),
    .B(_11047_),
    .X(_11048_));
 sky130_fd_sc_hd__nand3b_1 _21171_ (.A_N(_11048_),
    .B(_10835_),
    .C(_10836_),
    .Y(_11049_));
 sky130_fd_sc_hd__nand2_1 _21172_ (.A(_11046_),
    .B(_11049_),
    .Y(_11050_));
 sky130_fd_sc_hd__nand2_1 _21173_ (.A(_11050_),
    .B(_08857_),
    .Y(_11051_));
 sky130_fd_sc_hd__nor2_1 _21174_ (.A(_09215_),
    .B(_10683_),
    .Y(_11053_));
 sky130_fd_sc_hd__or2_1 _21175_ (.A(_06607_),
    .B(_11053_),
    .X(_11054_));
 sky130_fd_sc_hd__nand2_1 _21176_ (.A(_11054_),
    .B(_10328_),
    .Y(_11055_));
 sky130_fd_sc_hd__inv_2 _21177_ (.A(_11055_),
    .Y(_11056_));
 sky130_fd_sc_hd__nand2_1 _21178_ (.A(_10837_),
    .B(_11056_),
    .Y(_11057_));
 sky130_fd_sc_hd__nand3_1 _21179_ (.A(_10835_),
    .B(_10836_),
    .C(_11053_),
    .Y(_11058_));
 sky130_fd_sc_hd__nand2_1 _21180_ (.A(_11057_),
    .B(_11058_),
    .Y(_11059_));
 sky130_fd_sc_hd__nand2_1 _21181_ (.A(_11059_),
    .B(_06615_),
    .Y(_11060_));
 sky130_fd_sc_hd__nand2_1 _21182_ (.A(_11051_),
    .B(_11060_),
    .Y(_11061_));
 sky130_fd_sc_hd__inv_2 _21183_ (.A(_11061_),
    .Y(_11062_));
 sky130_fd_sc_hd__nand3_1 _21184_ (.A(_11057_),
    .B(_06620_),
    .C(_11058_),
    .Y(_11064_));
 sky130_fd_sc_hd__nand3_2 _21185_ (.A(_10837_),
    .B(_09228_),
    .C(_07004_),
    .Y(_11065_));
 sky130_fd_sc_hd__inv_2 _21186_ (.A(_11065_),
    .Y(_11066_));
 sky130_fd_sc_hd__nand3_2 _21187_ (.A(_11060_),
    .B(_11064_),
    .C(_11066_),
    .Y(_11067_));
 sky130_fd_sc_hd__nand2_1 _21188_ (.A(_11062_),
    .B(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__buf_6 _21189_ (.A(_08857_),
    .X(_11069_));
 sky130_fd_sc_hd__or2_1 _21190_ (.A(_11069_),
    .B(_11050_),
    .X(_11070_));
 sky130_fd_sc_hd__nand2_1 _21191_ (.A(_11068_),
    .B(_11070_),
    .Y(_11071_));
 sky130_fd_sc_hd__inv_2 _21192_ (.A(_11071_),
    .Y(_11072_));
 sky130_fd_sc_hd__clkinvlp_2 _21193_ (.A(_10934_),
    .Y(_11073_));
 sky130_fd_sc_hd__nand2_1 _21194_ (.A(_10838_),
    .B(_11073_),
    .Y(_11075_));
 sky130_fd_sc_hd__nand2_1 _21195_ (.A(_10921_),
    .B(_10938_),
    .Y(_11076_));
 sky130_fd_sc_hd__nand3_1 _21196_ (.A(_10918_),
    .B(_10937_),
    .C(_10919_),
    .Y(_11077_));
 sky130_fd_sc_hd__nand2_1 _21197_ (.A(_11076_),
    .B(_11077_),
    .Y(_11078_));
 sky130_fd_sc_hd__inv_2 _21198_ (.A(_11078_),
    .Y(_11079_));
 sky130_fd_sc_hd__nand3_1 _21199_ (.A(_10835_),
    .B(_10836_),
    .C(_11079_),
    .Y(_11080_));
 sky130_fd_sc_hd__nand2_1 _21200_ (.A(_11075_),
    .B(_11080_),
    .Y(_11081_));
 sky130_fd_sc_hd__nand2_1 _21201_ (.A(_11081_),
    .B(_06636_),
    .Y(_11082_));
 sky130_fd_sc_hd__nand3_2 _21202_ (.A(_11075_),
    .B(_06639_),
    .C(_11080_),
    .Y(_11083_));
 sky130_fd_sc_hd__nand2_2 _21203_ (.A(_11082_),
    .B(_11083_),
    .Y(_11084_));
 sky130_fd_sc_hd__inv_2 _21204_ (.A(_11084_),
    .Y(_11086_));
 sky130_fd_sc_hd__nand2_1 _21205_ (.A(_10838_),
    .B(_10916_),
    .Y(_11087_));
 sky130_fd_sc_hd__nand2_1 _21206_ (.A(_10919_),
    .B(_10917_),
    .Y(_11088_));
 sky130_fd_sc_hd__xor2_1 _21207_ (.A(_10914_),
    .B(_11088_),
    .X(_11089_));
 sky130_fd_sc_hd__nand3_1 _21208_ (.A(_10835_),
    .B(_10836_),
    .C(_11089_),
    .Y(_11090_));
 sky130_fd_sc_hd__nand2_1 _21209_ (.A(_11087_),
    .B(_11090_),
    .Y(_11091_));
 sky130_fd_sc_hd__nand2_1 _21210_ (.A(_11091_),
    .B(_06648_),
    .Y(_11092_));
 sky130_fd_sc_hd__nand3_2 _21211_ (.A(_11087_),
    .B(_06651_),
    .C(_11090_),
    .Y(_11093_));
 sky130_fd_sc_hd__nand2_1 _21212_ (.A(_11092_),
    .B(_11093_),
    .Y(_11094_));
 sky130_fd_sc_hd__inv_2 _21213_ (.A(_11094_),
    .Y(_11095_));
 sky130_fd_sc_hd__nand2_1 _21214_ (.A(_11086_),
    .B(_11095_),
    .Y(_11097_));
 sky130_fd_sc_hd__clkinvlp_2 _21215_ (.A(_10907_),
    .Y(_11098_));
 sky130_fd_sc_hd__nand2_1 _21216_ (.A(_10838_),
    .B(_11098_),
    .Y(_11099_));
 sky130_fd_sc_hd__or2_1 _21217_ (.A(_10912_),
    .B(_10902_),
    .X(_11100_));
 sky130_fd_sc_hd__nand2_1 _21218_ (.A(_11100_),
    .B(_10913_),
    .Y(_11101_));
 sky130_fd_sc_hd__inv_2 _21219_ (.A(_11101_),
    .Y(_11102_));
 sky130_fd_sc_hd__nand3_1 _21220_ (.A(_10835_),
    .B(_10836_),
    .C(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__nand2_1 _21221_ (.A(_11099_),
    .B(_11103_),
    .Y(_11104_));
 sky130_fd_sc_hd__buf_6 _21222_ (.A(_06033_),
    .X(_11105_));
 sky130_fd_sc_hd__nand2_1 _21223_ (.A(_11104_),
    .B(_11105_),
    .Y(_11106_));
 sky130_fd_sc_hd__nand3_1 _21224_ (.A(_11099_),
    .B(_07092_),
    .C(_11103_),
    .Y(_11108_));
 sky130_fd_sc_hd__nand2_1 _21225_ (.A(_11106_),
    .B(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__inv_2 _21226_ (.A(_11109_),
    .Y(_11110_));
 sky130_fd_sc_hd__nand2_1 _21227_ (.A(_10837_),
    .B(_10900_),
    .Y(_11111_));
 sky130_fd_sc_hd__nand2_1 _21228_ (.A(_10901_),
    .B(_10897_),
    .Y(_11112_));
 sky130_fd_sc_hd__xnor2_1 _21229_ (.A(_10893_),
    .B(_11112_),
    .Y(_11113_));
 sky130_fd_sc_hd__nand3_1 _21230_ (.A(_10835_),
    .B(_10836_),
    .C(_11113_),
    .Y(_11114_));
 sky130_fd_sc_hd__nand2_1 _21231_ (.A(_11111_),
    .B(_11114_),
    .Y(_11115_));
 sky130_fd_sc_hd__nand2_1 _21232_ (.A(_11115_),
    .B(_07102_),
    .Y(_11116_));
 sky130_fd_sc_hd__buf_4 _21233_ (.A(_06046_),
    .X(_11117_));
 sky130_fd_sc_hd__nand3_1 _21234_ (.A(_11111_),
    .B(_11117_),
    .C(_11114_),
    .Y(_11119_));
 sky130_fd_sc_hd__nand2_1 _21235_ (.A(_11116_),
    .B(_11119_),
    .Y(_11120_));
 sky130_fd_sc_hd__inv_4 _21236_ (.A(_11120_),
    .Y(_11121_));
 sky130_fd_sc_hd__nand2_1 _21237_ (.A(_11110_),
    .B(_11121_),
    .Y(_11122_));
 sky130_fd_sc_hd__nor2_1 _21238_ (.A(_11097_),
    .B(_11122_),
    .Y(_11123_));
 sky130_fd_sc_hd__nand2_1 _21239_ (.A(_11072_),
    .B(_11123_),
    .Y(_11124_));
 sky130_fd_sc_hd__inv_2 _21240_ (.A(_11108_),
    .Y(_11125_));
 sky130_fd_sc_hd__o21ai_1 _21241_ (.A1(_11116_),
    .A2(_11125_),
    .B1(_11106_),
    .Y(_11126_));
 sky130_fd_sc_hd__nor2_1 _21242_ (.A(_11084_),
    .B(_11094_),
    .Y(_11127_));
 sky130_fd_sc_hd__inv_2 _21243_ (.A(_11083_),
    .Y(_11128_));
 sky130_fd_sc_hd__o21ai_1 _21244_ (.A1(_11093_),
    .A2(_11128_),
    .B1(_11082_),
    .Y(_11130_));
 sky130_fd_sc_hd__a21oi_1 _21245_ (.A1(_11126_),
    .A2(_11127_),
    .B1(_11130_),
    .Y(_11131_));
 sky130_fd_sc_hd__nand2_2 _21246_ (.A(_11124_),
    .B(_11131_),
    .Y(_11132_));
 sky130_fd_sc_hd__nand2_1 _21247_ (.A(_10947_),
    .B(_10952_),
    .Y(_11133_));
 sky130_fd_sc_hd__or2_1 _21248_ (.A(_10952_),
    .B(_10947_),
    .X(_11134_));
 sky130_fd_sc_hd__nand3_1 _21249_ (.A(_10999_),
    .B(_11133_),
    .C(_11134_),
    .Y(_11135_));
 sky130_fd_sc_hd__nand2_1 _21250_ (.A(_10838_),
    .B(_10869_),
    .Y(_11136_));
 sky130_fd_sc_hd__nand2_1 _21251_ (.A(_11135_),
    .B(_11136_),
    .Y(_11137_));
 sky130_fd_sc_hd__nand2_1 _21252_ (.A(_11137_),
    .B(_06695_),
    .Y(_11138_));
 sky130_fd_sc_hd__nand3_2 _21253_ (.A(_11135_),
    .B(_06697_),
    .C(_11136_),
    .Y(_11139_));
 sky130_fd_sc_hd__nand2_2 _21254_ (.A(_11138_),
    .B(_11139_),
    .Y(_11141_));
 sky130_fd_sc_hd__inv_2 _21255_ (.A(_11141_),
    .Y(_11142_));
 sky130_fd_sc_hd__nand2_1 _21256_ (.A(_10932_),
    .B(_10940_),
    .Y(_11143_));
 sky130_fd_sc_hd__nand2_1 _21257_ (.A(_11076_),
    .B(_10936_),
    .Y(_11144_));
 sky130_fd_sc_hd__xor2_1 _21258_ (.A(_11143_),
    .B(_11144_),
    .X(_11145_));
 sky130_fd_sc_hd__nand2_1 _21259_ (.A(_11145_),
    .B(_11000_),
    .Y(_11146_));
 sky130_fd_sc_hd__nand2_1 _21260_ (.A(_10838_),
    .B(_10930_),
    .Y(_11147_));
 sky130_fd_sc_hd__nand2_1 _21261_ (.A(_11146_),
    .B(_11147_),
    .Y(_11148_));
 sky130_fd_sc_hd__nand2_1 _21262_ (.A(_11148_),
    .B(_09410_),
    .Y(_11149_));
 sky130_fd_sc_hd__nand3_2 _21263_ (.A(_11146_),
    .B(_08951_),
    .C(_11147_),
    .Y(_11150_));
 sky130_fd_sc_hd__nand2_1 _21264_ (.A(_11149_),
    .B(_11150_),
    .Y(_11152_));
 sky130_fd_sc_hd__inv_2 _21265_ (.A(_11152_),
    .Y(_11153_));
 sky130_fd_sc_hd__nand2_1 _21266_ (.A(_11142_),
    .B(_11153_),
    .Y(_11154_));
 sky130_fd_sc_hd__nand2_1 _21267_ (.A(_11133_),
    .B(_10870_),
    .Y(_11155_));
 sky130_fd_sc_hd__nand2_1 _21268_ (.A(_11155_),
    .B(_10949_),
    .Y(_11156_));
 sky130_fd_sc_hd__nand3_1 _21269_ (.A(_11133_),
    .B(_10948_),
    .C(_10870_),
    .Y(_11157_));
 sky130_fd_sc_hd__nand2_1 _21270_ (.A(_11156_),
    .B(_11157_),
    .Y(_11158_));
 sky130_fd_sc_hd__nand2_1 _21271_ (.A(_11158_),
    .B(_11000_),
    .Y(_11159_));
 sky130_fd_sc_hd__nand2_1 _21272_ (.A(_10838_),
    .B(_10864_),
    .Y(_11160_));
 sky130_fd_sc_hd__nand2_1 _21273_ (.A(_11159_),
    .B(_11160_),
    .Y(_11161_));
 sky130_fd_sc_hd__nand2_1 _21274_ (.A(_11161_),
    .B(_06721_),
    .Y(_11163_));
 sky130_fd_sc_hd__nand3_2 _21275_ (.A(_11159_),
    .B(_06723_),
    .C(_11160_),
    .Y(_11164_));
 sky130_fd_sc_hd__nand2_1 _21276_ (.A(_11163_),
    .B(_11164_),
    .Y(_11165_));
 sky130_fd_sc_hd__or2_1 _21277_ (.A(_10877_),
    .B(_11000_),
    .X(_11166_));
 sky130_fd_sc_hd__nand3_1 _21278_ (.A(_11022_),
    .B(_10879_),
    .C(_10875_),
    .Y(_11167_));
 sky130_fd_sc_hd__nand3_1 _21279_ (.A(_11024_),
    .B(_11000_),
    .C(_11167_),
    .Y(_11168_));
 sky130_fd_sc_hd__nand2_1 _21280_ (.A(_11166_),
    .B(_11168_),
    .Y(_11169_));
 sky130_fd_sc_hd__nand2_1 _21281_ (.A(_11169_),
    .B(_06731_),
    .Y(_11170_));
 sky130_fd_sc_hd__nand3_2 _21282_ (.A(_11166_),
    .B(_11168_),
    .C(_06733_),
    .Y(_11171_));
 sky130_fd_sc_hd__nand2_2 _21283_ (.A(_11170_),
    .B(_11171_),
    .Y(_11172_));
 sky130_fd_sc_hd__nor2_1 _21284_ (.A(_11165_),
    .B(_11172_),
    .Y(_11174_));
 sky130_fd_sc_hd__and2b_1 _21285_ (.A_N(_11154_),
    .B(_11174_),
    .X(_11175_));
 sky130_fd_sc_hd__nand2_1 _21286_ (.A(_11132_),
    .B(_11175_),
    .Y(_11176_));
 sky130_fd_sc_hd__inv_2 _21287_ (.A(_11139_),
    .Y(_11177_));
 sky130_fd_sc_hd__o21ai_2 _21288_ (.A1(_11150_),
    .A2(_11177_),
    .B1(_11138_),
    .Y(_11178_));
 sky130_fd_sc_hd__inv_2 _21289_ (.A(_11171_),
    .Y(_11179_));
 sky130_fd_sc_hd__o21ai_1 _21290_ (.A1(_11164_),
    .A2(_11179_),
    .B1(_11170_),
    .Y(_11180_));
 sky130_fd_sc_hd__a21oi_1 _21291_ (.A1(_11174_),
    .A2(_11178_),
    .B1(_11180_),
    .Y(_11181_));
 sky130_fd_sc_hd__nand2_2 _21292_ (.A(_11176_),
    .B(_11181_),
    .Y(_11182_));
 sky130_fd_sc_hd__nand2_1 _21293_ (.A(_11031_),
    .B(_11032_),
    .Y(_11183_));
 sky130_fd_sc_hd__buf_6 _21294_ (.A(_06159_),
    .X(_11185_));
 sky130_fd_sc_hd__nand2_1 _21295_ (.A(_11183_),
    .B(_11185_),
    .Y(_11186_));
 sky130_fd_sc_hd__nand2_1 _21296_ (.A(_11186_),
    .B(_11033_),
    .Y(_11187_));
 sky130_fd_sc_hd__nand2_1 _21297_ (.A(_11039_),
    .B(_11037_),
    .Y(_11188_));
 sky130_fd_sc_hd__nor2_1 _21298_ (.A(_11187_),
    .B(_11188_),
    .Y(_11189_));
 sky130_fd_sc_hd__nand3_1 _21299_ (.A(_11182_),
    .B(_11021_),
    .C(_11189_),
    .Y(_11190_));
 sky130_fd_sc_hd__nand2_2 _21300_ (.A(_11044_),
    .B(_11190_),
    .Y(_11191_));
 sky130_fd_sc_hd__nand2_1 _21301_ (.A(_10716_),
    .B(_10717_),
    .Y(_11192_));
 sky130_fd_sc_hd__inv_2 _21302_ (.A(_11192_),
    .Y(_11193_));
 sky130_fd_sc_hd__or2_1 _21303_ (.A(_11193_),
    .B(_10629_),
    .X(_11194_));
 sky130_fd_sc_hd__nand2_1 _21304_ (.A(_10629_),
    .B(_11193_),
    .Y(_11196_));
 sky130_fd_sc_hd__nand2_1 _21305_ (.A(_11194_),
    .B(_11196_),
    .Y(_11197_));
 sky130_fd_sc_hd__inv_2 _21306_ (.A(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__buf_6 _21307_ (.A(_06207_),
    .X(_11199_));
 sky130_fd_sc_hd__nand2_1 _21308_ (.A(_11198_),
    .B(_11199_),
    .Y(_11200_));
 sky130_fd_sc_hd__nand2_1 _21309_ (.A(_11197_),
    .B(_08465_),
    .Y(_11201_));
 sky130_fd_sc_hd__nand2_1 _21310_ (.A(_11200_),
    .B(_11201_),
    .Y(_11202_));
 sky130_fd_sc_hd__inv_2 _21311_ (.A(_11202_),
    .Y(_11203_));
 sky130_fd_sc_hd__nand2_1 _21312_ (.A(_10989_),
    .B(_10601_),
    .Y(_11204_));
 sky130_fd_sc_hd__inv_2 _21313_ (.A(_10590_),
    .Y(_11205_));
 sky130_fd_sc_hd__nand2_1 _21314_ (.A(_11204_),
    .B(_11205_),
    .Y(_11207_));
 sky130_fd_sc_hd__nand3_1 _21315_ (.A(_10989_),
    .B(_10590_),
    .C(_10601_),
    .Y(_11208_));
 sky130_fd_sc_hd__nand2_1 _21316_ (.A(_11207_),
    .B(_11208_),
    .Y(_11209_));
 sky130_fd_sc_hd__nand2_1 _21317_ (.A(_11209_),
    .B(_07905_),
    .Y(_11210_));
 sky130_fd_sc_hd__nand3_1 _21318_ (.A(_11207_),
    .B(_06772_),
    .C(_11208_),
    .Y(_11211_));
 sky130_fd_sc_hd__nand3_1 _21319_ (.A(_10996_),
    .B(_11210_),
    .C(_11211_),
    .Y(_11212_));
 sky130_fd_sc_hd__inv_2 _21320_ (.A(_11212_),
    .Y(_11213_));
 sky130_fd_sc_hd__nand3_1 _21321_ (.A(_10957_),
    .B(_10979_),
    .C(_11213_),
    .Y(_11214_));
 sky130_fd_sc_hd__inv_2 _21322_ (.A(_11210_),
    .Y(_11215_));
 sky130_fd_sc_hd__o21ai_1 _21323_ (.A1(_10993_),
    .A2(_11215_),
    .B1(_11211_),
    .Y(_11216_));
 sky130_fd_sc_hd__nor2_1 _21324_ (.A(_10982_),
    .B(_11212_),
    .Y(_11218_));
 sky130_fd_sc_hd__nor2_1 _21325_ (.A(_11216_),
    .B(_11218_),
    .Y(_11219_));
 sky130_fd_sc_hd__nand2_2 _21326_ (.A(_11214_),
    .B(_11219_),
    .Y(_11220_));
 sky130_fd_sc_hd__or2_1 _21327_ (.A(_11203_),
    .B(_11220_),
    .X(_11221_));
 sky130_fd_sc_hd__buf_6 _21328_ (.A(_11000_),
    .X(_11222_));
 sky130_fd_sc_hd__nand2_1 _21329_ (.A(_11220_),
    .B(_11203_),
    .Y(_11223_));
 sky130_fd_sc_hd__nand3_1 _21330_ (.A(_11221_),
    .B(_11222_),
    .C(_11223_),
    .Y(_11224_));
 sky130_fd_sc_hd__nand2_1 _21331_ (.A(\div1i.quot[10] ),
    .B(_11198_),
    .Y(_11225_));
 sky130_fd_sc_hd__nand2_1 _21332_ (.A(_11224_),
    .B(_11225_),
    .Y(_11226_));
 sky130_fd_sc_hd__xor2_2 _21333_ (.A(_06754_),
    .B(_11226_),
    .X(_11227_));
 sky130_fd_sc_hd__nand2_1 _21334_ (.A(_11210_),
    .B(_11211_),
    .Y(_11229_));
 sky130_fd_sc_hd__nand2_1 _21335_ (.A(_10998_),
    .B(_10993_),
    .Y(_11230_));
 sky130_fd_sc_hd__xor2_1 _21336_ (.A(_11229_),
    .B(_11230_),
    .X(_11231_));
 sky130_fd_sc_hd__nand2_1 _21337_ (.A(_11231_),
    .B(_11000_),
    .Y(_11232_));
 sky130_fd_sc_hd__nand2_1 _21338_ (.A(\div1i.quot[10] ),
    .B(_11209_),
    .Y(_11233_));
 sky130_fd_sc_hd__nand2_1 _21339_ (.A(_11232_),
    .B(_11233_),
    .Y(_11234_));
 sky130_fd_sc_hd__nand2_1 _21340_ (.A(_11234_),
    .B(_06797_),
    .Y(_11235_));
 sky130_fd_sc_hd__nand3_1 _21341_ (.A(_11232_),
    .B(_06799_),
    .C(_11233_),
    .Y(_11236_));
 sky130_fd_sc_hd__nand2_1 _21342_ (.A(_11235_),
    .B(_11236_),
    .Y(_11237_));
 sky130_fd_sc_hd__nor2_1 _21343_ (.A(_11227_),
    .B(_11237_),
    .Y(_11238_));
 sky130_fd_sc_hd__nand2_1 _21344_ (.A(_11191_),
    .B(_11238_),
    .Y(_11240_));
 sky130_fd_sc_hd__nand2_1 _21345_ (.A(_11226_),
    .B(_10138_),
    .Y(_11241_));
 sky130_fd_sc_hd__o21a_1 _21346_ (.A1(_11236_),
    .A2(_11227_),
    .B1(_11241_),
    .X(_11242_));
 sky130_fd_sc_hd__nand2_1 _21347_ (.A(_11240_),
    .B(_11242_),
    .Y(_11243_));
 sky130_fd_sc_hd__nand2_1 _21348_ (.A(_10629_),
    .B(_10719_),
    .Y(_11244_));
 sky130_fd_sc_hd__inv_2 _21349_ (.A(_10721_),
    .Y(_11245_));
 sky130_fd_sc_hd__a21o_1 _21350_ (.A1(_11244_),
    .A2(_11245_),
    .B1(_10700_),
    .X(_11246_));
 sky130_fd_sc_hd__nand3_1 _21351_ (.A(_11244_),
    .B(_10700_),
    .C(_11245_),
    .Y(_11247_));
 sky130_fd_sc_hd__nand2_1 _21352_ (.A(_11246_),
    .B(_11247_),
    .Y(_11248_));
 sky130_fd_sc_hd__nand2_1 _21353_ (.A(_11248_),
    .B(_07948_),
    .Y(_11249_));
 sky130_fd_sc_hd__nand3_2 _21354_ (.A(_11246_),
    .B(_06819_),
    .C(_11247_),
    .Y(_11251_));
 sky130_fd_sc_hd__nand2_1 _21355_ (.A(_11249_),
    .B(_11251_),
    .Y(_11252_));
 sky130_fd_sc_hd__inv_4 _21356_ (.A(_11252_),
    .Y(_11253_));
 sky130_fd_sc_hd__nand2_1 _21357_ (.A(_11196_),
    .B(_10717_),
    .Y(_11254_));
 sky130_fd_sc_hd__xor2_2 _21358_ (.A(_10709_),
    .B(_11254_),
    .X(_11255_));
 sky130_fd_sc_hd__inv_2 _21359_ (.A(_11255_),
    .Y(_11256_));
 sky130_fd_sc_hd__nand2_1 _21360_ (.A(_11256_),
    .B(_06827_),
    .Y(_11257_));
 sky130_fd_sc_hd__nand2_1 _21361_ (.A(_11255_),
    .B(_07957_),
    .Y(_11258_));
 sky130_fd_sc_hd__nand2_1 _21362_ (.A(_11257_),
    .B(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__or2_1 _21363_ (.A(_11202_),
    .B(_11259_),
    .X(_11260_));
 sky130_fd_sc_hd__inv_4 _21364_ (.A(_11260_),
    .Y(_11262_));
 sky130_fd_sc_hd__nand2_1 _21365_ (.A(_11220_),
    .B(_11262_),
    .Y(_11263_));
 sky130_fd_sc_hd__inv_2 _21366_ (.A(_11200_),
    .Y(_11264_));
 sky130_fd_sc_hd__a21boi_1 _21367_ (.A1(_11264_),
    .A2(_11258_),
    .B1_N(_11257_),
    .Y(_11265_));
 sky130_fd_sc_hd__nand2_1 _21368_ (.A(_11263_),
    .B(_11265_),
    .Y(_11266_));
 sky130_fd_sc_hd__or2_1 _21369_ (.A(_11253_),
    .B(_11266_),
    .X(_11267_));
 sky130_fd_sc_hd__nand2_1 _21370_ (.A(_11266_),
    .B(_11253_),
    .Y(_11268_));
 sky130_fd_sc_hd__nand3_1 _21371_ (.A(_11267_),
    .B(_11222_),
    .C(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__or2_1 _21372_ (.A(_11248_),
    .B(_11222_),
    .X(_11270_));
 sky130_fd_sc_hd__nand2_1 _21373_ (.A(_11269_),
    .B(_11270_),
    .Y(_11271_));
 sky130_fd_sc_hd__xor2_2 _21374_ (.A(_06809_),
    .B(_11271_),
    .X(_11273_));
 sky130_fd_sc_hd__nand2_1 _21375_ (.A(_11223_),
    .B(_11200_),
    .Y(_11274_));
 sky130_fd_sc_hd__xor2_1 _21376_ (.A(_11259_),
    .B(_11274_),
    .X(_11275_));
 sky130_fd_sc_hd__nand2_1 _21377_ (.A(_11275_),
    .B(_11222_),
    .Y(_11276_));
 sky130_fd_sc_hd__nand2_1 _21378_ (.A(\div1i.quot[10] ),
    .B(_11255_),
    .Y(_11277_));
 sky130_fd_sc_hd__nand2_1 _21379_ (.A(_11276_),
    .B(_11277_),
    .Y(_11278_));
 sky130_fd_sc_hd__or2_1 _21380_ (.A(_10173_),
    .B(_11278_),
    .X(_11279_));
 sky130_fd_sc_hd__nand2_1 _21381_ (.A(_11278_),
    .B(_10173_),
    .Y(_11280_));
 sky130_fd_sc_hd__nand2_1 _21382_ (.A(_11279_),
    .B(_11280_),
    .Y(_11281_));
 sky130_fd_sc_hd__nor2_1 _21383_ (.A(_11273_),
    .B(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__nand2_1 _21384_ (.A(_11243_),
    .B(_11282_),
    .Y(_11284_));
 sky130_fd_sc_hd__nand2_1 _21385_ (.A(_11271_),
    .B(_06856_),
    .Y(_11285_));
 sky130_fd_sc_hd__o21a_1 _21386_ (.A1(_11279_),
    .A2(_11273_),
    .B1(_11285_),
    .X(_11286_));
 sky130_fd_sc_hd__nand2_2 _21387_ (.A(_11284_),
    .B(_11286_),
    .Y(_11287_));
 sky130_fd_sc_hd__a21o_1 _21388_ (.A1(_10816_),
    .A2(_10818_),
    .B1(_10725_),
    .X(_11288_));
 sky130_fd_sc_hd__nand3_1 _21389_ (.A(_10725_),
    .B(_10816_),
    .C(_10818_),
    .Y(_11289_));
 sky130_fd_sc_hd__nand2_1 _21390_ (.A(_11288_),
    .B(_11289_),
    .Y(_11290_));
 sky130_fd_sc_hd__or2_1 _21391_ (.A(_10749_),
    .B(_11290_),
    .X(_11291_));
 sky130_fd_sc_hd__nand2_1 _21392_ (.A(_11290_),
    .B(_10749_),
    .Y(_11292_));
 sky130_fd_sc_hd__nand2_1 _21393_ (.A(_11291_),
    .B(_11292_),
    .Y(_11293_));
 sky130_fd_sc_hd__inv_4 _21394_ (.A(_11293_),
    .Y(_11295_));
 sky130_fd_sc_hd__nand2_1 _21395_ (.A(_11246_),
    .B(_10699_),
    .Y(_11296_));
 sky130_fd_sc_hd__inv_2 _21396_ (.A(_10691_),
    .Y(_11297_));
 sky130_fd_sc_hd__nand2_1 _21397_ (.A(_11296_),
    .B(_11297_),
    .Y(_11298_));
 sky130_fd_sc_hd__nand3_1 _21398_ (.A(_11246_),
    .B(_10691_),
    .C(_10699_),
    .Y(_11299_));
 sky130_fd_sc_hd__nand2_1 _21399_ (.A(_11298_),
    .B(_11299_),
    .Y(_11300_));
 sky130_fd_sc_hd__nand2_1 _21400_ (.A(_11300_),
    .B(_08001_),
    .Y(_11301_));
 sky130_fd_sc_hd__nand3_2 _21401_ (.A(_11298_),
    .B(_06874_),
    .C(_11299_),
    .Y(_11302_));
 sky130_fd_sc_hd__nand3_1 _21402_ (.A(_11301_),
    .B(_11253_),
    .C(_11302_),
    .Y(_11303_));
 sky130_fd_sc_hd__inv_2 _21403_ (.A(_11303_),
    .Y(_11304_));
 sky130_fd_sc_hd__nand3_1 _21404_ (.A(_11220_),
    .B(_11262_),
    .C(_11304_),
    .Y(_11306_));
 sky130_fd_sc_hd__clkinvlp_2 _21405_ (.A(_11251_),
    .Y(_11307_));
 sky130_fd_sc_hd__inv_2 _21406_ (.A(_11302_),
    .Y(_11308_));
 sky130_fd_sc_hd__a21o_1 _21407_ (.A1(_11301_),
    .A2(_11307_),
    .B1(_11308_),
    .X(_11309_));
 sky130_fd_sc_hd__nor2_1 _21408_ (.A(_11265_),
    .B(_11303_),
    .Y(_11310_));
 sky130_fd_sc_hd__nor2_1 _21409_ (.A(_11309_),
    .B(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__nand2_1 _21410_ (.A(_11306_),
    .B(_11311_),
    .Y(_11312_));
 sky130_fd_sc_hd__or2_1 _21411_ (.A(_11295_),
    .B(_11312_),
    .X(_11313_));
 sky130_fd_sc_hd__nand2_1 _21412_ (.A(_11312_),
    .B(_11295_),
    .Y(_11314_));
 sky130_fd_sc_hd__nand2_1 _21413_ (.A(_11313_),
    .B(_11314_),
    .Y(_11315_));
 sky130_fd_sc_hd__nand2_1 _21414_ (.A(_11315_),
    .B(_11222_),
    .Y(_11317_));
 sky130_fd_sc_hd__nand2_1 _21415_ (.A(\div1i.quot[10] ),
    .B(_11290_),
    .Y(_11318_));
 sky130_fd_sc_hd__nand2_1 _21416_ (.A(_11317_),
    .B(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__nand2_1 _21417_ (.A(_11319_),
    .B(_08020_),
    .Y(_11320_));
 sky130_fd_sc_hd__nand3_1 _21418_ (.A(_11317_),
    .B(_09664_),
    .C(_11318_),
    .Y(_11321_));
 sky130_fd_sc_hd__nand2_2 _21419_ (.A(_11320_),
    .B(_11321_),
    .Y(_11322_));
 sky130_fd_sc_hd__inv_2 _21420_ (.A(_11322_),
    .Y(_11323_));
 sky130_fd_sc_hd__nand2_1 _21421_ (.A(_11301_),
    .B(_11302_),
    .Y(_11324_));
 sky130_fd_sc_hd__nand2_1 _21422_ (.A(_11268_),
    .B(_11251_),
    .Y(_11325_));
 sky130_fd_sc_hd__xor2_1 _21423_ (.A(_11324_),
    .B(_11325_),
    .X(_11326_));
 sky130_fd_sc_hd__nand2_1 _21424_ (.A(_11326_),
    .B(_11222_),
    .Y(_11328_));
 sky130_fd_sc_hd__nand2_1 _21425_ (.A(_11300_),
    .B(\div1i.quot[10] ),
    .Y(_11329_));
 sky130_fd_sc_hd__nand2_1 _21426_ (.A(_11328_),
    .B(_11329_),
    .Y(_11330_));
 sky130_fd_sc_hd__nand2_1 _21427_ (.A(_11330_),
    .B(_06903_),
    .Y(_11331_));
 sky130_fd_sc_hd__nand3_2 _21428_ (.A(_11328_),
    .B(_06898_),
    .C(_11329_),
    .Y(_11332_));
 sky130_fd_sc_hd__nand3_1 _21429_ (.A(_11323_),
    .B(_11331_),
    .C(_11332_),
    .Y(_11333_));
 sky130_fd_sc_hd__nand2_1 _21430_ (.A(_11289_),
    .B(_10816_),
    .Y(_11334_));
 sky130_fd_sc_hd__xor2_2 _21431_ (.A(_10809_),
    .B(_11334_),
    .X(_11335_));
 sky130_fd_sc_hd__inv_2 _21432_ (.A(_11335_),
    .Y(_11336_));
 sky130_fd_sc_hd__nand2_1 _21433_ (.A(_11336_),
    .B(_07461_),
    .Y(_11337_));
 sky130_fd_sc_hd__nand2_1 _21434_ (.A(_11335_),
    .B(_08041_),
    .Y(_11339_));
 sky130_fd_sc_hd__nand2_1 _21435_ (.A(_11337_),
    .B(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__inv_2 _21436_ (.A(_11340_),
    .Y(_11341_));
 sky130_fd_sc_hd__nand2_1 _21437_ (.A(_11341_),
    .B(_11295_),
    .Y(_11342_));
 sky130_fd_sc_hd__inv_2 _21438_ (.A(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__nand2_1 _21439_ (.A(_11312_),
    .B(_11343_),
    .Y(_11344_));
 sky130_fd_sc_hd__o21a_1 _21440_ (.A1(_11291_),
    .A2(_11340_),
    .B1(_11337_),
    .X(_11345_));
 sky130_fd_sc_hd__nand2_1 _21441_ (.A(_11344_),
    .B(_11345_),
    .Y(_11346_));
 sky130_fd_sc_hd__a21oi_1 _21442_ (.A1(_10720_),
    .A2(_10724_),
    .B1(_10819_),
    .Y(_11347_));
 sky130_fd_sc_hd__or2_1 _21443_ (.A(_10823_),
    .B(_11347_),
    .X(_11348_));
 sky130_fd_sc_hd__or2_1 _21444_ (.A(_10774_),
    .B(_11348_),
    .X(_11350_));
 sky130_fd_sc_hd__nand2_1 _21445_ (.A(_11348_),
    .B(_10774_),
    .Y(_11351_));
 sky130_fd_sc_hd__nand2_1 _21446_ (.A(_11350_),
    .B(_11351_),
    .Y(_11352_));
 sky130_fd_sc_hd__inv_2 _21447_ (.A(_11352_),
    .Y(_11353_));
 sky130_fd_sc_hd__nand2_1 _21448_ (.A(_11353_),
    .B(_06936_),
    .Y(_11354_));
 sky130_fd_sc_hd__nand2_1 _21449_ (.A(_11352_),
    .B(_08611_),
    .Y(_11355_));
 sky130_fd_sc_hd__nand2_1 _21450_ (.A(_11354_),
    .B(_11355_),
    .Y(_11356_));
 sky130_fd_sc_hd__inv_2 _21451_ (.A(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__nand2_1 _21452_ (.A(_11346_),
    .B(_11357_),
    .Y(_11358_));
 sky130_fd_sc_hd__nand3_1 _21453_ (.A(_11344_),
    .B(_11345_),
    .C(_11356_),
    .Y(_11359_));
 sky130_fd_sc_hd__nand3_1 _21454_ (.A(_11358_),
    .B(_11222_),
    .C(_11359_),
    .Y(_11361_));
 sky130_fd_sc_hd__nand2_1 _21455_ (.A(_11353_),
    .B(\div1i.quot[10] ),
    .Y(_11362_));
 sky130_fd_sc_hd__nand2_1 _21456_ (.A(_11361_),
    .B(_11362_),
    .Y(_11363_));
 sky130_fd_sc_hd__nand2_1 _21457_ (.A(_11363_),
    .B(_06947_),
    .Y(_11364_));
 sky130_fd_sc_hd__nand3_1 _21458_ (.A(_11361_),
    .B(_06949_),
    .C(_11362_),
    .Y(_11365_));
 sky130_fd_sc_hd__nand2_4 _21459_ (.A(_11364_),
    .B(_11365_),
    .Y(_11366_));
 sky130_fd_sc_hd__nand2_1 _21460_ (.A(_11314_),
    .B(_11291_),
    .Y(_11367_));
 sky130_fd_sc_hd__nand2_1 _21461_ (.A(_11367_),
    .B(_11341_),
    .Y(_11368_));
 sky130_fd_sc_hd__nand3_1 _21462_ (.A(_11314_),
    .B(_11340_),
    .C(_11291_),
    .Y(_11369_));
 sky130_fd_sc_hd__nand2_1 _21463_ (.A(_11368_),
    .B(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__nand2_1 _21464_ (.A(_11370_),
    .B(_11222_),
    .Y(_11372_));
 sky130_fd_sc_hd__nand2_1 _21465_ (.A(_11335_),
    .B(\div1i.quot[10] ),
    .Y(_11373_));
 sky130_fd_sc_hd__nand2_1 _21466_ (.A(_11372_),
    .B(_11373_),
    .Y(_11374_));
 sky130_fd_sc_hd__nand2_1 _21467_ (.A(_11374_),
    .B(_07474_),
    .Y(_11375_));
 sky130_fd_sc_hd__buf_6 _21468_ (.A(_06366_),
    .X(_11376_));
 sky130_fd_sc_hd__nand3_1 _21469_ (.A(_11372_),
    .B(_11376_),
    .C(_11373_),
    .Y(_11377_));
 sky130_fd_sc_hd__nand2_2 _21470_ (.A(_11375_),
    .B(_11377_),
    .Y(_11378_));
 sky130_fd_sc_hd__nor2_4 _21471_ (.A(_11366_),
    .B(_11378_),
    .Y(_11379_));
 sky130_fd_sc_hd__clkinvlp_2 _21472_ (.A(_11379_),
    .Y(_11380_));
 sky130_fd_sc_hd__nor2_2 _21473_ (.A(_11333_),
    .B(_11380_),
    .Y(_11381_));
 sky130_fd_sc_hd__nand2_4 _21474_ (.A(_11287_),
    .B(_11381_),
    .Y(_11383_));
 sky130_fd_sc_hd__o21ai_1 _21475_ (.A1(_11332_),
    .A2(_11322_),
    .B1(_11321_),
    .Y(_11384_));
 sky130_fd_sc_hd__o21ai_1 _21476_ (.A1(_11377_),
    .A2(_11366_),
    .B1(_11364_),
    .Y(_11385_));
 sky130_fd_sc_hd__a21oi_2 _21477_ (.A1(_11384_),
    .A2(_11379_),
    .B1(_11385_),
    .Y(_11386_));
 sky130_fd_sc_hd__nand2_4 _21478_ (.A(_11383_),
    .B(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__nand2_1 _21479_ (.A(_11351_),
    .B(_10772_),
    .Y(_11388_));
 sky130_fd_sc_hd__xor2_2 _21480_ (.A(_10799_),
    .B(_11388_),
    .X(_11389_));
 sky130_fd_sc_hd__nand3_1 _21481_ (.A(_11358_),
    .B(_11222_),
    .C(_11354_),
    .Y(_11390_));
 sky130_fd_sc_hd__xnor2_2 _21482_ (.A(_11389_),
    .B(_11390_),
    .Y(_11391_));
 sky130_fd_sc_hd__nand2_8 _21483_ (.A(_11387_),
    .B(_11391_),
    .Y(_11392_));
 sky130_fd_sc_hd__clkinvlp_2 _21484_ (.A(_11391_),
    .Y(_11394_));
 sky130_fd_sc_hd__nand3_4 _21485_ (.A(_11383_),
    .B(_11386_),
    .C(_11394_),
    .Y(_11395_));
 sky130_fd_sc_hd__nand2_8 _21486_ (.A(_11392_),
    .B(_11395_),
    .Y(_11396_));
 sky130_fd_sc_hd__buf_8 _21487_ (.A(_11396_),
    .X(_11397_));
 sky130_fd_sc_hd__buf_8 _21488_ (.A(net227),
    .X(\div1i.quot[9] ));
 sky130_fd_sc_hd__nand2_1 _21489_ (.A(_11060_),
    .B(_11064_),
    .Y(_11398_));
 sky130_fd_sc_hd__nand2_1 _21490_ (.A(_11398_),
    .B(_11065_),
    .Y(_11399_));
 sky130_fd_sc_hd__nand2_1 _21491_ (.A(_11399_),
    .B(_11067_),
    .Y(_11400_));
 sky130_fd_sc_hd__inv_2 _21492_ (.A(_11400_),
    .Y(_11401_));
 sky130_fd_sc_hd__nand2_1 _21493_ (.A(_11397_),
    .B(_11401_),
    .Y(_11402_));
 sky130_fd_sc_hd__o21ai_2 _21494_ (.A1(_09215_),
    .A2(\div1i.quot[10] ),
    .B1(_09228_),
    .Y(_11404_));
 sky130_fd_sc_hd__nand2_1 _21495_ (.A(_11400_),
    .B(_06982_),
    .Y(_11405_));
 sky130_fd_sc_hd__nand3_1 _21496_ (.A(_11399_),
    .B(_06984_),
    .C(_11067_),
    .Y(_11406_));
 sky130_fd_sc_hd__nand2_1 _21497_ (.A(_11405_),
    .B(_11406_),
    .Y(_11407_));
 sky130_fd_sc_hd__xor2_1 _21498_ (.A(_11404_),
    .B(_11407_),
    .X(_11408_));
 sky130_fd_sc_hd__nand3b_1 _21499_ (.A_N(_11408_),
    .B(_11392_),
    .C(_11395_),
    .Y(_11409_));
 sky130_fd_sc_hd__nand2_1 _21500_ (.A(_11402_),
    .B(_11409_),
    .Y(_11410_));
 sky130_fd_sc_hd__nand2_1 _21501_ (.A(_11410_),
    .B(_11069_),
    .Y(_11411_));
 sky130_fd_sc_hd__clkbuf_4 _21502_ (.A(_06607_),
    .X(_11412_));
 sky130_fd_sc_hd__nor2_1 _21503_ (.A(_09215_),
    .B(_11222_),
    .Y(_11413_));
 sky130_fd_sc_hd__or2_1 _21504_ (.A(_11412_),
    .B(_11413_),
    .X(_11415_));
 sky130_fd_sc_hd__nand2_1 _21505_ (.A(_11415_),
    .B(_11065_),
    .Y(_11416_));
 sky130_fd_sc_hd__inv_2 _21506_ (.A(_11416_),
    .Y(_11417_));
 sky130_fd_sc_hd__nand2_2 _21507_ (.A(_11397_),
    .B(_11417_),
    .Y(_11418_));
 sky130_fd_sc_hd__nand3_1 _21508_ (.A(_11392_),
    .B(_11395_),
    .C(_11413_),
    .Y(_11419_));
 sky130_fd_sc_hd__nand2_2 _21509_ (.A(_11418_),
    .B(_11419_),
    .Y(_11420_));
 sky130_fd_sc_hd__buf_6 _21510_ (.A(_06615_),
    .X(_11421_));
 sky130_fd_sc_hd__nand2_4 _21511_ (.A(_11420_),
    .B(_11421_),
    .Y(_11422_));
 sky130_fd_sc_hd__nand2_2 _21512_ (.A(_11411_),
    .B(_11422_),
    .Y(_11423_));
 sky130_fd_sc_hd__inv_2 _21513_ (.A(_11423_),
    .Y(_11424_));
 sky130_fd_sc_hd__buf_6 _21514_ (.A(_06620_),
    .X(_11426_));
 sky130_fd_sc_hd__nand3_2 _21515_ (.A(_11418_),
    .B(_11426_),
    .C(_11419_),
    .Y(_11427_));
 sky130_fd_sc_hd__nand3_2 _21516_ (.A(_11397_),
    .B(_09228_),
    .C(_07004_),
    .Y(_11428_));
 sky130_fd_sc_hd__inv_2 _21517_ (.A(_11428_),
    .Y(_11429_));
 sky130_fd_sc_hd__nand3_4 _21518_ (.A(_11422_),
    .B(_11427_),
    .C(_11429_),
    .Y(_11430_));
 sky130_fd_sc_hd__or2_4 _21519_ (.A(_11069_),
    .B(_11410_),
    .X(_11431_));
 sky130_fd_sc_hd__inv_2 _21520_ (.A(_11431_),
    .Y(_11432_));
 sky130_fd_sc_hd__a21oi_2 _21521_ (.A1(_11424_),
    .A2(_11430_),
    .B1(_11432_),
    .Y(_11433_));
 sky130_fd_sc_hd__inv_2 _21522_ (.A(_11126_),
    .Y(_11434_));
 sky130_fd_sc_hd__o21ai_1 _21523_ (.A1(_11122_),
    .A2(_11071_),
    .B1(_11434_),
    .Y(_11435_));
 sky130_fd_sc_hd__or2_1 _21524_ (.A(_11095_),
    .B(_11435_),
    .X(_11437_));
 sky130_fd_sc_hd__nand2_1 _21525_ (.A(_11435_),
    .B(_11095_),
    .Y(_11438_));
 sky130_fd_sc_hd__nand2_1 _21526_ (.A(_11437_),
    .B(_11438_),
    .Y(_11439_));
 sky130_fd_sc_hd__inv_4 _21527_ (.A(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__nand2_1 _21528_ (.A(_11396_),
    .B(_11440_),
    .Y(_11441_));
 sky130_fd_sc_hd__nand2_1 _21529_ (.A(_11440_),
    .B(_07021_),
    .Y(_11442_));
 sky130_fd_sc_hd__nand2_1 _21530_ (.A(_11439_),
    .B(_07024_),
    .Y(_11443_));
 sky130_fd_sc_hd__nand2_1 _21531_ (.A(_11442_),
    .B(_11443_),
    .Y(_11444_));
 sky130_fd_sc_hd__inv_2 _21532_ (.A(_11444_),
    .Y(_11445_));
 sky130_fd_sc_hd__nand2_1 _21533_ (.A(_11072_),
    .B(_11121_),
    .Y(_11446_));
 sky130_fd_sc_hd__nand2_1 _21534_ (.A(_11071_),
    .B(_11120_),
    .Y(_11448_));
 sky130_fd_sc_hd__nand2_1 _21535_ (.A(_11446_),
    .B(_11448_),
    .Y(_11449_));
 sky130_fd_sc_hd__nand2_1 _21536_ (.A(_11449_),
    .B(_07031_),
    .Y(_11450_));
 sky130_fd_sc_hd__nand3_1 _21537_ (.A(_11446_),
    .B(_07034_),
    .C(_11448_),
    .Y(_11451_));
 sky130_fd_sc_hd__nand2_1 _21538_ (.A(_11450_),
    .B(_11451_),
    .Y(_11452_));
 sky130_fd_sc_hd__inv_2 _21539_ (.A(_11452_),
    .Y(_11453_));
 sky130_fd_sc_hd__inv_2 _21540_ (.A(_11406_),
    .Y(_11454_));
 sky130_fd_sc_hd__a21o_1 _21541_ (.A1(_11405_),
    .A2(_11404_),
    .B1(_11454_),
    .X(_11455_));
 sky130_fd_sc_hd__nand2_1 _21542_ (.A(_11070_),
    .B(_11051_),
    .Y(_11456_));
 sky130_fd_sc_hd__nand2_1 _21543_ (.A(_11067_),
    .B(_11060_),
    .Y(_11457_));
 sky130_fd_sc_hd__xor2_2 _21544_ (.A(_11456_),
    .B(_11457_),
    .X(_11459_));
 sky130_fd_sc_hd__nand2_1 _21545_ (.A(_11459_),
    .B(_07043_),
    .Y(_11460_));
 sky130_fd_sc_hd__nand2_1 _21546_ (.A(_11455_),
    .B(_11460_),
    .Y(_11461_));
 sky130_fd_sc_hd__inv_2 _21547_ (.A(_11459_),
    .Y(_11462_));
 sky130_fd_sc_hd__nand2_1 _21548_ (.A(_11462_),
    .B(_07048_),
    .Y(_11463_));
 sky130_fd_sc_hd__nand2_1 _21549_ (.A(_11461_),
    .B(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__nand2_1 _21550_ (.A(_11453_),
    .B(_11464_),
    .Y(_11465_));
 sky130_fd_sc_hd__nand2_1 _21551_ (.A(_11465_),
    .B(_11451_),
    .Y(_11466_));
 sky130_fd_sc_hd__nand2_1 _21552_ (.A(_11446_),
    .B(_11116_),
    .Y(_11467_));
 sky130_fd_sc_hd__xor2_1 _21553_ (.A(_11109_),
    .B(_11467_),
    .X(_11468_));
 sky130_fd_sc_hd__nand2_1 _21554_ (.A(_11468_),
    .B(_09823_),
    .Y(_11470_));
 sky130_fd_sc_hd__nand2_1 _21555_ (.A(_11466_),
    .B(_11470_),
    .Y(_11471_));
 sky130_fd_sc_hd__inv_2 _21556_ (.A(_11468_),
    .Y(_11472_));
 sky130_fd_sc_hd__nand2_1 _21557_ (.A(_11472_),
    .B(_08176_),
    .Y(_11473_));
 sky130_fd_sc_hd__nand2_1 _21558_ (.A(_11471_),
    .B(_11473_),
    .Y(_11474_));
 sky130_fd_sc_hd__or2_1 _21559_ (.A(_11445_),
    .B(_11474_),
    .X(_11475_));
 sky130_fd_sc_hd__nand2_1 _21560_ (.A(_11474_),
    .B(_11445_),
    .Y(_11476_));
 sky130_fd_sc_hd__nand2_1 _21561_ (.A(_11475_),
    .B(_11476_),
    .Y(_11477_));
 sky130_fd_sc_hd__inv_2 _21562_ (.A(_11477_),
    .Y(_11478_));
 sky130_fd_sc_hd__nand3_1 _21563_ (.A(_11392_),
    .B(_11395_),
    .C(_11478_),
    .Y(_11479_));
 sky130_fd_sc_hd__nand2_1 _21564_ (.A(_11441_),
    .B(_11479_),
    .Y(_11481_));
 sky130_fd_sc_hd__buf_6 _21565_ (.A(_06636_),
    .X(_11482_));
 sky130_fd_sc_hd__nand2_1 _21566_ (.A(_11481_),
    .B(_11482_),
    .Y(_11483_));
 sky130_fd_sc_hd__buf_6 _21567_ (.A(_06639_),
    .X(_11484_));
 sky130_fd_sc_hd__nand3_1 _21568_ (.A(_11441_),
    .B(_11484_),
    .C(_11479_),
    .Y(_11485_));
 sky130_fd_sc_hd__nand2_1 _21569_ (.A(_11483_),
    .B(_11485_),
    .Y(_11486_));
 sky130_fd_sc_hd__inv_2 _21570_ (.A(_11486_),
    .Y(_11487_));
 sky130_fd_sc_hd__nand2_1 _21571_ (.A(_11396_),
    .B(_11472_),
    .Y(_11488_));
 sky130_fd_sc_hd__nand2_1 _21572_ (.A(_11473_),
    .B(_11470_),
    .Y(_11489_));
 sky130_fd_sc_hd__xnor2_1 _21573_ (.A(_11466_),
    .B(_11489_),
    .Y(_11490_));
 sky130_fd_sc_hd__nand3_1 _21574_ (.A(_11392_),
    .B(_11395_),
    .C(_11490_),
    .Y(_11492_));
 sky130_fd_sc_hd__nand2_1 _21575_ (.A(_11488_),
    .B(_11492_),
    .Y(_11493_));
 sky130_fd_sc_hd__buf_6 _21576_ (.A(_06651_),
    .X(_11494_));
 sky130_fd_sc_hd__nand2_1 _21577_ (.A(_11493_),
    .B(_11494_),
    .Y(_11495_));
 sky130_fd_sc_hd__clkbuf_8 _21578_ (.A(_06648_),
    .X(_11496_));
 sky130_fd_sc_hd__nand3_1 _21579_ (.A(_11488_),
    .B(_11496_),
    .C(_11492_),
    .Y(_11497_));
 sky130_fd_sc_hd__nand2_2 _21580_ (.A(_11495_),
    .B(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__inv_2 _21581_ (.A(_11498_),
    .Y(_11499_));
 sky130_fd_sc_hd__nand2_1 _21582_ (.A(_11487_),
    .B(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__inv_2 _21583_ (.A(_11449_),
    .Y(_11501_));
 sky130_fd_sc_hd__nand2_1 _21584_ (.A(_11396_),
    .B(_11501_),
    .Y(_11503_));
 sky130_fd_sc_hd__or2_1 _21585_ (.A(_11464_),
    .B(_11453_),
    .X(_11504_));
 sky130_fd_sc_hd__nand2_1 _21586_ (.A(_11504_),
    .B(_11465_),
    .Y(_11505_));
 sky130_fd_sc_hd__inv_2 _21587_ (.A(_11505_),
    .Y(_11506_));
 sky130_fd_sc_hd__nand3_1 _21588_ (.A(_11392_),
    .B(_11395_),
    .C(_11506_),
    .Y(_11507_));
 sky130_fd_sc_hd__nand2_1 _21589_ (.A(_11503_),
    .B(_11507_),
    .Y(_11508_));
 sky130_fd_sc_hd__nand2_1 _21590_ (.A(_11508_),
    .B(_11105_),
    .Y(_11509_));
 sky130_fd_sc_hd__nand3_1 _21591_ (.A(_11503_),
    .B(_07092_),
    .C(_11507_),
    .Y(_11510_));
 sky130_fd_sc_hd__nand2_2 _21592_ (.A(_11509_),
    .B(_11510_),
    .Y(_11511_));
 sky130_fd_sc_hd__inv_2 _21593_ (.A(_11511_),
    .Y(_11512_));
 sky130_fd_sc_hd__nand2_1 _21594_ (.A(_11396_),
    .B(_11462_),
    .Y(_11514_));
 sky130_fd_sc_hd__nand2_1 _21595_ (.A(_11463_),
    .B(_11460_),
    .Y(_11515_));
 sky130_fd_sc_hd__xnor2_1 _21596_ (.A(_11455_),
    .B(_11515_),
    .Y(_11516_));
 sky130_fd_sc_hd__nand3_1 _21597_ (.A(_11392_),
    .B(_11395_),
    .C(_11516_),
    .Y(_11517_));
 sky130_fd_sc_hd__nand2_1 _21598_ (.A(_11514_),
    .B(_11517_),
    .Y(_11518_));
 sky130_fd_sc_hd__nand2_2 _21599_ (.A(_11518_),
    .B(_07102_),
    .Y(_11519_));
 sky130_fd_sc_hd__nand3_1 _21600_ (.A(_11514_),
    .B(_11117_),
    .C(_11517_),
    .Y(_11520_));
 sky130_fd_sc_hd__nand2_2 _21601_ (.A(_11519_),
    .B(_11520_),
    .Y(_11521_));
 sky130_fd_sc_hd__clkinvlp_2 _21602_ (.A(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__nand2_1 _21603_ (.A(_11512_),
    .B(_11522_),
    .Y(_11523_));
 sky130_fd_sc_hd__nor2_1 _21604_ (.A(_11500_),
    .B(_11523_),
    .Y(_11525_));
 sky130_fd_sc_hd__nand2_1 _21605_ (.A(_11433_),
    .B(_11525_),
    .Y(_11526_));
 sky130_fd_sc_hd__inv_2 _21606_ (.A(_11510_),
    .Y(_11527_));
 sky130_fd_sc_hd__o21ai_2 _21607_ (.A1(_11519_),
    .A2(_11527_),
    .B1(_11509_),
    .Y(_11528_));
 sky130_fd_sc_hd__nor2_1 _21608_ (.A(_11486_),
    .B(_11498_),
    .Y(_11529_));
 sky130_fd_sc_hd__inv_2 _21609_ (.A(_11485_),
    .Y(_11530_));
 sky130_fd_sc_hd__o21ai_1 _21610_ (.A1(_11495_),
    .A2(_11530_),
    .B1(_11483_),
    .Y(_11531_));
 sky130_fd_sc_hd__a21oi_1 _21611_ (.A1(_11528_),
    .A2(_11529_),
    .B1(_11531_),
    .Y(_11532_));
 sky130_fd_sc_hd__nand2_2 _21612_ (.A(_11526_),
    .B(_11532_),
    .Y(_11533_));
 sky130_fd_sc_hd__inv_2 _21613_ (.A(_11154_),
    .Y(_11534_));
 sky130_fd_sc_hd__nand2_1 _21614_ (.A(_11132_),
    .B(_11534_),
    .Y(_11536_));
 sky130_fd_sc_hd__inv_2 _21615_ (.A(_11178_),
    .Y(_11537_));
 sky130_fd_sc_hd__nand2_1 _21616_ (.A(_11536_),
    .B(_11537_),
    .Y(_11538_));
 sky130_fd_sc_hd__inv_2 _21617_ (.A(_11165_),
    .Y(_11539_));
 sky130_fd_sc_hd__nand2_1 _21618_ (.A(_11538_),
    .B(_11539_),
    .Y(_11540_));
 sky130_fd_sc_hd__nand3_1 _21619_ (.A(_11536_),
    .B(_11165_),
    .C(_11537_),
    .Y(_11541_));
 sky130_fd_sc_hd__nand2_1 _21620_ (.A(_11540_),
    .B(_11541_),
    .Y(_11542_));
 sky130_fd_sc_hd__inv_4 _21621_ (.A(_11542_),
    .Y(_11543_));
 sky130_fd_sc_hd__nand2_1 _21622_ (.A(_11543_),
    .B(_07128_),
    .Y(_11544_));
 sky130_fd_sc_hd__nand2_1 _21623_ (.A(_11542_),
    .B(_07130_),
    .Y(_11545_));
 sky130_fd_sc_hd__nand2_1 _21624_ (.A(_11544_),
    .B(_11545_),
    .Y(_11547_));
 sky130_fd_sc_hd__inv_2 _21625_ (.A(_11547_),
    .Y(_11548_));
 sky130_fd_sc_hd__nand2_1 _21626_ (.A(_11438_),
    .B(_11093_),
    .Y(_11549_));
 sky130_fd_sc_hd__nand2_1 _21627_ (.A(_11549_),
    .B(_11086_),
    .Y(_11550_));
 sky130_fd_sc_hd__nand3_1 _21628_ (.A(_11438_),
    .B(_11084_),
    .C(_11093_),
    .Y(_11551_));
 sky130_fd_sc_hd__nand2_1 _21629_ (.A(_11550_),
    .B(_11551_),
    .Y(_11552_));
 sky130_fd_sc_hd__or2_1 _21630_ (.A(_08738_),
    .B(_11552_),
    .X(_11553_));
 sky130_fd_sc_hd__nand2_1 _21631_ (.A(_11553_),
    .B(_11442_),
    .Y(_11554_));
 sky130_fd_sc_hd__inv_2 _21632_ (.A(_11554_),
    .Y(_11555_));
 sky130_fd_sc_hd__nand2_1 _21633_ (.A(_11476_),
    .B(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__nand2_2 _21634_ (.A(_11132_),
    .B(_11153_),
    .Y(_11558_));
 sky130_fd_sc_hd__nand2_2 _21635_ (.A(_11558_),
    .B(_11150_),
    .Y(_11559_));
 sky130_fd_sc_hd__xor2_2 _21636_ (.A(_11141_),
    .B(_11559_),
    .X(_11560_));
 sky130_fd_sc_hd__nand2_2 _21637_ (.A(_11560_),
    .B(_07146_),
    .Y(_11561_));
 sky130_fd_sc_hd__or2_1 _21638_ (.A(_11142_),
    .B(_11559_),
    .X(_11562_));
 sky130_fd_sc_hd__nand2_1 _21639_ (.A(_11559_),
    .B(_11142_),
    .Y(_11563_));
 sky130_fd_sc_hd__nand3_2 _21640_ (.A(_11562_),
    .B(_07149_),
    .C(_11563_),
    .Y(_11564_));
 sky130_fd_sc_hd__or2_1 _21641_ (.A(_11153_),
    .B(_11132_),
    .X(_11565_));
 sky130_fd_sc_hd__nand2_1 _21642_ (.A(_11565_),
    .B(_11558_),
    .Y(_11566_));
 sky130_fd_sc_hd__nand2_1 _21643_ (.A(_11566_),
    .B(_07155_),
    .Y(_11567_));
 sky130_fd_sc_hd__nand3_2 _21644_ (.A(_11565_),
    .B(_07157_),
    .C(_11558_),
    .Y(_11569_));
 sky130_fd_sc_hd__nand2_1 _21645_ (.A(_11567_),
    .B(_11569_),
    .Y(_11570_));
 sky130_fd_sc_hd__inv_2 _21646_ (.A(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__nand3_1 _21647_ (.A(_11561_),
    .B(_11564_),
    .C(_11571_),
    .Y(_11572_));
 sky130_fd_sc_hd__inv_2 _21648_ (.A(_11572_),
    .Y(_11573_));
 sky130_fd_sc_hd__nand2_1 _21649_ (.A(_11552_),
    .B(_08738_),
    .Y(_11574_));
 sky130_fd_sc_hd__nand3_2 _21650_ (.A(_11556_),
    .B(_11573_),
    .C(_11574_),
    .Y(_11575_));
 sky130_fd_sc_hd__clkinvlp_2 _21651_ (.A(_11569_),
    .Y(_11576_));
 sky130_fd_sc_hd__a21boi_2 _21652_ (.A1(_11561_),
    .A2(_11576_),
    .B1_N(_11564_),
    .Y(_11577_));
 sky130_fd_sc_hd__nand2_1 _21653_ (.A(_11575_),
    .B(_11577_),
    .Y(_11578_));
 sky130_fd_sc_hd__or2_1 _21654_ (.A(_11548_),
    .B(_11578_),
    .X(_11580_));
 sky130_fd_sc_hd__inv_6 _21655_ (.A(_11396_),
    .Y(_11581_));
 sky130_fd_sc_hd__nand2_1 _21656_ (.A(_11578_),
    .B(_11548_),
    .Y(_11582_));
 sky130_fd_sc_hd__nand3_1 _21657_ (.A(_11580_),
    .B(_11581_),
    .C(_11582_),
    .Y(_11583_));
 sky130_fd_sc_hd__nand2_1 _21658_ (.A(net227),
    .B(_11543_),
    .Y(_11584_));
 sky130_fd_sc_hd__nand2_1 _21659_ (.A(_11583_),
    .B(_11584_),
    .Y(_11585_));
 sky130_fd_sc_hd__buf_6 _21660_ (.A(_06731_),
    .X(_11586_));
 sky130_fd_sc_hd__nand2_1 _21661_ (.A(_11585_),
    .B(_11586_),
    .Y(_11587_));
 sky130_fd_sc_hd__buf_6 _21662_ (.A(_06733_),
    .X(_11588_));
 sky130_fd_sc_hd__nand3_1 _21663_ (.A(_11583_),
    .B(_11588_),
    .C(_11584_),
    .Y(_11589_));
 sky130_fd_sc_hd__nand2_2 _21664_ (.A(_11587_),
    .B(_11589_),
    .Y(_11591_));
 sky130_fd_sc_hd__nand3_1 _21665_ (.A(_11556_),
    .B(_11574_),
    .C(_11571_),
    .Y(_11592_));
 sky130_fd_sc_hd__nand2_1 _21666_ (.A(_11592_),
    .B(_11569_),
    .Y(_11593_));
 sky130_fd_sc_hd__nand3_1 _21667_ (.A(_11593_),
    .B(_11564_),
    .C(_11561_),
    .Y(_11594_));
 sky130_fd_sc_hd__nand2_1 _21668_ (.A(_11561_),
    .B(_11564_),
    .Y(_11595_));
 sky130_fd_sc_hd__nand3_1 _21669_ (.A(_11592_),
    .B(_11595_),
    .C(_11569_),
    .Y(_11596_));
 sky130_fd_sc_hd__a21o_1 _21670_ (.A1(_11594_),
    .A2(_11596_),
    .B1(_11397_),
    .X(_11597_));
 sky130_fd_sc_hd__nand2_2 _21671_ (.A(net227),
    .B(_11560_),
    .Y(_11598_));
 sky130_fd_sc_hd__nand2_1 _21672_ (.A(_11597_),
    .B(_11598_),
    .Y(_11599_));
 sky130_fd_sc_hd__buf_6 _21673_ (.A(_06721_),
    .X(_11600_));
 sky130_fd_sc_hd__nand2_1 _21674_ (.A(_11599_),
    .B(_11600_),
    .Y(_11602_));
 sky130_fd_sc_hd__clkbuf_8 _21675_ (.A(_06723_),
    .X(_11603_));
 sky130_fd_sc_hd__nand3_2 _21676_ (.A(_11597_),
    .B(_11603_),
    .C(_11598_),
    .Y(_11604_));
 sky130_fd_sc_hd__nand2_2 _21677_ (.A(_11602_),
    .B(_11604_),
    .Y(_11605_));
 sky130_fd_sc_hd__nor2_2 _21678_ (.A(_11591_),
    .B(_11605_),
    .Y(_11606_));
 sky130_fd_sc_hd__a21o_1 _21679_ (.A1(_11392_),
    .A2(_11395_),
    .B1(_11566_),
    .X(_11607_));
 sky130_fd_sc_hd__a21o_1 _21680_ (.A1(_11556_),
    .A2(_11574_),
    .B1(_11571_),
    .X(_11608_));
 sky130_fd_sc_hd__nand2_1 _21681_ (.A(_11608_),
    .B(_11592_),
    .Y(_11609_));
 sky130_fd_sc_hd__inv_2 _21682_ (.A(_11609_),
    .Y(_11610_));
 sky130_fd_sc_hd__nand2_1 _21683_ (.A(_11581_),
    .B(_11610_),
    .Y(_11611_));
 sky130_fd_sc_hd__nand2_1 _21684_ (.A(_11607_),
    .B(_11611_),
    .Y(_11613_));
 sky130_fd_sc_hd__buf_6 _21685_ (.A(_06695_),
    .X(_11614_));
 sky130_fd_sc_hd__nand2_1 _21686_ (.A(_11613_),
    .B(_11614_),
    .Y(_11615_));
 sky130_fd_sc_hd__buf_6 _21687_ (.A(_06697_),
    .X(_11616_));
 sky130_fd_sc_hd__nand3_1 _21688_ (.A(_11607_),
    .B(_11611_),
    .C(_11616_),
    .Y(_11617_));
 sky130_fd_sc_hd__nand2_2 _21689_ (.A(_11615_),
    .B(_11617_),
    .Y(_11618_));
 sky130_fd_sc_hd__nand2_1 _21690_ (.A(_11553_),
    .B(_11574_),
    .Y(_11619_));
 sky130_fd_sc_hd__nand2_1 _21691_ (.A(_11476_),
    .B(_11442_),
    .Y(_11620_));
 sky130_fd_sc_hd__xor2_1 _21692_ (.A(_11619_),
    .B(_11620_),
    .X(_11621_));
 sky130_fd_sc_hd__nand2_1 _21693_ (.A(_11581_),
    .B(_11621_),
    .Y(_11622_));
 sky130_fd_sc_hd__nand2_1 _21694_ (.A(_11397_),
    .B(_11552_),
    .Y(_11624_));
 sky130_fd_sc_hd__nand2_1 _21695_ (.A(_11622_),
    .B(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__nand2b_2 _21696_ (.A_N(_11625_),
    .B(_08951_),
    .Y(_11626_));
 sky130_fd_sc_hd__nand2_1 _21697_ (.A(_11625_),
    .B(_09410_),
    .Y(_11627_));
 sky130_fd_sc_hd__nand2_1 _21698_ (.A(_11626_),
    .B(_11627_),
    .Y(_11628_));
 sky130_fd_sc_hd__nor2_1 _21699_ (.A(_11618_),
    .B(_11628_),
    .Y(_11629_));
 sky130_fd_sc_hd__nand2_1 _21700_ (.A(_11606_),
    .B(_11629_),
    .Y(_11630_));
 sky130_fd_sc_hd__inv_2 _21701_ (.A(_11630_),
    .Y(_11631_));
 sky130_fd_sc_hd__nand2_1 _21702_ (.A(_11533_),
    .B(_11631_),
    .Y(_11632_));
 sky130_fd_sc_hd__o21ai_2 _21703_ (.A1(_11626_),
    .A2(_11618_),
    .B1(_11615_),
    .Y(_11633_));
 sky130_fd_sc_hd__o21ai_1 _21704_ (.A1(_11604_),
    .A2(_11591_),
    .B1(_11587_),
    .Y(_11635_));
 sky130_fd_sc_hd__a21oi_1 _21705_ (.A1(_11606_),
    .A2(_11633_),
    .B1(_11635_),
    .Y(_11636_));
 sky130_fd_sc_hd__nand2_2 _21706_ (.A(_11636_),
    .B(_11632_),
    .Y(_11637_));
 sky130_fd_sc_hd__inv_2 _21707_ (.A(_11575_),
    .Y(_11638_));
 sky130_fd_sc_hd__nand2_1 _21708_ (.A(_11540_),
    .B(_11164_),
    .Y(_11639_));
 sky130_fd_sc_hd__clkinvlp_2 _21709_ (.A(_11172_),
    .Y(_11640_));
 sky130_fd_sc_hd__nand2_1 _21710_ (.A(_11639_),
    .B(_11640_),
    .Y(_11641_));
 sky130_fd_sc_hd__nand3_1 _21711_ (.A(_11540_),
    .B(_11172_),
    .C(_11164_),
    .Y(_11642_));
 sky130_fd_sc_hd__nand2_1 _21712_ (.A(_11641_),
    .B(_11642_),
    .Y(_11643_));
 sky130_fd_sc_hd__nand2_1 _21713_ (.A(_11643_),
    .B(_07226_),
    .Y(_11644_));
 sky130_fd_sc_hd__nand3_1 _21714_ (.A(_11641_),
    .B(_07228_),
    .C(_11642_),
    .Y(_11646_));
 sky130_fd_sc_hd__nand3_1 _21715_ (.A(_11548_),
    .B(_11644_),
    .C(_11646_),
    .Y(_11647_));
 sky130_fd_sc_hd__inv_2 _21716_ (.A(_11647_),
    .Y(_11648_));
 sky130_fd_sc_hd__nand2_1 _21717_ (.A(_11638_),
    .B(_11648_),
    .Y(_11649_));
 sky130_fd_sc_hd__nor2_1 _21718_ (.A(_11577_),
    .B(_11647_),
    .Y(_11650_));
 sky130_fd_sc_hd__nand2_1 _21719_ (.A(_11644_),
    .B(_11646_),
    .Y(_11651_));
 sky130_fd_sc_hd__o21ai_1 _21720_ (.A1(_11544_),
    .A2(_11651_),
    .B1(_11646_),
    .Y(_11652_));
 sky130_fd_sc_hd__nor2_1 _21721_ (.A(_11650_),
    .B(_11652_),
    .Y(_11653_));
 sky130_fd_sc_hd__nand2_1 _21722_ (.A(_11649_),
    .B(_11653_),
    .Y(_11654_));
 sky130_fd_sc_hd__inv_2 _21723_ (.A(_11188_),
    .Y(_11655_));
 sky130_fd_sc_hd__inv_2 _21724_ (.A(_11187_),
    .Y(_11657_));
 sky130_fd_sc_hd__nand2_1 _21725_ (.A(_11182_),
    .B(_11657_),
    .Y(_11658_));
 sky130_fd_sc_hd__nand2_1 _21726_ (.A(_11658_),
    .B(_11033_),
    .Y(_11659_));
 sky130_fd_sc_hd__or2_1 _21727_ (.A(_11655_),
    .B(_11659_),
    .X(_11660_));
 sky130_fd_sc_hd__nand2_1 _21728_ (.A(_11659_),
    .B(_11655_),
    .Y(_11661_));
 sky130_fd_sc_hd__nand2_1 _21729_ (.A(_11660_),
    .B(_11661_),
    .Y(_11662_));
 sky130_fd_sc_hd__nand2_1 _21730_ (.A(_11662_),
    .B(_07247_),
    .Y(_11663_));
 sky130_fd_sc_hd__nand3_1 _21731_ (.A(_11660_),
    .B(_07249_),
    .C(_11661_),
    .Y(_11664_));
 sky130_fd_sc_hd__nand2_1 _21732_ (.A(_11663_),
    .B(_11664_),
    .Y(_11665_));
 sky130_fd_sc_hd__inv_2 _21733_ (.A(_11665_),
    .Y(_11666_));
 sky130_fd_sc_hd__or2_1 _21734_ (.A(_11657_),
    .B(_11182_),
    .X(_11668_));
 sky130_fd_sc_hd__nand2_1 _21735_ (.A(_11668_),
    .B(_11658_),
    .Y(_11669_));
 sky130_fd_sc_hd__inv_4 _21736_ (.A(_11669_),
    .Y(_11670_));
 sky130_fd_sc_hd__buf_6 _21737_ (.A(_06521_),
    .X(_11671_));
 sky130_fd_sc_hd__nand2_1 _21738_ (.A(_11670_),
    .B(_11671_),
    .Y(_11672_));
 sky130_fd_sc_hd__nand2_1 _21739_ (.A(_11669_),
    .B(_07677_),
    .Y(_11673_));
 sky130_fd_sc_hd__nand2_1 _21740_ (.A(_11672_),
    .B(_11673_),
    .Y(_11674_));
 sky130_fd_sc_hd__inv_2 _21741_ (.A(_11674_),
    .Y(_11675_));
 sky130_fd_sc_hd__nand2_1 _21742_ (.A(_11666_),
    .B(_11675_),
    .Y(_11676_));
 sky130_fd_sc_hd__inv_2 _21743_ (.A(_11676_),
    .Y(_11677_));
 sky130_fd_sc_hd__nand2_1 _21744_ (.A(_11654_),
    .B(_11677_),
    .Y(_11679_));
 sky130_fd_sc_hd__inv_2 _21745_ (.A(_11672_),
    .Y(_11680_));
 sky130_fd_sc_hd__a21boi_2 _21746_ (.A1(_11663_),
    .A2(_11680_),
    .B1_N(_11664_),
    .Y(_11681_));
 sky130_fd_sc_hd__nand2_1 _21747_ (.A(_11679_),
    .B(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__nand2_1 _21748_ (.A(_11182_),
    .B(_11189_),
    .Y(_11683_));
 sky130_fd_sc_hd__inv_2 _21749_ (.A(_11040_),
    .Y(_11684_));
 sky130_fd_sc_hd__nand2_1 _21750_ (.A(_11683_),
    .B(_11684_),
    .Y(_11685_));
 sky130_fd_sc_hd__inv_2 _21751_ (.A(_11020_),
    .Y(_11686_));
 sky130_fd_sc_hd__nand2_1 _21752_ (.A(_11685_),
    .B(_11686_),
    .Y(_11687_));
 sky130_fd_sc_hd__nand3_1 _21753_ (.A(_11683_),
    .B(_11684_),
    .C(_11020_),
    .Y(_11688_));
 sky130_fd_sc_hd__nand2_1 _21754_ (.A(_11687_),
    .B(_11688_),
    .Y(_11690_));
 sky130_fd_sc_hd__nand2_1 _21755_ (.A(_11690_),
    .B(_07276_),
    .Y(_11691_));
 sky130_fd_sc_hd__nand3_1 _21756_ (.A(_11687_),
    .B(_11688_),
    .C(_07278_),
    .Y(_11692_));
 sky130_fd_sc_hd__nand2_1 _21757_ (.A(_11691_),
    .B(_11692_),
    .Y(_11693_));
 sky130_fd_sc_hd__inv_2 _21758_ (.A(_11693_),
    .Y(_11694_));
 sky130_fd_sc_hd__nand2_1 _21759_ (.A(_11682_),
    .B(_11694_),
    .Y(_11695_));
 sky130_fd_sc_hd__nand3_1 _21760_ (.A(_11679_),
    .B(_11693_),
    .C(_11681_),
    .Y(_11696_));
 sky130_fd_sc_hd__nand3_1 _21761_ (.A(_11695_),
    .B(_11581_),
    .C(_11696_),
    .Y(_11697_));
 sky130_fd_sc_hd__or2_1 _21762_ (.A(_11690_),
    .B(_11581_),
    .X(_11698_));
 sky130_fd_sc_hd__nand2_1 _21763_ (.A(_11697_),
    .B(_11698_),
    .Y(_11699_));
 sky130_fd_sc_hd__buf_6 _21764_ (.A(_06554_),
    .X(_11701_));
 sky130_fd_sc_hd__nand2_1 _21765_ (.A(_11699_),
    .B(_11701_),
    .Y(_11702_));
 sky130_fd_sc_hd__buf_6 _21766_ (.A(_06556_),
    .X(_11703_));
 sky130_fd_sc_hd__nand3_1 _21767_ (.A(_11697_),
    .B(_11703_),
    .C(_11698_),
    .Y(_11704_));
 sky130_fd_sc_hd__nand2_1 _21768_ (.A(_11702_),
    .B(_11704_),
    .Y(_11705_));
 sky130_fd_sc_hd__nand2_1 _21769_ (.A(_11654_),
    .B(_11675_),
    .Y(_11706_));
 sky130_fd_sc_hd__nand2_1 _21770_ (.A(_11706_),
    .B(_11672_),
    .Y(_11707_));
 sky130_fd_sc_hd__nand2_1 _21771_ (.A(_11707_),
    .B(_11666_),
    .Y(_11708_));
 sky130_fd_sc_hd__nand3_1 _21772_ (.A(_11706_),
    .B(_11665_),
    .C(_11672_),
    .Y(_11709_));
 sky130_fd_sc_hd__nand2_1 _21773_ (.A(_11708_),
    .B(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__nand2_1 _21774_ (.A(_11710_),
    .B(_11581_),
    .Y(_11712_));
 sky130_fd_sc_hd__nand2_1 _21775_ (.A(\div1i.quot[9] ),
    .B(_11662_),
    .Y(_11713_));
 sky130_fd_sc_hd__nand2_1 _21776_ (.A(_11712_),
    .B(_11713_),
    .Y(_11714_));
 sky130_fd_sc_hd__buf_6 _21777_ (.A(_06568_),
    .X(_11715_));
 sky130_fd_sc_hd__nand2_1 _21778_ (.A(_11714_),
    .B(_11715_),
    .Y(_11716_));
 sky130_fd_sc_hd__clkbuf_8 _21779_ (.A(_06570_),
    .X(_11717_));
 sky130_fd_sc_hd__nand3_2 _21780_ (.A(_11712_),
    .B(_11717_),
    .C(_11713_),
    .Y(_11718_));
 sky130_fd_sc_hd__nand2_2 _21781_ (.A(_11716_),
    .B(_11718_),
    .Y(_11719_));
 sky130_fd_sc_hd__nor2_2 _21782_ (.A(_11705_),
    .B(_11719_),
    .Y(_11720_));
 sky130_fd_sc_hd__or2_1 _21783_ (.A(_11675_),
    .B(_11654_),
    .X(_11721_));
 sky130_fd_sc_hd__nand3_1 _21784_ (.A(_11721_),
    .B(_11581_),
    .C(_11706_),
    .Y(_11723_));
 sky130_fd_sc_hd__nand2_1 _21785_ (.A(net227),
    .B(_11670_),
    .Y(_11724_));
 sky130_fd_sc_hd__nand2_1 _21786_ (.A(_11723_),
    .B(_11724_),
    .Y(_11725_));
 sky130_fd_sc_hd__nand2_1 _21787_ (.A(_11725_),
    .B(_06149_),
    .Y(_11726_));
 sky130_fd_sc_hd__nand3_1 _21788_ (.A(_11723_),
    .B(_09944_),
    .C(_11724_),
    .Y(_11727_));
 sky130_fd_sc_hd__nand2_1 _21789_ (.A(_11726_),
    .B(_11727_),
    .Y(_11728_));
 sky130_fd_sc_hd__nand2_1 _21790_ (.A(_11582_),
    .B(_11544_),
    .Y(_11729_));
 sky130_fd_sc_hd__xor2_1 _21791_ (.A(_11651_),
    .B(_11729_),
    .X(_11730_));
 sky130_fd_sc_hd__buf_6 _21792_ (.A(_11581_),
    .X(_11731_));
 sky130_fd_sc_hd__nand2_1 _21793_ (.A(_11730_),
    .B(_11731_),
    .Y(_11732_));
 sky130_fd_sc_hd__nand2_1 _21794_ (.A(\div1i.quot[9] ),
    .B(_11643_),
    .Y(_11734_));
 sky130_fd_sc_hd__nand2_1 _21795_ (.A(_11732_),
    .B(_11734_),
    .Y(_11735_));
 sky130_fd_sc_hd__nand2_1 _21796_ (.A(_11735_),
    .B(_11185_),
    .Y(_11736_));
 sky130_fd_sc_hd__nand3_1 _21797_ (.A(_11732_),
    .B(_07318_),
    .C(_11734_),
    .Y(_11737_));
 sky130_fd_sc_hd__nand2_1 _21798_ (.A(_11736_),
    .B(_11737_),
    .Y(_11738_));
 sky130_fd_sc_hd__nor2_2 _21799_ (.A(_11728_),
    .B(_11738_),
    .Y(_11739_));
 sky130_fd_sc_hd__nand2_1 _21800_ (.A(_11720_),
    .B(_11739_),
    .Y(_11740_));
 sky130_fd_sc_hd__inv_2 _21801_ (.A(_11740_),
    .Y(_11741_));
 sky130_fd_sc_hd__nand2_2 _21802_ (.A(_11637_),
    .B(_11741_),
    .Y(_11742_));
 sky130_fd_sc_hd__o21ai_1 _21803_ (.A1(_11737_),
    .A2(_11728_),
    .B1(_11726_),
    .Y(_11743_));
 sky130_fd_sc_hd__o21ai_1 _21804_ (.A1(_11718_),
    .A2(_11705_),
    .B1(_11702_),
    .Y(_11745_));
 sky130_fd_sc_hd__a21oi_2 _21805_ (.A1(_11720_),
    .A2(_11743_),
    .B1(_11745_),
    .Y(_11746_));
 sky130_fd_sc_hd__nand2_4 _21806_ (.A(_11742_),
    .B(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__nand2_1 _21807_ (.A(_11687_),
    .B(_11018_),
    .Y(_11748_));
 sky130_fd_sc_hd__inv_2 _21808_ (.A(_11007_),
    .Y(_11749_));
 sky130_fd_sc_hd__nand2_1 _21809_ (.A(_11748_),
    .B(_11749_),
    .Y(_11750_));
 sky130_fd_sc_hd__nand3_1 _21810_ (.A(_11687_),
    .B(_11007_),
    .C(_11018_),
    .Y(_11751_));
 sky130_fd_sc_hd__nand2_1 _21811_ (.A(_11750_),
    .B(_11751_),
    .Y(_11752_));
 sky130_fd_sc_hd__nand2_1 _21812_ (.A(_11752_),
    .B(_07905_),
    .Y(_11753_));
 sky130_fd_sc_hd__buf_6 _21813_ (.A(_06772_),
    .X(_11754_));
 sky130_fd_sc_hd__nand3_1 _21814_ (.A(_11750_),
    .B(_11754_),
    .C(_11751_),
    .Y(_11756_));
 sky130_fd_sc_hd__nand3_1 _21815_ (.A(_11753_),
    .B(_11756_),
    .C(_11694_),
    .Y(_11757_));
 sky130_fd_sc_hd__nor2_1 _21816_ (.A(_11757_),
    .B(_11676_),
    .Y(_11758_));
 sky130_fd_sc_hd__nand2_2 _21817_ (.A(_11654_),
    .B(_11758_),
    .Y(_11759_));
 sky130_fd_sc_hd__nor2_1 _21818_ (.A(_11757_),
    .B(_11681_),
    .Y(_11760_));
 sky130_fd_sc_hd__nand2_1 _21819_ (.A(_11753_),
    .B(_11756_),
    .Y(_11761_));
 sky130_fd_sc_hd__o21ai_1 _21820_ (.A1(_11692_),
    .A2(_11761_),
    .B1(_11756_),
    .Y(_11762_));
 sky130_fd_sc_hd__nor2_2 _21821_ (.A(_11760_),
    .B(_11762_),
    .Y(_11763_));
 sky130_fd_sc_hd__nand2_2 _21822_ (.A(_11759_),
    .B(_11763_),
    .Y(_11764_));
 sky130_fd_sc_hd__clkinvlp_2 _21823_ (.A(_11227_),
    .Y(_11765_));
 sky130_fd_sc_hd__inv_2 _21824_ (.A(_11237_),
    .Y(_11767_));
 sky130_fd_sc_hd__nand2_1 _21825_ (.A(_11191_),
    .B(_11767_),
    .Y(_11768_));
 sky130_fd_sc_hd__nand2_1 _21826_ (.A(_11768_),
    .B(_11236_),
    .Y(_11769_));
 sky130_fd_sc_hd__or2_1 _21827_ (.A(_11765_),
    .B(_11769_),
    .X(_11770_));
 sky130_fd_sc_hd__nand2_1 _21828_ (.A(_11769_),
    .B(_11765_),
    .Y(_11771_));
 sky130_fd_sc_hd__nand2_1 _21829_ (.A(_11770_),
    .B(_11771_),
    .Y(_11772_));
 sky130_fd_sc_hd__nand2_1 _21830_ (.A(_11772_),
    .B(_07957_),
    .Y(_11773_));
 sky130_fd_sc_hd__buf_6 _21831_ (.A(_06827_),
    .X(_11774_));
 sky130_fd_sc_hd__nand3_1 _21832_ (.A(_11770_),
    .B(_11774_),
    .C(_11771_),
    .Y(_11775_));
 sky130_fd_sc_hd__nand2_1 _21833_ (.A(_11773_),
    .B(_11775_),
    .Y(_11776_));
 sky130_fd_sc_hd__or2_1 _21834_ (.A(_11767_),
    .B(_11191_),
    .X(_11778_));
 sky130_fd_sc_hd__nand2_1 _21835_ (.A(_11778_),
    .B(_11768_),
    .Y(_11779_));
 sky130_fd_sc_hd__inv_2 _21836_ (.A(_11779_),
    .Y(_11780_));
 sky130_fd_sc_hd__nand2_1 _21837_ (.A(_11780_),
    .B(_11199_),
    .Y(_11781_));
 sky130_fd_sc_hd__nand2_1 _21838_ (.A(_11779_),
    .B(_08465_),
    .Y(_11782_));
 sky130_fd_sc_hd__nand2_1 _21839_ (.A(_11781_),
    .B(_11782_),
    .Y(_11783_));
 sky130_fd_sc_hd__inv_2 _21840_ (.A(_11783_),
    .Y(_11784_));
 sky130_fd_sc_hd__nand2b_1 _21841_ (.A_N(_11776_),
    .B(_11784_),
    .Y(_11785_));
 sky130_fd_sc_hd__inv_2 _21842_ (.A(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__nand2_1 _21843_ (.A(_11764_),
    .B(_11786_),
    .Y(_11787_));
 sky130_fd_sc_hd__inv_2 _21844_ (.A(_11781_),
    .Y(_11789_));
 sky130_fd_sc_hd__a21boi_2 _21845_ (.A1(_11773_),
    .A2(_11789_),
    .B1_N(_11775_),
    .Y(_11790_));
 sky130_fd_sc_hd__nand2_1 _21846_ (.A(_11787_),
    .B(_11790_),
    .Y(_11791_));
 sky130_fd_sc_hd__inv_2 _21847_ (.A(_11281_),
    .Y(_11792_));
 sky130_fd_sc_hd__nand2_1 _21848_ (.A(_11243_),
    .B(_11792_),
    .Y(_11793_));
 sky130_fd_sc_hd__nand3_1 _21849_ (.A(_11240_),
    .B(_11242_),
    .C(_11281_),
    .Y(_11794_));
 sky130_fd_sc_hd__nand2_1 _21850_ (.A(_11793_),
    .B(_11794_),
    .Y(_11795_));
 sky130_fd_sc_hd__inv_2 _21851_ (.A(_11795_),
    .Y(_11796_));
 sky130_fd_sc_hd__buf_6 _21852_ (.A(_06819_),
    .X(_11797_));
 sky130_fd_sc_hd__nand2_1 _21853_ (.A(_11796_),
    .B(_11797_),
    .Y(_11798_));
 sky130_fd_sc_hd__nand2_1 _21854_ (.A(_11795_),
    .B(_07948_),
    .Y(_11800_));
 sky130_fd_sc_hd__nand2_1 _21855_ (.A(_11798_),
    .B(_11800_),
    .Y(_11801_));
 sky130_fd_sc_hd__inv_2 _21856_ (.A(_11801_),
    .Y(_11802_));
 sky130_fd_sc_hd__nand2_1 _21857_ (.A(_11791_),
    .B(_11802_),
    .Y(_11803_));
 sky130_fd_sc_hd__nand3_1 _21858_ (.A(_11787_),
    .B(_11801_),
    .C(_11790_),
    .Y(_11804_));
 sky130_fd_sc_hd__nand3_1 _21859_ (.A(_11803_),
    .B(_11731_),
    .C(_11804_),
    .Y(_11805_));
 sky130_fd_sc_hd__nand2_1 _21860_ (.A(\div1i.quot[9] ),
    .B(_11796_),
    .Y(_11806_));
 sky130_fd_sc_hd__nand2_1 _21861_ (.A(_11805_),
    .B(_11806_),
    .Y(_11807_));
 sky130_fd_sc_hd__buf_6 _21862_ (.A(_06856_),
    .X(_11808_));
 sky130_fd_sc_hd__nand2_1 _21863_ (.A(_11807_),
    .B(_11808_),
    .Y(_11809_));
 sky130_fd_sc_hd__buf_8 _21864_ (.A(_06809_),
    .X(_11811_));
 sky130_fd_sc_hd__nand3_1 _21865_ (.A(_11805_),
    .B(_11811_),
    .C(_11806_),
    .Y(_11812_));
 sky130_fd_sc_hd__nand2_1 _21866_ (.A(_11809_),
    .B(_11812_),
    .Y(_11813_));
 sky130_fd_sc_hd__nand2_1 _21867_ (.A(_11764_),
    .B(_11784_),
    .Y(_11814_));
 sky130_fd_sc_hd__nand2_1 _21868_ (.A(_11814_),
    .B(_11781_),
    .Y(_11815_));
 sky130_fd_sc_hd__xor2_1 _21869_ (.A(_11776_),
    .B(_11815_),
    .X(_11816_));
 sky130_fd_sc_hd__nand2_1 _21870_ (.A(_11816_),
    .B(_11731_),
    .Y(_11817_));
 sky130_fd_sc_hd__nand2_1 _21871_ (.A(\div1i.quot[9] ),
    .B(_11772_),
    .Y(_11818_));
 sky130_fd_sc_hd__nand2_1 _21872_ (.A(_11817_),
    .B(_11818_),
    .Y(_11819_));
 sky130_fd_sc_hd__nand2_1 _21873_ (.A(_11819_),
    .B(_10173_),
    .Y(_11820_));
 sky130_fd_sc_hd__nand3_2 _21874_ (.A(_11817_),
    .B(_07400_),
    .C(_11818_),
    .Y(_11822_));
 sky130_fd_sc_hd__nand2_1 _21875_ (.A(_11820_),
    .B(_11822_),
    .Y(_11823_));
 sky130_fd_sc_hd__nor2_1 _21876_ (.A(_11813_),
    .B(_11823_),
    .Y(_11824_));
 sky130_fd_sc_hd__nand3_1 _21877_ (.A(_11759_),
    .B(_11783_),
    .C(_11763_),
    .Y(_11825_));
 sky130_fd_sc_hd__nand3_1 _21878_ (.A(_11814_),
    .B(_11581_),
    .C(_11825_),
    .Y(_11826_));
 sky130_fd_sc_hd__nand2_1 _21879_ (.A(net227),
    .B(_11780_),
    .Y(_11827_));
 sky130_fd_sc_hd__nand2_1 _21880_ (.A(_11826_),
    .B(_11827_),
    .Y(_11828_));
 sky130_fd_sc_hd__or2_1 _21881_ (.A(_10138_),
    .B(_11828_),
    .X(_11829_));
 sky130_fd_sc_hd__nand2_1 _21882_ (.A(_11828_),
    .B(_10138_),
    .Y(_11830_));
 sky130_fd_sc_hd__nand2_2 _21883_ (.A(_11829_),
    .B(_11830_),
    .Y(_11831_));
 sky130_fd_sc_hd__nand2_1 _21884_ (.A(_11695_),
    .B(_11692_),
    .Y(_11833_));
 sky130_fd_sc_hd__xor2_1 _21885_ (.A(_11761_),
    .B(_11833_),
    .X(_11834_));
 sky130_fd_sc_hd__nand2_1 _21886_ (.A(_11834_),
    .B(_11731_),
    .Y(_11835_));
 sky130_fd_sc_hd__nand2_1 _21887_ (.A(\div1i.quot[9] ),
    .B(_11752_),
    .Y(_11836_));
 sky130_fd_sc_hd__nand2_1 _21888_ (.A(_11835_),
    .B(_11836_),
    .Y(_11837_));
 sky130_fd_sc_hd__buf_6 _21889_ (.A(_06797_),
    .X(_11838_));
 sky130_fd_sc_hd__nand2_1 _21890_ (.A(_11837_),
    .B(_11838_),
    .Y(_11839_));
 sky130_fd_sc_hd__buf_6 _21891_ (.A(_06799_),
    .X(_11840_));
 sky130_fd_sc_hd__nand3_2 _21892_ (.A(_11835_),
    .B(_11840_),
    .C(_11836_),
    .Y(_11841_));
 sky130_fd_sc_hd__nand3b_2 _21893_ (.A_N(_11831_),
    .B(_11839_),
    .C(_11841_),
    .Y(_11842_));
 sky130_fd_sc_hd__inv_4 _21894_ (.A(_11842_),
    .Y(_11844_));
 sky130_fd_sc_hd__nand3_4 _21895_ (.A(_11747_),
    .B(_11824_),
    .C(_11844_),
    .Y(_11845_));
 sky130_fd_sc_hd__inv_2 _21896_ (.A(_11830_),
    .Y(_11846_));
 sky130_fd_sc_hd__o21bai_2 _21897_ (.A1(_11831_),
    .A2(_11841_),
    .B1_N(_11846_),
    .Y(_11847_));
 sky130_fd_sc_hd__o21ai_1 _21898_ (.A1(_11813_),
    .A2(_11822_),
    .B1(_11809_),
    .Y(_11848_));
 sky130_fd_sc_hd__a21oi_1 _21899_ (.A1(_11824_),
    .A2(_11847_),
    .B1(_11848_),
    .Y(_11849_));
 sky130_fd_sc_hd__nand2_2 _21900_ (.A(_11845_),
    .B(_11849_),
    .Y(_11850_));
 sky130_fd_sc_hd__nand2_1 _21901_ (.A(_11793_),
    .B(_11279_),
    .Y(_11851_));
 sky130_fd_sc_hd__inv_2 _21902_ (.A(_11273_),
    .Y(_11852_));
 sky130_fd_sc_hd__nand2_1 _21903_ (.A(_11851_),
    .B(_11852_),
    .Y(_11853_));
 sky130_fd_sc_hd__nand3_1 _21904_ (.A(_11793_),
    .B(_11273_),
    .C(_11279_),
    .Y(_11855_));
 sky130_fd_sc_hd__nand2_1 _21905_ (.A(_11853_),
    .B(_11855_),
    .Y(_11856_));
 sky130_fd_sc_hd__nand2_1 _21906_ (.A(_11856_),
    .B(_08001_),
    .Y(_11857_));
 sky130_fd_sc_hd__buf_6 _21907_ (.A(_06874_),
    .X(_11858_));
 sky130_fd_sc_hd__nand3_1 _21908_ (.A(_11853_),
    .B(_11858_),
    .C(_11855_),
    .Y(_11859_));
 sky130_fd_sc_hd__nand3_1 _21909_ (.A(_11802_),
    .B(_11857_),
    .C(_11859_),
    .Y(_11860_));
 sky130_fd_sc_hd__inv_2 _21910_ (.A(_11860_),
    .Y(_11861_));
 sky130_fd_sc_hd__nand3_2 _21911_ (.A(_11764_),
    .B(_11786_),
    .C(_11861_),
    .Y(_11862_));
 sky130_fd_sc_hd__inv_2 _21912_ (.A(_11857_),
    .Y(_11863_));
 sky130_fd_sc_hd__o21ai_1 _21913_ (.A1(_11798_),
    .A2(_11863_),
    .B1(_11859_),
    .Y(_11864_));
 sky130_fd_sc_hd__nor2_1 _21914_ (.A(_11790_),
    .B(_11860_),
    .Y(_11866_));
 sky130_fd_sc_hd__nor2_1 _21915_ (.A(_11864_),
    .B(_11866_),
    .Y(_11867_));
 sky130_fd_sc_hd__nand2_1 _21916_ (.A(_11862_),
    .B(_11867_),
    .Y(_11868_));
 sky130_fd_sc_hd__inv_2 _21917_ (.A(_11287_),
    .Y(_11869_));
 sky130_fd_sc_hd__nand2_1 _21918_ (.A(_11331_),
    .B(_11332_),
    .Y(_11870_));
 sky130_fd_sc_hd__nand2_1 _21919_ (.A(_11869_),
    .B(_11870_),
    .Y(_11871_));
 sky130_fd_sc_hd__inv_2 _21920_ (.A(_11870_),
    .Y(_11872_));
 sky130_fd_sc_hd__nand2_1 _21921_ (.A(_11287_),
    .B(_11872_),
    .Y(_11873_));
 sky130_fd_sc_hd__nand2_1 _21922_ (.A(_11871_),
    .B(_11873_),
    .Y(_11874_));
 sky130_fd_sc_hd__nand2_1 _21923_ (.A(_11874_),
    .B(_10749_),
    .Y(_11875_));
 sky130_fd_sc_hd__nand3_2 _21924_ (.A(_11871_),
    .B(_08554_),
    .C(_11873_),
    .Y(_11877_));
 sky130_fd_sc_hd__nand2_1 _21925_ (.A(_11875_),
    .B(_11877_),
    .Y(_11878_));
 sky130_fd_sc_hd__inv_2 _21926_ (.A(_11878_),
    .Y(_11879_));
 sky130_fd_sc_hd__nand2_1 _21927_ (.A(_11868_),
    .B(_11879_),
    .Y(_11880_));
 sky130_fd_sc_hd__nand3_1 _21928_ (.A(_11862_),
    .B(_11867_),
    .C(_11878_),
    .Y(_11881_));
 sky130_fd_sc_hd__nand3_1 _21929_ (.A(_11880_),
    .B(_11731_),
    .C(_11881_),
    .Y(_11882_));
 sky130_fd_sc_hd__or2_1 _21930_ (.A(_11874_),
    .B(_11581_),
    .X(_11883_));
 sky130_fd_sc_hd__nand2_1 _21931_ (.A(_11882_),
    .B(_11883_),
    .Y(_11884_));
 sky130_fd_sc_hd__or2_1 _21932_ (.A(_09664_),
    .B(_11884_),
    .X(_11885_));
 sky130_fd_sc_hd__nand2_1 _21933_ (.A(_11884_),
    .B(_09664_),
    .Y(_11886_));
 sky130_fd_sc_hd__nand2_1 _21934_ (.A(_11885_),
    .B(_11886_),
    .Y(_11888_));
 sky130_fd_sc_hd__inv_2 _21935_ (.A(_11888_),
    .Y(_11889_));
 sky130_fd_sc_hd__nand2_1 _21936_ (.A(_11857_),
    .B(_11859_),
    .Y(_11890_));
 sky130_fd_sc_hd__nand2_1 _21937_ (.A(_11803_),
    .B(_11798_),
    .Y(_11891_));
 sky130_fd_sc_hd__xor2_1 _21938_ (.A(_11890_),
    .B(_11891_),
    .X(_11892_));
 sky130_fd_sc_hd__nand2_1 _21939_ (.A(_11892_),
    .B(_11731_),
    .Y(_11893_));
 sky130_fd_sc_hd__nand2_1 _21940_ (.A(\div1i.quot[9] ),
    .B(_11856_),
    .Y(_11894_));
 sky130_fd_sc_hd__nand2_1 _21941_ (.A(_11893_),
    .B(_11894_),
    .Y(_11895_));
 sky130_fd_sc_hd__buf_6 _21942_ (.A(_06903_),
    .X(_11896_));
 sky130_fd_sc_hd__nand2_1 _21943_ (.A(_11895_),
    .B(_11896_),
    .Y(_11897_));
 sky130_fd_sc_hd__clkbuf_8 _21944_ (.A(_06898_),
    .X(_11899_));
 sky130_fd_sc_hd__nand3_2 _21945_ (.A(_11893_),
    .B(_11899_),
    .C(_11894_),
    .Y(_11900_));
 sky130_fd_sc_hd__nand3_1 _21946_ (.A(_11889_),
    .B(_11897_),
    .C(_11900_),
    .Y(_11901_));
 sky130_fd_sc_hd__nand2_1 _21947_ (.A(_11880_),
    .B(_11877_),
    .Y(_11902_));
 sky130_fd_sc_hd__nand2_1 _21948_ (.A(_11873_),
    .B(_11332_),
    .Y(_11903_));
 sky130_fd_sc_hd__xor2_2 _21949_ (.A(_11322_),
    .B(_11903_),
    .X(_11904_));
 sky130_fd_sc_hd__inv_2 _21950_ (.A(_11904_),
    .Y(_11905_));
 sky130_fd_sc_hd__nand2_1 _21951_ (.A(_11905_),
    .B(_07461_),
    .Y(_11906_));
 sky130_fd_sc_hd__nand2_1 _21952_ (.A(_11904_),
    .B(_08041_),
    .Y(_11907_));
 sky130_fd_sc_hd__nand2_1 _21953_ (.A(_11906_),
    .B(_11907_),
    .Y(_11908_));
 sky130_fd_sc_hd__inv_2 _21954_ (.A(_11908_),
    .Y(_11910_));
 sky130_fd_sc_hd__nand2_1 _21955_ (.A(_11902_),
    .B(_11910_),
    .Y(_11911_));
 sky130_fd_sc_hd__nand3_1 _21956_ (.A(_11880_),
    .B(_11908_),
    .C(_11877_),
    .Y(_11912_));
 sky130_fd_sc_hd__nand2_1 _21957_ (.A(_11911_),
    .B(_11912_),
    .Y(_11913_));
 sky130_fd_sc_hd__nand2_1 _21958_ (.A(_11913_),
    .B(_11731_),
    .Y(_11914_));
 sky130_fd_sc_hd__nand2_1 _21959_ (.A(_11904_),
    .B(\div1i.quot[9] ),
    .Y(_11915_));
 sky130_fd_sc_hd__nand2_1 _21960_ (.A(_11914_),
    .B(_11915_),
    .Y(_11916_));
 sky130_fd_sc_hd__nand2_1 _21961_ (.A(_11916_),
    .B(_07474_),
    .Y(_11917_));
 sky130_fd_sc_hd__nand3_2 _21962_ (.A(_11914_),
    .B(_11376_),
    .C(_11915_),
    .Y(_11918_));
 sky130_fd_sc_hd__nand2_1 _21963_ (.A(_11917_),
    .B(_11918_),
    .Y(_11919_));
 sky130_fd_sc_hd__inv_2 _21964_ (.A(_11919_),
    .Y(_11921_));
 sky130_fd_sc_hd__nand3_1 _21965_ (.A(_11906_),
    .B(_11907_),
    .C(_11879_),
    .Y(_11922_));
 sky130_fd_sc_hd__inv_2 _21966_ (.A(_11922_),
    .Y(_11923_));
 sky130_fd_sc_hd__nand2_1 _21967_ (.A(_11923_),
    .B(_11868_),
    .Y(_11924_));
 sky130_fd_sc_hd__inv_2 _21968_ (.A(_11907_),
    .Y(_11925_));
 sky130_fd_sc_hd__o21a_1 _21969_ (.A1(_11877_),
    .A2(_11925_),
    .B1(_11906_),
    .X(_11926_));
 sky130_fd_sc_hd__nand2_1 _21970_ (.A(_11924_),
    .B(_11926_),
    .Y(_11927_));
 sky130_fd_sc_hd__inv_2 _21971_ (.A(_11378_),
    .Y(_11928_));
 sky130_fd_sc_hd__o21bai_1 _21972_ (.A1(_11333_),
    .A2(_11869_),
    .B1_N(_11384_),
    .Y(_11929_));
 sky130_fd_sc_hd__or2_1 _21973_ (.A(_11928_),
    .B(_11929_),
    .X(_11930_));
 sky130_fd_sc_hd__nand2_1 _21974_ (.A(_11929_),
    .B(_11928_),
    .Y(_11932_));
 sky130_fd_sc_hd__nand2_1 _21975_ (.A(_11930_),
    .B(_11932_),
    .Y(_11933_));
 sky130_fd_sc_hd__inv_2 _21976_ (.A(_11933_),
    .Y(_11934_));
 sky130_fd_sc_hd__buf_6 _21977_ (.A(_06936_),
    .X(_11935_));
 sky130_fd_sc_hd__nand2_1 _21978_ (.A(_11934_),
    .B(_11935_),
    .Y(_11936_));
 sky130_fd_sc_hd__nand2_1 _21979_ (.A(_11933_),
    .B(_08611_),
    .Y(_11937_));
 sky130_fd_sc_hd__nand2_1 _21980_ (.A(_11936_),
    .B(_11937_),
    .Y(_11938_));
 sky130_fd_sc_hd__inv_2 _21981_ (.A(_11938_),
    .Y(_11939_));
 sky130_fd_sc_hd__nand2_1 _21982_ (.A(_11927_),
    .B(_11939_),
    .Y(_11940_));
 sky130_fd_sc_hd__nand3_1 _21983_ (.A(_11924_),
    .B(_11926_),
    .C(_11938_),
    .Y(_11941_));
 sky130_fd_sc_hd__nand3_2 _21984_ (.A(_11940_),
    .B(_11941_),
    .C(_11731_),
    .Y(_11943_));
 sky130_fd_sc_hd__nand2_1 _21985_ (.A(_11934_),
    .B(\div1i.quot[9] ),
    .Y(_11944_));
 sky130_fd_sc_hd__nand2_1 _21986_ (.A(_11943_),
    .B(_11944_),
    .Y(_11945_));
 sky130_fd_sc_hd__buf_6 _21987_ (.A(_06947_),
    .X(_11946_));
 sky130_fd_sc_hd__nand2_1 _21988_ (.A(_11945_),
    .B(_11946_),
    .Y(_11947_));
 sky130_fd_sc_hd__buf_6 _21989_ (.A(_06949_),
    .X(_11948_));
 sky130_fd_sc_hd__nand3_2 _21990_ (.A(_11943_),
    .B(_11948_),
    .C(_11944_),
    .Y(_11949_));
 sky130_fd_sc_hd__nand2_4 _21991_ (.A(_11949_),
    .B(_11947_),
    .Y(_11950_));
 sky130_fd_sc_hd__inv_2 _21992_ (.A(_11950_),
    .Y(_11951_));
 sky130_fd_sc_hd__nand2_1 _21993_ (.A(_11921_),
    .B(_11951_),
    .Y(_11952_));
 sky130_fd_sc_hd__nor2_1 _21994_ (.A(_11901_),
    .B(_11952_),
    .Y(_11954_));
 sky130_fd_sc_hd__nand2_4 _21995_ (.A(_11850_),
    .B(_11954_),
    .Y(_11955_));
 sky130_fd_sc_hd__o21ai_1 _21996_ (.A1(_11888_),
    .A2(_11900_),
    .B1(_11886_),
    .Y(_11956_));
 sky130_fd_sc_hd__nor2_1 _21997_ (.A(_11950_),
    .B(_11919_),
    .Y(_11957_));
 sky130_fd_sc_hd__inv_2 _21998_ (.A(_11949_),
    .Y(_11958_));
 sky130_fd_sc_hd__o21ai_1 _21999_ (.A1(_11918_),
    .A2(_11958_),
    .B1(_11947_),
    .Y(_11959_));
 sky130_fd_sc_hd__a21oi_2 _22000_ (.A1(_11956_),
    .A2(_11957_),
    .B1(_11959_),
    .Y(_11960_));
 sky130_fd_sc_hd__nand2_2 _22001_ (.A(_11960_),
    .B(_11955_),
    .Y(_11961_));
 sky130_fd_sc_hd__nand2_2 _22002_ (.A(_11932_),
    .B(_11377_),
    .Y(_11962_));
 sky130_fd_sc_hd__xor2_4 _22003_ (.A(_11366_),
    .B(_11962_),
    .X(_11963_));
 sky130_fd_sc_hd__nand3_2 _22004_ (.A(_11940_),
    .B(_11731_),
    .C(_11936_),
    .Y(_11965_));
 sky130_fd_sc_hd__xor2_4 _22005_ (.A(_11963_),
    .B(_11965_),
    .X(_11966_));
 sky130_fd_sc_hd__clkinvlp_2 _22006_ (.A(_11966_),
    .Y(_11967_));
 sky130_fd_sc_hd__nand2_4 _22007_ (.A(_11961_),
    .B(_11967_),
    .Y(_11968_));
 sky130_fd_sc_hd__nand3_4 _22008_ (.A(_11955_),
    .B(_11960_),
    .C(_11966_),
    .Y(_11969_));
 sky130_fd_sc_hd__nand2_8 _22009_ (.A(_11968_),
    .B(_11969_),
    .Y(_11970_));
 sky130_fd_sc_hd__buf_8 _22010_ (.A(_11970_),
    .X(_11971_));
 sky130_fd_sc_hd__buf_6 _22011_ (.A(net242),
    .X(\div1i.quot[8] ));
 sky130_fd_sc_hd__nand2_1 _22012_ (.A(_11533_),
    .B(_11629_),
    .Y(_11972_));
 sky130_fd_sc_hd__inv_2 _22013_ (.A(_11633_),
    .Y(_11973_));
 sky130_fd_sc_hd__nand2_1 _22014_ (.A(_11972_),
    .B(_11973_),
    .Y(_11975_));
 sky130_fd_sc_hd__inv_2 _22015_ (.A(_11605_),
    .Y(_11976_));
 sky130_fd_sc_hd__nand2_1 _22016_ (.A(_11975_),
    .B(_11976_),
    .Y(_11977_));
 sky130_fd_sc_hd__nand2_1 _22017_ (.A(_11977_),
    .B(_11604_),
    .Y(_11978_));
 sky130_fd_sc_hd__inv_2 _22018_ (.A(_11591_),
    .Y(_11979_));
 sky130_fd_sc_hd__nand2_1 _22019_ (.A(_11978_),
    .B(_11979_),
    .Y(_11980_));
 sky130_fd_sc_hd__nand3_1 _22020_ (.A(_11977_),
    .B(_11591_),
    .C(_11604_),
    .Y(_11981_));
 sky130_fd_sc_hd__nand2_1 _22021_ (.A(_11980_),
    .B(_11981_),
    .Y(_11982_));
 sky130_fd_sc_hd__buf_6 _22022_ (.A(_07226_),
    .X(_11983_));
 sky130_fd_sc_hd__nand2_2 _22023_ (.A(_11982_),
    .B(_11983_),
    .Y(_11984_));
 sky130_fd_sc_hd__buf_6 _22024_ (.A(_07128_),
    .X(_11986_));
 sky130_fd_sc_hd__nand3_1 _22025_ (.A(_11972_),
    .B(_11605_),
    .C(_11973_),
    .Y(_11987_));
 sky130_fd_sc_hd__nand3_2 _22026_ (.A(_11977_),
    .B(_11986_),
    .C(_11987_),
    .Y(_11988_));
 sky130_fd_sc_hd__clkinvlp_2 _22027_ (.A(_11988_),
    .Y(_11989_));
 sky130_fd_sc_hd__buf_6 _22028_ (.A(_07228_),
    .X(_11990_));
 sky130_fd_sc_hd__nand3_2 _22029_ (.A(_11980_),
    .B(_11990_),
    .C(_11981_),
    .Y(_11991_));
 sky130_fd_sc_hd__nand3_1 _22030_ (.A(_11984_),
    .B(_11989_),
    .C(_11991_),
    .Y(_11992_));
 sky130_fd_sc_hd__nand2_1 _22031_ (.A(_11992_),
    .B(_11991_),
    .Y(_11993_));
 sky130_fd_sc_hd__inv_2 _22032_ (.A(_11628_),
    .Y(_11994_));
 sky130_fd_sc_hd__nand2_1 _22033_ (.A(_11533_),
    .B(_11994_),
    .Y(_11995_));
 sky130_fd_sc_hd__nand2_1 _22034_ (.A(_11995_),
    .B(_11626_),
    .Y(_11997_));
 sky130_fd_sc_hd__inv_2 _22035_ (.A(_11618_),
    .Y(_11998_));
 sky130_fd_sc_hd__nand2_1 _22036_ (.A(_11997_),
    .B(_11998_),
    .Y(_11999_));
 sky130_fd_sc_hd__nand3_1 _22037_ (.A(_11995_),
    .B(_11618_),
    .C(_11626_),
    .Y(_12000_));
 sky130_fd_sc_hd__nand2_1 _22038_ (.A(_11999_),
    .B(_12000_),
    .Y(_12001_));
 sky130_fd_sc_hd__buf_6 _22039_ (.A(_07146_),
    .X(_12002_));
 sky130_fd_sc_hd__nand2_1 _22040_ (.A(_12001_),
    .B(_12002_),
    .Y(_12003_));
 sky130_fd_sc_hd__or2_1 _22041_ (.A(_11994_),
    .B(_11533_),
    .X(_12004_));
 sky130_fd_sc_hd__nand2_1 _22042_ (.A(_12004_),
    .B(_11995_),
    .Y(_12005_));
 sky130_fd_sc_hd__inv_2 _22043_ (.A(_12005_),
    .Y(_12006_));
 sky130_fd_sc_hd__buf_6 _22044_ (.A(_07157_),
    .X(_12008_));
 sky130_fd_sc_hd__nand2_1 _22045_ (.A(_12006_),
    .B(_12008_),
    .Y(_12009_));
 sky130_fd_sc_hd__inv_2 _22046_ (.A(_12009_),
    .Y(_12010_));
 sky130_fd_sc_hd__inv_2 _22047_ (.A(_12001_),
    .Y(_12011_));
 sky130_fd_sc_hd__buf_6 _22048_ (.A(_07149_),
    .X(_12012_));
 sky130_fd_sc_hd__nand2_1 _22049_ (.A(_12011_),
    .B(_12012_),
    .Y(_12013_));
 sky130_fd_sc_hd__inv_2 _22050_ (.A(_12013_),
    .Y(_12014_));
 sky130_fd_sc_hd__a21oi_2 _22051_ (.A1(_12003_),
    .A2(_12010_),
    .B1(_12014_),
    .Y(_12015_));
 sky130_fd_sc_hd__nand2_1 _22052_ (.A(_11977_),
    .B(_11987_),
    .Y(_12016_));
 sky130_fd_sc_hd__buf_6 _22053_ (.A(_07130_),
    .X(_12017_));
 sky130_fd_sc_hd__nand2_1 _22054_ (.A(_12016_),
    .B(_12017_),
    .Y(_12019_));
 sky130_fd_sc_hd__nand2_1 _22055_ (.A(_12019_),
    .B(_11988_),
    .Y(_12020_));
 sky130_fd_sc_hd__inv_2 _22056_ (.A(_12020_),
    .Y(_12021_));
 sky130_fd_sc_hd__nand3_1 _22057_ (.A(_11984_),
    .B(_12021_),
    .C(_11991_),
    .Y(_12022_));
 sky130_fd_sc_hd__nor2_1 _22058_ (.A(_12015_),
    .B(_12022_),
    .Y(_12023_));
 sky130_fd_sc_hd__nor2_1 _22059_ (.A(_11993_),
    .B(_12023_),
    .Y(_12024_));
 sky130_fd_sc_hd__inv_2 _22060_ (.A(_12022_),
    .Y(_12025_));
 sky130_fd_sc_hd__nand2_1 _22061_ (.A(_11422_),
    .B(_11427_),
    .Y(_12026_));
 sky130_fd_sc_hd__nand2_1 _22062_ (.A(_12026_),
    .B(_11428_),
    .Y(_12027_));
 sky130_fd_sc_hd__nand2_1 _22063_ (.A(_12027_),
    .B(_11430_),
    .Y(_12028_));
 sky130_fd_sc_hd__buf_6 _22064_ (.A(_06982_),
    .X(_12030_));
 sky130_fd_sc_hd__nand2_1 _22065_ (.A(_12028_),
    .B(_12030_),
    .Y(_12031_));
 sky130_fd_sc_hd__buf_6 _22066_ (.A(_09215_),
    .X(_12032_));
 sky130_fd_sc_hd__buf_6 _22067_ (.A(_09228_),
    .X(_12033_));
 sky130_fd_sc_hd__o21ai_1 _22068_ (.A1(_12032_),
    .A2(\div1i.quot[9] ),
    .B1(_12033_),
    .Y(_12034_));
 sky130_fd_sc_hd__buf_6 _22069_ (.A(_06984_),
    .X(_12035_));
 sky130_fd_sc_hd__nand3_1 _22070_ (.A(_12027_),
    .B(_12035_),
    .C(_11430_),
    .Y(_12036_));
 sky130_fd_sc_hd__inv_2 _22071_ (.A(_12036_),
    .Y(_12037_));
 sky130_fd_sc_hd__a21o_1 _22072_ (.A1(_12031_),
    .A2(_12034_),
    .B1(_12037_),
    .X(_12038_));
 sky130_fd_sc_hd__nand2_1 _22073_ (.A(_11431_),
    .B(_11411_),
    .Y(_12039_));
 sky130_fd_sc_hd__nand2_1 _22074_ (.A(_11430_),
    .B(_11422_),
    .Y(_12041_));
 sky130_fd_sc_hd__xor2_1 _22075_ (.A(_12039_),
    .B(_12041_),
    .X(_12042_));
 sky130_fd_sc_hd__buf_6 _22076_ (.A(_07043_),
    .X(_12043_));
 sky130_fd_sc_hd__nand2_1 _22077_ (.A(_12042_),
    .B(_12043_),
    .Y(_12044_));
 sky130_fd_sc_hd__nand2_1 _22078_ (.A(_12038_),
    .B(_12044_),
    .Y(_12045_));
 sky130_fd_sc_hd__inv_2 _22079_ (.A(_12042_),
    .Y(_12046_));
 sky130_fd_sc_hd__buf_6 _22080_ (.A(_07048_),
    .X(_12047_));
 sky130_fd_sc_hd__nand2_1 _22081_ (.A(_12046_),
    .B(_12047_),
    .Y(_12048_));
 sky130_fd_sc_hd__nand2_1 _22082_ (.A(_12045_),
    .B(_12048_),
    .Y(_12049_));
 sky130_fd_sc_hd__nand2_1 _22083_ (.A(_11424_),
    .B(_11430_),
    .Y(_12050_));
 sky130_fd_sc_hd__nand2_1 _22084_ (.A(_12050_),
    .B(_11431_),
    .Y(_12052_));
 sky130_fd_sc_hd__nand2_1 _22085_ (.A(_12052_),
    .B(_11521_),
    .Y(_12053_));
 sky130_fd_sc_hd__nand3_1 _22086_ (.A(_12050_),
    .B(_11431_),
    .C(_11522_),
    .Y(_12054_));
 sky130_fd_sc_hd__nand2_1 _22087_ (.A(_12053_),
    .B(_12054_),
    .Y(_12055_));
 sky130_fd_sc_hd__buf_6 _22088_ (.A(_07031_),
    .X(_12056_));
 sky130_fd_sc_hd__nand2_1 _22089_ (.A(_12055_),
    .B(_12056_),
    .Y(_12057_));
 sky130_fd_sc_hd__buf_6 _22090_ (.A(_07034_),
    .X(_12058_));
 sky130_fd_sc_hd__nand3_1 _22091_ (.A(_12053_),
    .B(_12058_),
    .C(_12054_),
    .Y(_12059_));
 sky130_fd_sc_hd__nand2_1 _22092_ (.A(_12057_),
    .B(_12059_),
    .Y(_12060_));
 sky130_fd_sc_hd__inv_2 _22093_ (.A(_12060_),
    .Y(_12061_));
 sky130_fd_sc_hd__nand2_1 _22094_ (.A(_12049_),
    .B(_12061_),
    .Y(_12063_));
 sky130_fd_sc_hd__nand2_1 _22095_ (.A(_12063_),
    .B(_12059_),
    .Y(_12064_));
 sky130_fd_sc_hd__nand2_1 _22096_ (.A(_12054_),
    .B(_11519_),
    .Y(_12065_));
 sky130_fd_sc_hd__xor2_2 _22097_ (.A(_11511_),
    .B(_12065_),
    .X(_12066_));
 sky130_fd_sc_hd__nand2_1 _22098_ (.A(_12066_),
    .B(_09823_),
    .Y(_12067_));
 sky130_fd_sc_hd__nand2_1 _22099_ (.A(_12064_),
    .B(_12067_),
    .Y(_12068_));
 sky130_fd_sc_hd__or2_1 _22100_ (.A(_09823_),
    .B(_12066_),
    .X(_12069_));
 sky130_fd_sc_hd__nand2_1 _22101_ (.A(_12068_),
    .B(_12069_),
    .Y(_12070_));
 sky130_fd_sc_hd__nor2_1 _22102_ (.A(_11511_),
    .B(_11521_),
    .Y(_12071_));
 sky130_fd_sc_hd__nand3_1 _22103_ (.A(_12050_),
    .B(_12071_),
    .C(_11431_),
    .Y(_12072_));
 sky130_fd_sc_hd__inv_2 _22104_ (.A(_11528_),
    .Y(_12074_));
 sky130_fd_sc_hd__nand2_1 _22105_ (.A(_12072_),
    .B(_12074_),
    .Y(_12075_));
 sky130_fd_sc_hd__nand2_1 _22106_ (.A(_12075_),
    .B(_11499_),
    .Y(_12076_));
 sky130_fd_sc_hd__nand2_1 _22107_ (.A(_12076_),
    .B(_11495_),
    .Y(_12077_));
 sky130_fd_sc_hd__nand2_1 _22108_ (.A(_12077_),
    .B(_11487_),
    .Y(_12078_));
 sky130_fd_sc_hd__nand3_1 _22109_ (.A(_12076_),
    .B(_11486_),
    .C(_11495_),
    .Y(_12079_));
 sky130_fd_sc_hd__nand2_1 _22110_ (.A(_12078_),
    .B(_12079_),
    .Y(_12080_));
 sky130_fd_sc_hd__nand2_1 _22111_ (.A(_12080_),
    .B(_08738_),
    .Y(_12081_));
 sky130_fd_sc_hd__nand3_1 _22112_ (.A(_12072_),
    .B(_11498_),
    .C(_12074_),
    .Y(_12082_));
 sky130_fd_sc_hd__nand2_1 _22113_ (.A(_12076_),
    .B(_12082_),
    .Y(_12083_));
 sky130_fd_sc_hd__buf_6 _22114_ (.A(_07024_),
    .X(_12085_));
 sky130_fd_sc_hd__nand2_1 _22115_ (.A(_12083_),
    .B(_12085_),
    .Y(_12086_));
 sky130_fd_sc_hd__buf_6 _22116_ (.A(_07021_),
    .X(_12087_));
 sky130_fd_sc_hd__nand3_2 _22117_ (.A(_12076_),
    .B(_12087_),
    .C(_12082_),
    .Y(_12088_));
 sky130_fd_sc_hd__nand2_1 _22118_ (.A(_12086_),
    .B(_12088_),
    .Y(_12089_));
 sky130_fd_sc_hd__inv_2 _22119_ (.A(_12089_),
    .Y(_12090_));
 sky130_fd_sc_hd__nand3_1 _22120_ (.A(_12078_),
    .B(_10939_),
    .C(_12079_),
    .Y(_12091_));
 sky130_fd_sc_hd__nand3_1 _22121_ (.A(_12081_),
    .B(_12090_),
    .C(_12091_),
    .Y(_12092_));
 sky130_fd_sc_hd__inv_2 _22122_ (.A(_12092_),
    .Y(_12093_));
 sky130_fd_sc_hd__nand2_1 _22123_ (.A(_12070_),
    .B(_12093_),
    .Y(_12094_));
 sky130_fd_sc_hd__inv_2 _22124_ (.A(_12088_),
    .Y(_12096_));
 sky130_fd_sc_hd__a21boi_1 _22125_ (.A1(_12081_),
    .A2(_12096_),
    .B1_N(_12091_),
    .Y(_12097_));
 sky130_fd_sc_hd__nand2_1 _22126_ (.A(_12094_),
    .B(_12097_),
    .Y(_12098_));
 sky130_fd_sc_hd__nand2_1 _22127_ (.A(_12013_),
    .B(_12003_),
    .Y(_12099_));
 sky130_fd_sc_hd__inv_2 _22128_ (.A(_12099_),
    .Y(_12100_));
 sky130_fd_sc_hd__buf_6 _22129_ (.A(_07155_),
    .X(_12101_));
 sky130_fd_sc_hd__nand2_1 _22130_ (.A(_12005_),
    .B(_12101_),
    .Y(_12102_));
 sky130_fd_sc_hd__nand2_1 _22131_ (.A(_12009_),
    .B(_12102_),
    .Y(_12103_));
 sky130_fd_sc_hd__inv_4 _22132_ (.A(_12103_),
    .Y(_12104_));
 sky130_fd_sc_hd__nand2_1 _22133_ (.A(_12100_),
    .B(_12104_),
    .Y(_12105_));
 sky130_fd_sc_hd__inv_2 _22134_ (.A(_12105_),
    .Y(_12107_));
 sky130_fd_sc_hd__nand3_1 _22135_ (.A(_12025_),
    .B(_12098_),
    .C(_12107_),
    .Y(_12108_));
 sky130_fd_sc_hd__nand2_2 _22136_ (.A(_12024_),
    .B(_12108_),
    .Y(_12109_));
 sky130_fd_sc_hd__inv_2 _22137_ (.A(_11728_),
    .Y(_12110_));
 sky130_fd_sc_hd__inv_2 _22138_ (.A(_11738_),
    .Y(_12111_));
 sky130_fd_sc_hd__nand2_1 _22139_ (.A(_11637_),
    .B(_12111_),
    .Y(_12112_));
 sky130_fd_sc_hd__nand2_1 _22140_ (.A(_12112_),
    .B(_11737_),
    .Y(_12113_));
 sky130_fd_sc_hd__or2_1 _22141_ (.A(_12110_),
    .B(_12113_),
    .X(_12114_));
 sky130_fd_sc_hd__nand2_1 _22142_ (.A(_12113_),
    .B(_12110_),
    .Y(_12115_));
 sky130_fd_sc_hd__nand2_1 _22143_ (.A(_12114_),
    .B(_12115_),
    .Y(_12116_));
 sky130_fd_sc_hd__buf_6 _22144_ (.A(_07247_),
    .X(_12118_));
 sky130_fd_sc_hd__nand2_1 _22145_ (.A(_12116_),
    .B(_12118_),
    .Y(_12119_));
 sky130_fd_sc_hd__buf_6 _22146_ (.A(_07249_),
    .X(_12120_));
 sky130_fd_sc_hd__nand3_1 _22147_ (.A(_12114_),
    .B(_12120_),
    .C(_12115_),
    .Y(_12121_));
 sky130_fd_sc_hd__nand2_1 _22148_ (.A(_12119_),
    .B(_12121_),
    .Y(_12122_));
 sky130_fd_sc_hd__inv_2 _22149_ (.A(_12122_),
    .Y(_12123_));
 sky130_fd_sc_hd__or2_1 _22150_ (.A(_12111_),
    .B(_11637_),
    .X(_12124_));
 sky130_fd_sc_hd__nand2_1 _22151_ (.A(_12124_),
    .B(_12112_),
    .Y(_12125_));
 sky130_fd_sc_hd__inv_2 _22152_ (.A(_12125_),
    .Y(_12126_));
 sky130_fd_sc_hd__nand2_1 _22153_ (.A(_12126_),
    .B(_11671_),
    .Y(_12127_));
 sky130_fd_sc_hd__nand2_1 _22154_ (.A(_12125_),
    .B(_07677_),
    .Y(_12129_));
 sky130_fd_sc_hd__nand2_1 _22155_ (.A(_12127_),
    .B(_12129_),
    .Y(_12130_));
 sky130_fd_sc_hd__inv_2 _22156_ (.A(_12130_),
    .Y(_12131_));
 sky130_fd_sc_hd__nand2_1 _22157_ (.A(_12123_),
    .B(_12131_),
    .Y(_12132_));
 sky130_fd_sc_hd__inv_2 _22158_ (.A(_12132_),
    .Y(_12133_));
 sky130_fd_sc_hd__nand2_1 _22159_ (.A(_12109_),
    .B(_12133_),
    .Y(_12134_));
 sky130_fd_sc_hd__inv_2 _22160_ (.A(_12127_),
    .Y(_12135_));
 sky130_fd_sc_hd__a21boi_2 _22161_ (.A1(_12119_),
    .A2(_12135_),
    .B1_N(_12121_),
    .Y(_12136_));
 sky130_fd_sc_hd__nand2_1 _22162_ (.A(_12134_),
    .B(_12136_),
    .Y(_12137_));
 sky130_fd_sc_hd__nand2_1 _22163_ (.A(_11637_),
    .B(_11739_),
    .Y(_12138_));
 sky130_fd_sc_hd__inv_2 _22164_ (.A(_11743_),
    .Y(_12140_));
 sky130_fd_sc_hd__nand2_1 _22165_ (.A(_12138_),
    .B(_12140_),
    .Y(_12141_));
 sky130_fd_sc_hd__inv_2 _22166_ (.A(_11719_),
    .Y(_12142_));
 sky130_fd_sc_hd__nand2_1 _22167_ (.A(_12141_),
    .B(_12142_),
    .Y(_12143_));
 sky130_fd_sc_hd__nand3_1 _22168_ (.A(_12138_),
    .B(_11719_),
    .C(_12140_),
    .Y(_12144_));
 sky130_fd_sc_hd__nand2_1 _22169_ (.A(_12143_),
    .B(_12144_),
    .Y(_12145_));
 sky130_fd_sc_hd__inv_2 _22170_ (.A(_12145_),
    .Y(_12146_));
 sky130_fd_sc_hd__buf_6 _22171_ (.A(_07278_),
    .X(_12147_));
 sky130_fd_sc_hd__nand2_1 _22172_ (.A(_12146_),
    .B(_12147_),
    .Y(_12148_));
 sky130_fd_sc_hd__buf_6 _22173_ (.A(_07276_),
    .X(_12149_));
 sky130_fd_sc_hd__nand2_1 _22174_ (.A(_12145_),
    .B(_12149_),
    .Y(_12151_));
 sky130_fd_sc_hd__nand2_1 _22175_ (.A(_12148_),
    .B(_12151_),
    .Y(_12152_));
 sky130_fd_sc_hd__inv_2 _22176_ (.A(_12152_),
    .Y(_12153_));
 sky130_fd_sc_hd__nand2_1 _22177_ (.A(_12137_),
    .B(_12153_),
    .Y(_12154_));
 sky130_fd_sc_hd__inv_6 _22178_ (.A(_11970_),
    .Y(_12155_));
 sky130_fd_sc_hd__nand3_1 _22179_ (.A(_12134_),
    .B(_12152_),
    .C(_12136_),
    .Y(_12156_));
 sky130_fd_sc_hd__nand3_1 _22180_ (.A(_12154_),
    .B(_12155_),
    .C(_12156_),
    .Y(_12157_));
 sky130_fd_sc_hd__nand2_1 _22181_ (.A(net242),
    .B(_12146_),
    .Y(_12158_));
 sky130_fd_sc_hd__nand2_1 _22182_ (.A(_12157_),
    .B(_12158_),
    .Y(_12159_));
 sky130_fd_sc_hd__nand2_1 _22183_ (.A(_12159_),
    .B(_11701_),
    .Y(_12160_));
 sky130_fd_sc_hd__nand3_1 _22184_ (.A(_12157_),
    .B(_11703_),
    .C(_12158_),
    .Y(_12162_));
 sky130_fd_sc_hd__nand2_1 _22185_ (.A(_12160_),
    .B(_12162_),
    .Y(_12163_));
 sky130_fd_sc_hd__nand2_1 _22186_ (.A(_12109_),
    .B(_12131_),
    .Y(_12164_));
 sky130_fd_sc_hd__nand2_1 _22187_ (.A(_12164_),
    .B(_12127_),
    .Y(_12165_));
 sky130_fd_sc_hd__nand2_1 _22188_ (.A(_12165_),
    .B(_12123_),
    .Y(_12166_));
 sky130_fd_sc_hd__nand3_1 _22189_ (.A(_12164_),
    .B(_12122_),
    .C(_12127_),
    .Y(_12167_));
 sky130_fd_sc_hd__nand2_1 _22190_ (.A(_12166_),
    .B(_12167_),
    .Y(_12168_));
 sky130_fd_sc_hd__nand2_1 _22191_ (.A(_12168_),
    .B(_12155_),
    .Y(_12169_));
 sky130_fd_sc_hd__nand2_1 _22192_ (.A(net242),
    .B(_12116_),
    .Y(_12170_));
 sky130_fd_sc_hd__nand2_1 _22193_ (.A(_12169_),
    .B(_12170_),
    .Y(_12171_));
 sky130_fd_sc_hd__nand2_1 _22194_ (.A(_12171_),
    .B(_11715_),
    .Y(_12173_));
 sky130_fd_sc_hd__nand3_2 _22195_ (.A(_12169_),
    .B(_11717_),
    .C(_12170_),
    .Y(_12174_));
 sky130_fd_sc_hd__nand2_1 _22196_ (.A(_12173_),
    .B(_12174_),
    .Y(_12175_));
 sky130_fd_sc_hd__nor2_1 _22197_ (.A(_12163_),
    .B(_12175_),
    .Y(_12176_));
 sky130_fd_sc_hd__nand2_1 _22198_ (.A(_12107_),
    .B(_12098_),
    .Y(_12177_));
 sky130_fd_sc_hd__nand2_1 _22199_ (.A(_12177_),
    .B(_12015_),
    .Y(_12178_));
 sky130_fd_sc_hd__nand2_1 _22200_ (.A(_12178_),
    .B(_12021_),
    .Y(_12179_));
 sky130_fd_sc_hd__nand2_1 _22201_ (.A(_12179_),
    .B(_11988_),
    .Y(_12180_));
 sky130_fd_sc_hd__nand3_1 _22202_ (.A(_12180_),
    .B(_11991_),
    .C(_11984_),
    .Y(_12181_));
 sky130_fd_sc_hd__nand2_1 _22203_ (.A(_11984_),
    .B(_11991_),
    .Y(_12182_));
 sky130_fd_sc_hd__nand3_1 _22204_ (.A(_12179_),
    .B(_11988_),
    .C(_12182_),
    .Y(_12184_));
 sky130_fd_sc_hd__nand2_1 _22205_ (.A(_12181_),
    .B(_12184_),
    .Y(_12185_));
 sky130_fd_sc_hd__nand2_1 _22206_ (.A(_12185_),
    .B(_12155_),
    .Y(_12186_));
 sky130_fd_sc_hd__buf_6 _22207_ (.A(_07318_),
    .X(_12187_));
 sky130_fd_sc_hd__nand2_1 _22208_ (.A(net242),
    .B(_11982_),
    .Y(_12188_));
 sky130_fd_sc_hd__nand3_2 _22209_ (.A(_12186_),
    .B(_12187_),
    .C(_12188_),
    .Y(_12189_));
 sky130_fd_sc_hd__or2_1 _22210_ (.A(_12131_),
    .B(_12109_),
    .X(_12190_));
 sky130_fd_sc_hd__nand3_1 _22211_ (.A(_12190_),
    .B(_12155_),
    .C(_12164_),
    .Y(_12191_));
 sky130_fd_sc_hd__nand2_1 _22212_ (.A(net242),
    .B(_12126_),
    .Y(_12192_));
 sky130_fd_sc_hd__nand3_1 _22213_ (.A(_12191_),
    .B(_09944_),
    .C(_12192_),
    .Y(_12193_));
 sky130_fd_sc_hd__inv_2 _22214_ (.A(_12193_),
    .Y(_12195_));
 sky130_fd_sc_hd__a21o_1 _22215_ (.A1(_12191_),
    .A2(_12192_),
    .B1(_09944_),
    .X(_12196_));
 sky130_fd_sc_hd__o21ai_2 _22216_ (.A1(_12189_),
    .A2(_12195_),
    .B1(_12196_),
    .Y(_12197_));
 sky130_fd_sc_hd__inv_2 _22217_ (.A(_12162_),
    .Y(_12198_));
 sky130_fd_sc_hd__o21ai_1 _22218_ (.A1(_12174_),
    .A2(_12198_),
    .B1(_12160_),
    .Y(_12199_));
 sky130_fd_sc_hd__a21oi_1 _22219_ (.A1(_12176_),
    .A2(_12197_),
    .B1(_12199_),
    .Y(_12200_));
 sky130_fd_sc_hd__inv_2 _22220_ (.A(_12028_),
    .Y(_12201_));
 sky130_fd_sc_hd__nand2_1 _22221_ (.A(_11971_),
    .B(_12201_),
    .Y(_12202_));
 sky130_fd_sc_hd__nand2_1 _22222_ (.A(_12031_),
    .B(_12036_),
    .Y(_12203_));
 sky130_fd_sc_hd__xor2_1 _22223_ (.A(_12034_),
    .B(_12203_),
    .X(_12204_));
 sky130_fd_sc_hd__nand3b_1 _22224_ (.A_N(_12204_),
    .B(_11968_),
    .C(_11969_),
    .Y(_12206_));
 sky130_fd_sc_hd__nand2_1 _22225_ (.A(_12202_),
    .B(_12206_),
    .Y(_12207_));
 sky130_fd_sc_hd__nand2_1 _22226_ (.A(_12207_),
    .B(_11069_),
    .Y(_12208_));
 sky130_fd_sc_hd__nor2_1 _22227_ (.A(_12032_),
    .B(_11731_),
    .Y(_12209_));
 sky130_fd_sc_hd__or2_1 _22228_ (.A(_11412_),
    .B(_12209_),
    .X(_12210_));
 sky130_fd_sc_hd__nand2_1 _22229_ (.A(_12210_),
    .B(_11428_),
    .Y(_12211_));
 sky130_fd_sc_hd__inv_2 _22230_ (.A(_12211_),
    .Y(_12212_));
 sky130_fd_sc_hd__nand2_1 _22231_ (.A(_11970_),
    .B(_12212_),
    .Y(_12213_));
 sky130_fd_sc_hd__nand3_1 _22232_ (.A(_11968_),
    .B(_11969_),
    .C(_12209_),
    .Y(_12214_));
 sky130_fd_sc_hd__nand2_1 _22233_ (.A(_12213_),
    .B(_12214_),
    .Y(_12215_));
 sky130_fd_sc_hd__nand2_2 _22234_ (.A(_12215_),
    .B(_11421_),
    .Y(_12217_));
 sky130_fd_sc_hd__nand2_1 _22235_ (.A(_12208_),
    .B(_12217_),
    .Y(_12218_));
 sky130_fd_sc_hd__inv_2 _22236_ (.A(_12218_),
    .Y(_12219_));
 sky130_fd_sc_hd__nand3_1 _22237_ (.A(_12213_),
    .B(_11426_),
    .C(_12214_),
    .Y(_12220_));
 sky130_fd_sc_hd__buf_6 _22238_ (.A(_07004_),
    .X(_12221_));
 sky130_fd_sc_hd__nand3_2 _22239_ (.A(_11971_),
    .B(_12033_),
    .C(_12221_),
    .Y(_12222_));
 sky130_fd_sc_hd__inv_2 _22240_ (.A(_12222_),
    .Y(_12223_));
 sky130_fd_sc_hd__nand3_4 _22241_ (.A(_12217_),
    .B(_12220_),
    .C(_12223_),
    .Y(_12224_));
 sky130_fd_sc_hd__or2_4 _22242_ (.A(_11069_),
    .B(_12207_),
    .X(_12225_));
 sky130_fd_sc_hd__a21boi_2 _22243_ (.A1(_12219_),
    .A2(_12224_),
    .B1_N(_12225_),
    .Y(_12226_));
 sky130_fd_sc_hd__clkinvlp_2 _22244_ (.A(_12083_),
    .Y(_12228_));
 sky130_fd_sc_hd__nand2_1 _22245_ (.A(_11970_),
    .B(_12228_),
    .Y(_12229_));
 sky130_fd_sc_hd__nand2_1 _22246_ (.A(_12070_),
    .B(_12090_),
    .Y(_12230_));
 sky130_fd_sc_hd__nand3_1 _22247_ (.A(_12068_),
    .B(_12089_),
    .C(_12069_),
    .Y(_12231_));
 sky130_fd_sc_hd__nand2_1 _22248_ (.A(_12230_),
    .B(_12231_),
    .Y(_12232_));
 sky130_fd_sc_hd__inv_2 _22249_ (.A(_12232_),
    .Y(_12233_));
 sky130_fd_sc_hd__nand3_1 _22250_ (.A(_11968_),
    .B(_11969_),
    .C(_12233_),
    .Y(_12234_));
 sky130_fd_sc_hd__nand2_1 _22251_ (.A(_12229_),
    .B(_12234_),
    .Y(_12235_));
 sky130_fd_sc_hd__nand2_1 _22252_ (.A(_12235_),
    .B(_11482_),
    .Y(_12236_));
 sky130_fd_sc_hd__nand3_1 _22253_ (.A(_12229_),
    .B(_11484_),
    .C(_12234_),
    .Y(_12237_));
 sky130_fd_sc_hd__nand2_1 _22254_ (.A(_12236_),
    .B(_12237_),
    .Y(_12239_));
 sky130_fd_sc_hd__clkinvlp_2 _22255_ (.A(_12239_),
    .Y(_12240_));
 sky130_fd_sc_hd__nand2_1 _22256_ (.A(_11971_),
    .B(_12066_),
    .Y(_12241_));
 sky130_fd_sc_hd__nand2_1 _22257_ (.A(_12069_),
    .B(_12067_),
    .Y(_12242_));
 sky130_fd_sc_hd__xor2_1 _22258_ (.A(_12064_),
    .B(_12242_),
    .X(_12243_));
 sky130_fd_sc_hd__nand3_1 _22259_ (.A(_11968_),
    .B(_11969_),
    .C(_12243_),
    .Y(_12244_));
 sky130_fd_sc_hd__nand2_1 _22260_ (.A(_12241_),
    .B(_12244_),
    .Y(_12245_));
 sky130_fd_sc_hd__nand2_1 _22261_ (.A(_12245_),
    .B(_11496_),
    .Y(_12246_));
 sky130_fd_sc_hd__nand3_2 _22262_ (.A(_12241_),
    .B(_11494_),
    .C(_12244_),
    .Y(_12247_));
 sky130_fd_sc_hd__nand2_1 _22263_ (.A(_12246_),
    .B(_12247_),
    .Y(_12248_));
 sky130_fd_sc_hd__inv_2 _22264_ (.A(_12248_),
    .Y(_12250_));
 sky130_fd_sc_hd__nand2_1 _22265_ (.A(_12240_),
    .B(_12250_),
    .Y(_12251_));
 sky130_fd_sc_hd__inv_2 _22266_ (.A(_12055_),
    .Y(_12252_));
 sky130_fd_sc_hd__nand2_1 _22267_ (.A(_11970_),
    .B(_12252_),
    .Y(_12253_));
 sky130_fd_sc_hd__or2_1 _22268_ (.A(_12061_),
    .B(_12049_),
    .X(_12254_));
 sky130_fd_sc_hd__nand2_1 _22269_ (.A(_12254_),
    .B(_12063_),
    .Y(_12255_));
 sky130_fd_sc_hd__clkinvlp_2 _22270_ (.A(_12255_),
    .Y(_12256_));
 sky130_fd_sc_hd__nand3_1 _22271_ (.A(_11968_),
    .B(_11969_),
    .C(_12256_),
    .Y(_12257_));
 sky130_fd_sc_hd__nand2_1 _22272_ (.A(_12253_),
    .B(_12257_),
    .Y(_12258_));
 sky130_fd_sc_hd__nand2_1 _22273_ (.A(_12258_),
    .B(_11105_),
    .Y(_12259_));
 sky130_fd_sc_hd__buf_6 _22274_ (.A(_07092_),
    .X(_12261_));
 sky130_fd_sc_hd__nand3_1 _22275_ (.A(_12253_),
    .B(_12261_),
    .C(_12257_),
    .Y(_12262_));
 sky130_fd_sc_hd__nand2_1 _22276_ (.A(_12259_),
    .B(_12262_),
    .Y(_12263_));
 sky130_fd_sc_hd__inv_2 _22277_ (.A(_12263_),
    .Y(_12264_));
 sky130_fd_sc_hd__nand2_1 _22278_ (.A(_11970_),
    .B(_12046_),
    .Y(_12265_));
 sky130_fd_sc_hd__nand2_1 _22279_ (.A(_12048_),
    .B(_12044_),
    .Y(_12266_));
 sky130_fd_sc_hd__xnor2_1 _22280_ (.A(_12038_),
    .B(_12266_),
    .Y(_12267_));
 sky130_fd_sc_hd__nand3_1 _22281_ (.A(_11968_),
    .B(_11969_),
    .C(_12267_),
    .Y(_12268_));
 sky130_fd_sc_hd__nand2_1 _22282_ (.A(_12265_),
    .B(_12268_),
    .Y(_12269_));
 sky130_fd_sc_hd__buf_6 _22283_ (.A(_07102_),
    .X(_12270_));
 sky130_fd_sc_hd__nand2_1 _22284_ (.A(_12269_),
    .B(_12270_),
    .Y(_12272_));
 sky130_fd_sc_hd__nand3_1 _22285_ (.A(_12265_),
    .B(_11117_),
    .C(_12268_),
    .Y(_12273_));
 sky130_fd_sc_hd__nand2_1 _22286_ (.A(_12272_),
    .B(_12273_),
    .Y(_12274_));
 sky130_fd_sc_hd__inv_2 _22287_ (.A(_12274_),
    .Y(_12275_));
 sky130_fd_sc_hd__nand2_1 _22288_ (.A(_12264_),
    .B(_12275_),
    .Y(_12276_));
 sky130_fd_sc_hd__nor2_1 _22289_ (.A(_12251_),
    .B(_12276_),
    .Y(_12277_));
 sky130_fd_sc_hd__nand2_1 _22290_ (.A(_12226_),
    .B(_12277_),
    .Y(_12278_));
 sky130_fd_sc_hd__inv_2 _22291_ (.A(_12262_),
    .Y(_12279_));
 sky130_fd_sc_hd__o21ai_2 _22292_ (.A1(_12272_),
    .A2(_12279_),
    .B1(_12259_),
    .Y(_12280_));
 sky130_fd_sc_hd__nor2_1 _22293_ (.A(_12239_),
    .B(_12248_),
    .Y(_12281_));
 sky130_fd_sc_hd__clkinvlp_2 _22294_ (.A(_12237_),
    .Y(_12283_));
 sky130_fd_sc_hd__o21ai_1 _22295_ (.A1(_12247_),
    .A2(_12283_),
    .B1(_12236_),
    .Y(_12284_));
 sky130_fd_sc_hd__a21oi_1 _22296_ (.A1(_12280_),
    .A2(_12281_),
    .B1(_12284_),
    .Y(_12285_));
 sky130_fd_sc_hd__nand2_2 _22297_ (.A(_12278_),
    .B(_12285_),
    .Y(_12286_));
 sky130_fd_sc_hd__nand2_1 _22298_ (.A(_12098_),
    .B(_12104_),
    .Y(_12287_));
 sky130_fd_sc_hd__or2_1 _22299_ (.A(_12104_),
    .B(_12098_),
    .X(_12288_));
 sky130_fd_sc_hd__nand3_1 _22300_ (.A(_12155_),
    .B(_12287_),
    .C(_12288_),
    .Y(_12289_));
 sky130_fd_sc_hd__nand2_1 _22301_ (.A(_11970_),
    .B(_12006_),
    .Y(_12290_));
 sky130_fd_sc_hd__nand2_1 _22302_ (.A(_12289_),
    .B(_12290_),
    .Y(_12291_));
 sky130_fd_sc_hd__nand2_1 _22303_ (.A(_12291_),
    .B(_11614_),
    .Y(_12292_));
 sky130_fd_sc_hd__nand3_1 _22304_ (.A(_12289_),
    .B(_11616_),
    .C(_12290_),
    .Y(_12294_));
 sky130_fd_sc_hd__nand2_1 _22305_ (.A(_12292_),
    .B(_12294_),
    .Y(_12295_));
 sky130_fd_sc_hd__inv_2 _22306_ (.A(_12295_),
    .Y(_12296_));
 sky130_fd_sc_hd__nand2_1 _22307_ (.A(_12081_),
    .B(_12091_),
    .Y(_12297_));
 sky130_fd_sc_hd__nand2_1 _22308_ (.A(_12230_),
    .B(_12088_),
    .Y(_12298_));
 sky130_fd_sc_hd__xor2_1 _22309_ (.A(_12297_),
    .B(_12298_),
    .X(_12299_));
 sky130_fd_sc_hd__nand2_1 _22310_ (.A(_12299_),
    .B(_12155_),
    .Y(_12300_));
 sky130_fd_sc_hd__nand2_1 _22311_ (.A(_11971_),
    .B(_12080_),
    .Y(_12301_));
 sky130_fd_sc_hd__nand2_1 _22312_ (.A(_12300_),
    .B(_12301_),
    .Y(_12302_));
 sky130_fd_sc_hd__nand2_1 _22313_ (.A(_12302_),
    .B(_09410_),
    .Y(_12303_));
 sky130_fd_sc_hd__nand3_2 _22314_ (.A(_12300_),
    .B(_08951_),
    .C(_12301_),
    .Y(_12305_));
 sky130_fd_sc_hd__nand2_1 _22315_ (.A(_12303_),
    .B(_12305_),
    .Y(_12306_));
 sky130_fd_sc_hd__inv_2 _22316_ (.A(_12306_),
    .Y(_12307_));
 sky130_fd_sc_hd__nand2_1 _22317_ (.A(_12296_),
    .B(_12307_),
    .Y(_12308_));
 sky130_fd_sc_hd__nand2_1 _22318_ (.A(_12287_),
    .B(_12009_),
    .Y(_12309_));
 sky130_fd_sc_hd__nand2_1 _22319_ (.A(_12309_),
    .B(_12100_),
    .Y(_12310_));
 sky130_fd_sc_hd__nand3_1 _22320_ (.A(_12287_),
    .B(_12099_),
    .C(_12009_),
    .Y(_12311_));
 sky130_fd_sc_hd__nand2_1 _22321_ (.A(_12310_),
    .B(_12311_),
    .Y(_12312_));
 sky130_fd_sc_hd__nand2_1 _22322_ (.A(_12312_),
    .B(_12155_),
    .Y(_12313_));
 sky130_fd_sc_hd__nand2_1 _22323_ (.A(_11971_),
    .B(_12001_),
    .Y(_12314_));
 sky130_fd_sc_hd__nand2_1 _22324_ (.A(_12313_),
    .B(_12314_),
    .Y(_12316_));
 sky130_fd_sc_hd__nand2_1 _22325_ (.A(_12316_),
    .B(_11600_),
    .Y(_12317_));
 sky130_fd_sc_hd__nand3_2 _22326_ (.A(_12313_),
    .B(_11603_),
    .C(_12314_),
    .Y(_12318_));
 sky130_fd_sc_hd__nand2_1 _22327_ (.A(_12317_),
    .B(_12318_),
    .Y(_12319_));
 sky130_fd_sc_hd__or2_1 _22328_ (.A(_12016_),
    .B(_12155_),
    .X(_12320_));
 sky130_fd_sc_hd__nand3_1 _22329_ (.A(_12177_),
    .B(_12020_),
    .C(_12015_),
    .Y(_12321_));
 sky130_fd_sc_hd__nand3_1 _22330_ (.A(_12179_),
    .B(_12155_),
    .C(_12321_),
    .Y(_12322_));
 sky130_fd_sc_hd__nand2_1 _22331_ (.A(_12320_),
    .B(_12322_),
    .Y(_12323_));
 sky130_fd_sc_hd__nand2_1 _22332_ (.A(_12323_),
    .B(_11586_),
    .Y(_12324_));
 sky130_fd_sc_hd__nand3_1 _22333_ (.A(_12320_),
    .B(_12322_),
    .C(_11588_),
    .Y(_12325_));
 sky130_fd_sc_hd__nand2_2 _22334_ (.A(_12324_),
    .B(_12325_),
    .Y(_12327_));
 sky130_fd_sc_hd__nor2_1 _22335_ (.A(_12319_),
    .B(_12327_),
    .Y(_12328_));
 sky130_fd_sc_hd__nor2b_1 _22336_ (.A(_12308_),
    .B_N(_12328_),
    .Y(_12329_));
 sky130_fd_sc_hd__nand2_1 _22337_ (.A(_12286_),
    .B(_12329_),
    .Y(_12330_));
 sky130_fd_sc_hd__clkinvlp_2 _22338_ (.A(_12294_),
    .Y(_12331_));
 sky130_fd_sc_hd__o21ai_2 _22339_ (.A1(_12305_),
    .A2(_12331_),
    .B1(_12292_),
    .Y(_12332_));
 sky130_fd_sc_hd__inv_2 _22340_ (.A(_12325_),
    .Y(_12333_));
 sky130_fd_sc_hd__o21ai_1 _22341_ (.A1(_12318_),
    .A2(_12333_),
    .B1(_12324_),
    .Y(_12334_));
 sky130_fd_sc_hd__a21oi_1 _22342_ (.A1(_12328_),
    .A2(_12332_),
    .B1(_12334_),
    .Y(_12335_));
 sky130_fd_sc_hd__nand2_2 _22343_ (.A(_12330_),
    .B(_12335_),
    .Y(_12336_));
 sky130_fd_sc_hd__nand2_1 _22344_ (.A(_12186_),
    .B(_12188_),
    .Y(_12338_));
 sky130_fd_sc_hd__nand2_1 _22345_ (.A(_12338_),
    .B(_11185_),
    .Y(_12339_));
 sky130_fd_sc_hd__nand2_1 _22346_ (.A(_12339_),
    .B(_12189_),
    .Y(_12340_));
 sky130_fd_sc_hd__nand2_1 _22347_ (.A(_12196_),
    .B(_12193_),
    .Y(_12341_));
 sky130_fd_sc_hd__nor2_1 _22348_ (.A(_12340_),
    .B(_12341_),
    .Y(_12342_));
 sky130_fd_sc_hd__nand3_1 _22349_ (.A(_12336_),
    .B(_12176_),
    .C(_12342_),
    .Y(_12343_));
 sky130_fd_sc_hd__nand2_2 _22350_ (.A(_12200_),
    .B(_12343_),
    .Y(_12344_));
 sky130_fd_sc_hd__nand2_1 _22351_ (.A(_11839_),
    .B(_11841_),
    .Y(_12345_));
 sky130_fd_sc_hd__inv_2 _22352_ (.A(_12345_),
    .Y(_12346_));
 sky130_fd_sc_hd__or2_1 _22353_ (.A(_12346_),
    .B(_11747_),
    .X(_12347_));
 sky130_fd_sc_hd__nand2_1 _22354_ (.A(_11747_),
    .B(_12346_),
    .Y(_12349_));
 sky130_fd_sc_hd__nand2_1 _22355_ (.A(_12347_),
    .B(_12349_),
    .Y(_12350_));
 sky130_fd_sc_hd__inv_2 _22356_ (.A(_12350_),
    .Y(_12351_));
 sky130_fd_sc_hd__nand2_1 _22357_ (.A(_12351_),
    .B(_11199_),
    .Y(_12352_));
 sky130_fd_sc_hd__nand2_1 _22358_ (.A(_12350_),
    .B(_08465_),
    .Y(_12353_));
 sky130_fd_sc_hd__nand2_1 _22359_ (.A(_12352_),
    .B(_12353_),
    .Y(_12354_));
 sky130_fd_sc_hd__inv_2 _22360_ (.A(_12354_),
    .Y(_12355_));
 sky130_fd_sc_hd__nand2_1 _22361_ (.A(_12143_),
    .B(_11718_),
    .Y(_12356_));
 sky130_fd_sc_hd__inv_2 _22362_ (.A(_11705_),
    .Y(_12357_));
 sky130_fd_sc_hd__nand2_1 _22363_ (.A(_12356_),
    .B(_12357_),
    .Y(_12358_));
 sky130_fd_sc_hd__nand3_1 _22364_ (.A(_12143_),
    .B(_11705_),
    .C(_11718_),
    .Y(_12360_));
 sky130_fd_sc_hd__nand2_1 _22365_ (.A(_12358_),
    .B(_12360_),
    .Y(_12361_));
 sky130_fd_sc_hd__nand2_1 _22366_ (.A(_12361_),
    .B(_07905_),
    .Y(_12362_));
 sky130_fd_sc_hd__nand3_1 _22367_ (.A(_12358_),
    .B(_11754_),
    .C(_12360_),
    .Y(_12363_));
 sky130_fd_sc_hd__nand3_1 _22368_ (.A(_12153_),
    .B(_12362_),
    .C(_12363_),
    .Y(_12364_));
 sky130_fd_sc_hd__inv_2 _22369_ (.A(_12364_),
    .Y(_12365_));
 sky130_fd_sc_hd__nand3_1 _22370_ (.A(_12109_),
    .B(_12133_),
    .C(_12365_),
    .Y(_12366_));
 sky130_fd_sc_hd__inv_2 _22371_ (.A(_12362_),
    .Y(_12367_));
 sky130_fd_sc_hd__o21ai_1 _22372_ (.A1(_12148_),
    .A2(_12367_),
    .B1(_12363_),
    .Y(_12368_));
 sky130_fd_sc_hd__nor2_1 _22373_ (.A(_12136_),
    .B(_12364_),
    .Y(_12369_));
 sky130_fd_sc_hd__nor2_1 _22374_ (.A(_12368_),
    .B(_12369_),
    .Y(_12371_));
 sky130_fd_sc_hd__nand2_2 _22375_ (.A(_12366_),
    .B(_12371_),
    .Y(_12372_));
 sky130_fd_sc_hd__or2_1 _22376_ (.A(_12355_),
    .B(_12372_),
    .X(_12373_));
 sky130_fd_sc_hd__buf_6 _22377_ (.A(_12155_),
    .X(_12374_));
 sky130_fd_sc_hd__nand2_1 _22378_ (.A(_12372_),
    .B(_12355_),
    .Y(_12375_));
 sky130_fd_sc_hd__nand3_1 _22379_ (.A(_12373_),
    .B(_12374_),
    .C(_12375_),
    .Y(_12376_));
 sky130_fd_sc_hd__nand2_1 _22380_ (.A(\div1i.quot[8] ),
    .B(_12351_),
    .Y(_12377_));
 sky130_fd_sc_hd__nand2_1 _22381_ (.A(_12376_),
    .B(_12377_),
    .Y(_12378_));
 sky130_fd_sc_hd__xor2_2 _22382_ (.A(_06754_),
    .B(_12378_),
    .X(_12379_));
 sky130_fd_sc_hd__nand2_1 _22383_ (.A(_12362_),
    .B(_12363_),
    .Y(_12380_));
 sky130_fd_sc_hd__nand2_1 _22384_ (.A(_12154_),
    .B(_12148_),
    .Y(_12382_));
 sky130_fd_sc_hd__xor2_1 _22385_ (.A(_12380_),
    .B(_12382_),
    .X(_12383_));
 sky130_fd_sc_hd__nand2_1 _22386_ (.A(_12383_),
    .B(_12374_),
    .Y(_12384_));
 sky130_fd_sc_hd__nand2_1 _22387_ (.A(\div1i.quot[8] ),
    .B(_12361_),
    .Y(_12385_));
 sky130_fd_sc_hd__nand2_1 _22388_ (.A(_12384_),
    .B(_12385_),
    .Y(_12386_));
 sky130_fd_sc_hd__nand2_1 _22389_ (.A(_12386_),
    .B(_11838_),
    .Y(_12387_));
 sky130_fd_sc_hd__nand3_1 _22390_ (.A(_12384_),
    .B(_11840_),
    .C(_12385_),
    .Y(_12388_));
 sky130_fd_sc_hd__nand2_1 _22391_ (.A(_12387_),
    .B(_12388_),
    .Y(_12389_));
 sky130_fd_sc_hd__nor2_1 _22392_ (.A(_12379_),
    .B(_12389_),
    .Y(_12390_));
 sky130_fd_sc_hd__nand2_1 _22393_ (.A(_12344_),
    .B(_12390_),
    .Y(_12391_));
 sky130_fd_sc_hd__nand2_1 _22394_ (.A(_12378_),
    .B(_10138_),
    .Y(_12393_));
 sky130_fd_sc_hd__o21a_1 _22395_ (.A1(_12388_),
    .A2(_12379_),
    .B1(_12393_),
    .X(_12394_));
 sky130_fd_sc_hd__nand2_1 _22396_ (.A(_12391_),
    .B(_12394_),
    .Y(_12395_));
 sky130_fd_sc_hd__nand2_1 _22397_ (.A(_11747_),
    .B(_11844_),
    .Y(_12396_));
 sky130_fd_sc_hd__inv_2 _22398_ (.A(_11847_),
    .Y(_12397_));
 sky130_fd_sc_hd__a21o_1 _22399_ (.A1(_12396_),
    .A2(_12397_),
    .B1(_11823_),
    .X(_12398_));
 sky130_fd_sc_hd__nand3_1 _22400_ (.A(_12396_),
    .B(_11823_),
    .C(_12397_),
    .Y(_12399_));
 sky130_fd_sc_hd__nand2_1 _22401_ (.A(_12398_),
    .B(_12399_),
    .Y(_12400_));
 sky130_fd_sc_hd__inv_2 _22402_ (.A(_12400_),
    .Y(_12401_));
 sky130_fd_sc_hd__nand2_1 _22403_ (.A(_12401_),
    .B(_11797_),
    .Y(_12402_));
 sky130_fd_sc_hd__nand2_1 _22404_ (.A(_12400_),
    .B(_07948_),
    .Y(_12404_));
 sky130_fd_sc_hd__nand2_1 _22405_ (.A(_12402_),
    .B(_12404_),
    .Y(_12405_));
 sky130_fd_sc_hd__inv_4 _22406_ (.A(_12405_),
    .Y(_12406_));
 sky130_fd_sc_hd__nand2_1 _22407_ (.A(_12349_),
    .B(_11841_),
    .Y(_12407_));
 sky130_fd_sc_hd__xor2_2 _22408_ (.A(_11831_),
    .B(_12407_),
    .X(_12408_));
 sky130_fd_sc_hd__inv_2 _22409_ (.A(_12408_),
    .Y(_12409_));
 sky130_fd_sc_hd__nand2_1 _22410_ (.A(_12409_),
    .B(_11774_),
    .Y(_12410_));
 sky130_fd_sc_hd__nand2_1 _22411_ (.A(_12408_),
    .B(_07957_),
    .Y(_12411_));
 sky130_fd_sc_hd__nand2_1 _22412_ (.A(_12410_),
    .B(_12411_),
    .Y(_12412_));
 sky130_fd_sc_hd__or2_1 _22413_ (.A(_12354_),
    .B(_12412_),
    .X(_12413_));
 sky130_fd_sc_hd__inv_4 _22414_ (.A(_12413_),
    .Y(_12415_));
 sky130_fd_sc_hd__nand2_1 _22415_ (.A(_12372_),
    .B(_12415_),
    .Y(_12416_));
 sky130_fd_sc_hd__inv_2 _22416_ (.A(_12352_),
    .Y(_12417_));
 sky130_fd_sc_hd__a21boi_1 _22417_ (.A1(_12417_),
    .A2(_12411_),
    .B1_N(_12410_),
    .Y(_12418_));
 sky130_fd_sc_hd__nand2_1 _22418_ (.A(_12416_),
    .B(_12418_),
    .Y(_12419_));
 sky130_fd_sc_hd__or2_1 _22419_ (.A(_12406_),
    .B(_12419_),
    .X(_12420_));
 sky130_fd_sc_hd__nand2_1 _22420_ (.A(_12419_),
    .B(_12406_),
    .Y(_12421_));
 sky130_fd_sc_hd__nand3_1 _22421_ (.A(_12420_),
    .B(_12374_),
    .C(_12421_),
    .Y(_12422_));
 sky130_fd_sc_hd__nand2_1 _22422_ (.A(\div1i.quot[8] ),
    .B(_12401_),
    .Y(_12423_));
 sky130_fd_sc_hd__nand2_1 _22423_ (.A(_12422_),
    .B(_12423_),
    .Y(_12424_));
 sky130_fd_sc_hd__xor2_2 _22424_ (.A(_11811_),
    .B(_12424_),
    .X(_12426_));
 sky130_fd_sc_hd__nand2_1 _22425_ (.A(_12375_),
    .B(_12352_),
    .Y(_12427_));
 sky130_fd_sc_hd__xor2_1 _22426_ (.A(_12412_),
    .B(_12427_),
    .X(_12428_));
 sky130_fd_sc_hd__nand2_1 _22427_ (.A(_12428_),
    .B(_12374_),
    .Y(_12429_));
 sky130_fd_sc_hd__nand2_1 _22428_ (.A(\div1i.quot[8] ),
    .B(_12408_),
    .Y(_12430_));
 sky130_fd_sc_hd__nand2_1 _22429_ (.A(_12429_),
    .B(_12430_),
    .Y(_12431_));
 sky130_fd_sc_hd__or2_1 _22430_ (.A(_10173_),
    .B(_12431_),
    .X(_12432_));
 sky130_fd_sc_hd__nand2_1 _22431_ (.A(_12431_),
    .B(_10173_),
    .Y(_12433_));
 sky130_fd_sc_hd__nand2_1 _22432_ (.A(_12432_),
    .B(_12433_),
    .Y(_12434_));
 sky130_fd_sc_hd__nor2_1 _22433_ (.A(_12426_),
    .B(_12434_),
    .Y(_12435_));
 sky130_fd_sc_hd__nand2_1 _22434_ (.A(_12395_),
    .B(_12435_),
    .Y(_12437_));
 sky130_fd_sc_hd__nand2_1 _22435_ (.A(_12424_),
    .B(_11808_),
    .Y(_12438_));
 sky130_fd_sc_hd__o21a_1 _22436_ (.A1(_12432_),
    .A2(_12426_),
    .B1(_12438_),
    .X(_12439_));
 sky130_fd_sc_hd__nand2_2 _22437_ (.A(_12437_),
    .B(_12439_),
    .Y(_12440_));
 sky130_fd_sc_hd__nand2_1 _22438_ (.A(_11897_),
    .B(_11900_),
    .Y(_12441_));
 sky130_fd_sc_hd__nand2b_1 _22439_ (.A_N(_11850_),
    .B(_12441_),
    .Y(_12442_));
 sky130_fd_sc_hd__nand2b_1 _22440_ (.A_N(_12441_),
    .B(_11850_),
    .Y(_12443_));
 sky130_fd_sc_hd__nand2_1 _22441_ (.A(_12442_),
    .B(_12443_),
    .Y(_12444_));
 sky130_fd_sc_hd__or2_1 _22442_ (.A(_10749_),
    .B(_12444_),
    .X(_12445_));
 sky130_fd_sc_hd__nand2_1 _22443_ (.A(_12444_),
    .B(_10749_),
    .Y(_12446_));
 sky130_fd_sc_hd__nand2_1 _22444_ (.A(_12445_),
    .B(_12446_),
    .Y(_12448_));
 sky130_fd_sc_hd__inv_4 _22445_ (.A(_12448_),
    .Y(_12449_));
 sky130_fd_sc_hd__nand2_1 _22446_ (.A(_12398_),
    .B(_11822_),
    .Y(_12450_));
 sky130_fd_sc_hd__inv_2 _22447_ (.A(_11813_),
    .Y(_12451_));
 sky130_fd_sc_hd__nand2_1 _22448_ (.A(_12450_),
    .B(_12451_),
    .Y(_12452_));
 sky130_fd_sc_hd__nand3_1 _22449_ (.A(_12398_),
    .B(_11822_),
    .C(_11813_),
    .Y(_12453_));
 sky130_fd_sc_hd__nand2_1 _22450_ (.A(_12452_),
    .B(_12453_),
    .Y(_12454_));
 sky130_fd_sc_hd__nand2_1 _22451_ (.A(_12454_),
    .B(_08001_),
    .Y(_12455_));
 sky130_fd_sc_hd__nand3_2 _22452_ (.A(_12452_),
    .B(_11858_),
    .C(_12453_),
    .Y(_12456_));
 sky130_fd_sc_hd__nand3_1 _22453_ (.A(_12406_),
    .B(_12455_),
    .C(_12456_),
    .Y(_12457_));
 sky130_fd_sc_hd__inv_2 _22454_ (.A(_12457_),
    .Y(_12459_));
 sky130_fd_sc_hd__nand3_1 _22455_ (.A(_12372_),
    .B(_12415_),
    .C(_12459_),
    .Y(_12460_));
 sky130_fd_sc_hd__inv_2 _22456_ (.A(_12402_),
    .Y(_12461_));
 sky130_fd_sc_hd__inv_2 _22457_ (.A(_12456_),
    .Y(_12462_));
 sky130_fd_sc_hd__a21o_1 _22458_ (.A1(_12455_),
    .A2(_12461_),
    .B1(_12462_),
    .X(_12463_));
 sky130_fd_sc_hd__nor2_1 _22459_ (.A(_12418_),
    .B(_12457_),
    .Y(_12464_));
 sky130_fd_sc_hd__nor2_1 _22460_ (.A(_12463_),
    .B(_12464_),
    .Y(_12465_));
 sky130_fd_sc_hd__nand2_1 _22461_ (.A(_12460_),
    .B(_12465_),
    .Y(_12466_));
 sky130_fd_sc_hd__or2_1 _22462_ (.A(_12449_),
    .B(_12466_),
    .X(_12467_));
 sky130_fd_sc_hd__nand2_1 _22463_ (.A(_12466_),
    .B(_12449_),
    .Y(_12468_));
 sky130_fd_sc_hd__nand2_1 _22464_ (.A(_12467_),
    .B(_12468_),
    .Y(_12470_));
 sky130_fd_sc_hd__nand2_1 _22465_ (.A(_12470_),
    .B(_12374_),
    .Y(_12471_));
 sky130_fd_sc_hd__nand2_1 _22466_ (.A(\div1i.quot[8] ),
    .B(_12444_),
    .Y(_12472_));
 sky130_fd_sc_hd__nand2_1 _22467_ (.A(_12471_),
    .B(_12472_),
    .Y(_12473_));
 sky130_fd_sc_hd__nand2_1 _22468_ (.A(_12473_),
    .B(_08020_),
    .Y(_12474_));
 sky130_fd_sc_hd__nand3_1 _22469_ (.A(_12471_),
    .B(_09664_),
    .C(_12472_),
    .Y(_12475_));
 sky130_fd_sc_hd__nand2_2 _22470_ (.A(_12474_),
    .B(_12475_),
    .Y(_12476_));
 sky130_fd_sc_hd__inv_2 _22471_ (.A(_12476_),
    .Y(_12477_));
 sky130_fd_sc_hd__nand2_1 _22472_ (.A(_12455_),
    .B(_12456_),
    .Y(_12478_));
 sky130_fd_sc_hd__nand2_1 _22473_ (.A(_12421_),
    .B(_12402_),
    .Y(_12479_));
 sky130_fd_sc_hd__xor2_1 _22474_ (.A(_12478_),
    .B(_12479_),
    .X(_12481_));
 sky130_fd_sc_hd__nand2_1 _22475_ (.A(_12481_),
    .B(_12374_),
    .Y(_12482_));
 sky130_fd_sc_hd__nand2_1 _22476_ (.A(_12454_),
    .B(\div1i.quot[8] ),
    .Y(_12483_));
 sky130_fd_sc_hd__nand2_1 _22477_ (.A(_12482_),
    .B(_12483_),
    .Y(_12484_));
 sky130_fd_sc_hd__nand2_1 _22478_ (.A(_12484_),
    .B(_11896_),
    .Y(_12485_));
 sky130_fd_sc_hd__nand3_2 _22479_ (.A(_12482_),
    .B(_11899_),
    .C(_12483_),
    .Y(_12486_));
 sky130_fd_sc_hd__nand3_1 _22480_ (.A(_12477_),
    .B(_12485_),
    .C(_12486_),
    .Y(_12487_));
 sky130_fd_sc_hd__nand2_1 _22481_ (.A(_12468_),
    .B(_12445_),
    .Y(_12488_));
 sky130_fd_sc_hd__nand2_1 _22482_ (.A(_12443_),
    .B(_11900_),
    .Y(_12489_));
 sky130_fd_sc_hd__or2_1 _22483_ (.A(_11889_),
    .B(_12489_),
    .X(_12490_));
 sky130_fd_sc_hd__nand2_1 _22484_ (.A(_12489_),
    .B(_11889_),
    .Y(_12492_));
 sky130_fd_sc_hd__nand2_1 _22485_ (.A(_12490_),
    .B(_12492_),
    .Y(_12493_));
 sky130_fd_sc_hd__nand2_1 _22486_ (.A(_12493_),
    .B(_08041_),
    .Y(_12494_));
 sky130_fd_sc_hd__buf_6 _22487_ (.A(_07461_),
    .X(_12495_));
 sky130_fd_sc_hd__nand3_1 _22488_ (.A(_12490_),
    .B(_12495_),
    .C(_12492_),
    .Y(_12496_));
 sky130_fd_sc_hd__nand2_1 _22489_ (.A(_12494_),
    .B(_12496_),
    .Y(_12497_));
 sky130_fd_sc_hd__inv_2 _22490_ (.A(_12497_),
    .Y(_12498_));
 sky130_fd_sc_hd__nand2_1 _22491_ (.A(_12488_),
    .B(_12498_),
    .Y(_12499_));
 sky130_fd_sc_hd__nand3_1 _22492_ (.A(_12468_),
    .B(_12497_),
    .C(_12445_),
    .Y(_12500_));
 sky130_fd_sc_hd__nand2_1 _22493_ (.A(_12499_),
    .B(_12500_),
    .Y(_12501_));
 sky130_fd_sc_hd__nand2_1 _22494_ (.A(_12501_),
    .B(_12374_),
    .Y(_12503_));
 sky130_fd_sc_hd__nand2_1 _22495_ (.A(_12493_),
    .B(\div1i.quot[8] ),
    .Y(_12504_));
 sky130_fd_sc_hd__nand2_1 _22496_ (.A(_12503_),
    .B(_12504_),
    .Y(_12505_));
 sky130_fd_sc_hd__buf_4 _22497_ (.A(_07474_),
    .X(_12506_));
 sky130_fd_sc_hd__nand2_1 _22498_ (.A(_12505_),
    .B(_12506_),
    .Y(_12507_));
 sky130_fd_sc_hd__nand3_1 _22499_ (.A(_12503_),
    .B(_11376_),
    .C(_12504_),
    .Y(_12508_));
 sky130_fd_sc_hd__nand2_1 _22500_ (.A(_12507_),
    .B(_12508_),
    .Y(_12509_));
 sky130_fd_sc_hd__inv_2 _22501_ (.A(_12509_),
    .Y(_12510_));
 sky130_fd_sc_hd__nand2_1 _22502_ (.A(_12498_),
    .B(_12449_),
    .Y(_12511_));
 sky130_fd_sc_hd__inv_2 _22503_ (.A(_12511_),
    .Y(_12512_));
 sky130_fd_sc_hd__nand2_1 _22504_ (.A(_12466_),
    .B(_12512_),
    .Y(_12514_));
 sky130_fd_sc_hd__o21a_1 _22505_ (.A1(_12445_),
    .A2(_12497_),
    .B1(_12496_),
    .X(_12515_));
 sky130_fd_sc_hd__nand2_1 _22506_ (.A(_12514_),
    .B(_12515_),
    .Y(_12516_));
 sky130_fd_sc_hd__a21oi_1 _22507_ (.A1(_11845_),
    .A2(_11849_),
    .B1(_11901_),
    .Y(_12517_));
 sky130_fd_sc_hd__or2_1 _22508_ (.A(_11956_),
    .B(_12517_),
    .X(_12518_));
 sky130_fd_sc_hd__or2_1 _22509_ (.A(_11921_),
    .B(_12518_),
    .X(_12519_));
 sky130_fd_sc_hd__nand2_1 _22510_ (.A(_12518_),
    .B(_11921_),
    .Y(_12520_));
 sky130_fd_sc_hd__nand2_1 _22511_ (.A(_12519_),
    .B(_12520_),
    .Y(_12521_));
 sky130_fd_sc_hd__inv_2 _22512_ (.A(_12521_),
    .Y(_12522_));
 sky130_fd_sc_hd__nand2_1 _22513_ (.A(_12522_),
    .B(_11935_),
    .Y(_12523_));
 sky130_fd_sc_hd__nand2_1 _22514_ (.A(_12521_),
    .B(_08611_),
    .Y(_12525_));
 sky130_fd_sc_hd__nand2_1 _22515_ (.A(_12523_),
    .B(_12525_),
    .Y(_12526_));
 sky130_fd_sc_hd__inv_2 _22516_ (.A(_12526_),
    .Y(_12527_));
 sky130_fd_sc_hd__nand2_1 _22517_ (.A(_12516_),
    .B(_12527_),
    .Y(_12528_));
 sky130_fd_sc_hd__nand3_1 _22518_ (.A(_12514_),
    .B(_12515_),
    .C(_12526_),
    .Y(_12529_));
 sky130_fd_sc_hd__nand3_1 _22519_ (.A(_12528_),
    .B(_12374_),
    .C(_12529_),
    .Y(_12530_));
 sky130_fd_sc_hd__nand2_1 _22520_ (.A(_12522_),
    .B(\div1i.quot[8] ),
    .Y(_12531_));
 sky130_fd_sc_hd__nand2_1 _22521_ (.A(_12530_),
    .B(_12531_),
    .Y(_12532_));
 sky130_fd_sc_hd__nand2_1 _22522_ (.A(_12532_),
    .B(_11946_),
    .Y(_12533_));
 sky130_fd_sc_hd__nand3_1 _22523_ (.A(_12530_),
    .B(_11948_),
    .C(_12531_),
    .Y(_12534_));
 sky130_fd_sc_hd__nand2_4 _22524_ (.A(_12533_),
    .B(_12534_),
    .Y(_12536_));
 sky130_fd_sc_hd__inv_2 _22525_ (.A(_12536_),
    .Y(_12537_));
 sky130_fd_sc_hd__nand2_1 _22526_ (.A(_12510_),
    .B(_12537_),
    .Y(_12538_));
 sky130_fd_sc_hd__nor2_1 _22527_ (.A(_12487_),
    .B(_12538_),
    .Y(_12539_));
 sky130_fd_sc_hd__nand2_4 _22528_ (.A(_12440_),
    .B(_12539_),
    .Y(_12540_));
 sky130_fd_sc_hd__o21ai_1 _22529_ (.A1(_12486_),
    .A2(_12476_),
    .B1(_12475_),
    .Y(_12541_));
 sky130_fd_sc_hd__nor2_1 _22530_ (.A(_12536_),
    .B(_12509_),
    .Y(_12542_));
 sky130_fd_sc_hd__o21ai_1 _22531_ (.A1(_12508_),
    .A2(_12536_),
    .B1(_12533_),
    .Y(_12543_));
 sky130_fd_sc_hd__a21oi_2 _22532_ (.A1(_12541_),
    .A2(_12542_),
    .B1(_12543_),
    .Y(_12544_));
 sky130_fd_sc_hd__nand2_4 _22533_ (.A(_12540_),
    .B(_12544_),
    .Y(_12545_));
 sky130_fd_sc_hd__nand2_2 _22534_ (.A(_12520_),
    .B(_11918_),
    .Y(_12547_));
 sky130_fd_sc_hd__xor2_4 _22535_ (.A(_11950_),
    .B(_12547_),
    .X(_12548_));
 sky130_fd_sc_hd__nand3_2 _22536_ (.A(_12528_),
    .B(_12374_),
    .C(_12523_),
    .Y(_12549_));
 sky130_fd_sc_hd__xnor2_4 _22537_ (.A(_12548_),
    .B(_12549_),
    .Y(_12550_));
 sky130_fd_sc_hd__nand2_8 _22538_ (.A(_12545_),
    .B(_12550_),
    .Y(_12551_));
 sky130_fd_sc_hd__inv_2 _22539_ (.A(_12550_),
    .Y(_12552_));
 sky130_fd_sc_hd__nand3_4 _22540_ (.A(_12540_),
    .B(_12544_),
    .C(_12552_),
    .Y(_12553_));
 sky130_fd_sc_hd__nand2_8 _22541_ (.A(_12551_),
    .B(_12553_),
    .Y(_12554_));
 sky130_fd_sc_hd__buf_8 _22542_ (.A(_12554_),
    .X(_12555_));
 sky130_fd_sc_hd__buf_8 _22543_ (.A(net223),
    .X(\div1i.quot[7] ));
 sky130_fd_sc_hd__nand2_1 _22544_ (.A(_12217_),
    .B(_12220_),
    .Y(_12557_));
 sky130_fd_sc_hd__nand2_1 _22545_ (.A(_12557_),
    .B(_12222_),
    .Y(_12558_));
 sky130_fd_sc_hd__nand2_1 _22546_ (.A(_12558_),
    .B(_12224_),
    .Y(_12559_));
 sky130_fd_sc_hd__inv_2 _22547_ (.A(_12559_),
    .Y(_12560_));
 sky130_fd_sc_hd__nand2_1 _22548_ (.A(_12555_),
    .B(_12560_),
    .Y(_12561_));
 sky130_fd_sc_hd__o21ai_2 _22549_ (.A1(_12032_),
    .A2(\div1i.quot[8] ),
    .B1(_12033_),
    .Y(_12562_));
 sky130_fd_sc_hd__nand2_1 _22550_ (.A(_12559_),
    .B(_12030_),
    .Y(_12563_));
 sky130_fd_sc_hd__nand3_1 _22551_ (.A(_12558_),
    .B(_12035_),
    .C(_12224_),
    .Y(_12564_));
 sky130_fd_sc_hd__nand2_1 _22552_ (.A(_12563_),
    .B(_12564_),
    .Y(_12565_));
 sky130_fd_sc_hd__xor2_1 _22553_ (.A(_12562_),
    .B(_12565_),
    .X(_12566_));
 sky130_fd_sc_hd__nand3b_1 _22554_ (.A_N(_12566_),
    .B(_12551_),
    .C(_12553_),
    .Y(_12568_));
 sky130_fd_sc_hd__nand2_1 _22555_ (.A(_12561_),
    .B(_12568_),
    .Y(_12569_));
 sky130_fd_sc_hd__nand2_2 _22556_ (.A(_12569_),
    .B(_11069_),
    .Y(_12570_));
 sky130_fd_sc_hd__nor2_1 _22557_ (.A(_12032_),
    .B(_12374_),
    .Y(_12571_));
 sky130_fd_sc_hd__or2_1 _22558_ (.A(_11412_),
    .B(_12571_),
    .X(_12572_));
 sky130_fd_sc_hd__nand2_1 _22559_ (.A(_12572_),
    .B(_12222_),
    .Y(_12573_));
 sky130_fd_sc_hd__inv_2 _22560_ (.A(_12573_),
    .Y(_12574_));
 sky130_fd_sc_hd__nand2_2 _22561_ (.A(_12555_),
    .B(_12574_),
    .Y(_12575_));
 sky130_fd_sc_hd__nand3_1 _22562_ (.A(_12551_),
    .B(_12553_),
    .C(_12571_),
    .Y(_12576_));
 sky130_fd_sc_hd__nand2_2 _22563_ (.A(_12575_),
    .B(_12576_),
    .Y(_12577_));
 sky130_fd_sc_hd__nand2_4 _22564_ (.A(_12577_),
    .B(_11421_),
    .Y(_12579_));
 sky130_fd_sc_hd__nand2_2 _22565_ (.A(_12570_),
    .B(_12579_),
    .Y(_12580_));
 sky130_fd_sc_hd__inv_2 _22566_ (.A(_12580_),
    .Y(_12581_));
 sky130_fd_sc_hd__nand3_2 _22567_ (.A(_12575_),
    .B(_11426_),
    .C(_12576_),
    .Y(_12582_));
 sky130_fd_sc_hd__nand3_2 _22568_ (.A(_12555_),
    .B(_12033_),
    .C(_12221_),
    .Y(_12583_));
 sky130_fd_sc_hd__inv_2 _22569_ (.A(_12583_),
    .Y(_12584_));
 sky130_fd_sc_hd__nand3_4 _22570_ (.A(_12579_),
    .B(_12582_),
    .C(_12584_),
    .Y(_12585_));
 sky130_fd_sc_hd__or2_4 _22571_ (.A(_11069_),
    .B(_12569_),
    .X(_12586_));
 sky130_fd_sc_hd__inv_2 _22572_ (.A(_12586_),
    .Y(_12587_));
 sky130_fd_sc_hd__a21oi_1 _22573_ (.A1(_12581_),
    .A2(_12585_),
    .B1(_12587_),
    .Y(_12588_));
 sky130_fd_sc_hd__nand2_1 _22574_ (.A(_12219_),
    .B(_12224_),
    .Y(_12590_));
 sky130_fd_sc_hd__nand2_1 _22575_ (.A(_12590_),
    .B(_12225_),
    .Y(_12591_));
 sky130_fd_sc_hd__inv_2 _22576_ (.A(_12280_),
    .Y(_12592_));
 sky130_fd_sc_hd__o21ai_1 _22577_ (.A1(_12276_),
    .A2(_12591_),
    .B1(_12592_),
    .Y(_12593_));
 sky130_fd_sc_hd__or2_1 _22578_ (.A(_12250_),
    .B(_12593_),
    .X(_12594_));
 sky130_fd_sc_hd__nand2_1 _22579_ (.A(_12593_),
    .B(_12250_),
    .Y(_12595_));
 sky130_fd_sc_hd__nand2_1 _22580_ (.A(_12594_),
    .B(_12595_),
    .Y(_12596_));
 sky130_fd_sc_hd__inv_2 _22581_ (.A(_12596_),
    .Y(_12597_));
 sky130_fd_sc_hd__nand2_1 _22582_ (.A(_12554_),
    .B(_12597_),
    .Y(_12598_));
 sky130_fd_sc_hd__nand2_1 _22583_ (.A(_12597_),
    .B(_12087_),
    .Y(_12599_));
 sky130_fd_sc_hd__nand2_1 _22584_ (.A(_12596_),
    .B(_12085_),
    .Y(_12601_));
 sky130_fd_sc_hd__nand2_1 _22585_ (.A(_12599_),
    .B(_12601_),
    .Y(_12602_));
 sky130_fd_sc_hd__inv_2 _22586_ (.A(_12602_),
    .Y(_12603_));
 sky130_fd_sc_hd__nand2_1 _22587_ (.A(_12226_),
    .B(_12275_),
    .Y(_12604_));
 sky130_fd_sc_hd__nand2_1 _22588_ (.A(_12591_),
    .B(_12274_),
    .Y(_12605_));
 sky130_fd_sc_hd__nand2_1 _22589_ (.A(_12604_),
    .B(_12605_),
    .Y(_12606_));
 sky130_fd_sc_hd__nand2_1 _22590_ (.A(_12606_),
    .B(_12056_),
    .Y(_12607_));
 sky130_fd_sc_hd__nand3_1 _22591_ (.A(_12604_),
    .B(_12058_),
    .C(_12605_),
    .Y(_12608_));
 sky130_fd_sc_hd__nand2_1 _22592_ (.A(_12607_),
    .B(_12608_),
    .Y(_12609_));
 sky130_fd_sc_hd__inv_2 _22593_ (.A(_12609_),
    .Y(_12610_));
 sky130_fd_sc_hd__inv_2 _22594_ (.A(_12564_),
    .Y(_12612_));
 sky130_fd_sc_hd__a21o_1 _22595_ (.A1(_12563_),
    .A2(_12562_),
    .B1(_12612_),
    .X(_12613_));
 sky130_fd_sc_hd__nand2_1 _22596_ (.A(_12225_),
    .B(_12208_),
    .Y(_12614_));
 sky130_fd_sc_hd__nand2_1 _22597_ (.A(_12224_),
    .B(_12217_),
    .Y(_12615_));
 sky130_fd_sc_hd__xor2_2 _22598_ (.A(_12614_),
    .B(_12615_),
    .X(_12616_));
 sky130_fd_sc_hd__nand2_1 _22599_ (.A(_12616_),
    .B(_12043_),
    .Y(_12617_));
 sky130_fd_sc_hd__nand2_1 _22600_ (.A(_12613_),
    .B(_12617_),
    .Y(_12618_));
 sky130_fd_sc_hd__inv_2 _22601_ (.A(_12616_),
    .Y(_12619_));
 sky130_fd_sc_hd__nand2_1 _22602_ (.A(_12619_),
    .B(_12047_),
    .Y(_12620_));
 sky130_fd_sc_hd__nand2_1 _22603_ (.A(_12618_),
    .B(_12620_),
    .Y(_12621_));
 sky130_fd_sc_hd__nand2_1 _22604_ (.A(_12610_),
    .B(_12621_),
    .Y(_12623_));
 sky130_fd_sc_hd__nand2_1 _22605_ (.A(_12623_),
    .B(_12608_),
    .Y(_12624_));
 sky130_fd_sc_hd__nand2_1 _22606_ (.A(_12604_),
    .B(_12272_),
    .Y(_12625_));
 sky130_fd_sc_hd__xor2_1 _22607_ (.A(_12263_),
    .B(_12625_),
    .X(_12626_));
 sky130_fd_sc_hd__nand2_1 _22608_ (.A(_12626_),
    .B(_09823_),
    .Y(_12627_));
 sky130_fd_sc_hd__nand2_1 _22609_ (.A(_12624_),
    .B(_12627_),
    .Y(_12628_));
 sky130_fd_sc_hd__inv_2 _22610_ (.A(_12626_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand2_1 _22611_ (.A(_12629_),
    .B(_08176_),
    .Y(_12630_));
 sky130_fd_sc_hd__nand2_1 _22612_ (.A(_12628_),
    .B(_12630_),
    .Y(_12631_));
 sky130_fd_sc_hd__or2_1 _22613_ (.A(_12603_),
    .B(_12631_),
    .X(_12632_));
 sky130_fd_sc_hd__nand2_1 _22614_ (.A(_12631_),
    .B(_12603_),
    .Y(_12634_));
 sky130_fd_sc_hd__nand2_1 _22615_ (.A(_12632_),
    .B(_12634_),
    .Y(_12635_));
 sky130_fd_sc_hd__inv_2 _22616_ (.A(_12635_),
    .Y(_12636_));
 sky130_fd_sc_hd__nand3_1 _22617_ (.A(_12551_),
    .B(_12553_),
    .C(_12636_),
    .Y(_12637_));
 sky130_fd_sc_hd__nand2_1 _22618_ (.A(_12598_),
    .B(_12637_),
    .Y(_12638_));
 sky130_fd_sc_hd__nand2_1 _22619_ (.A(_12638_),
    .B(_11482_),
    .Y(_12639_));
 sky130_fd_sc_hd__nand3_1 _22620_ (.A(_12598_),
    .B(_11484_),
    .C(_12637_),
    .Y(_12640_));
 sky130_fd_sc_hd__nand2_1 _22621_ (.A(_12639_),
    .B(_12640_),
    .Y(_12641_));
 sky130_fd_sc_hd__inv_2 _22622_ (.A(_12641_),
    .Y(_12642_));
 sky130_fd_sc_hd__nand2_1 _22623_ (.A(_12554_),
    .B(_12629_),
    .Y(_12643_));
 sky130_fd_sc_hd__nand2_1 _22624_ (.A(_12630_),
    .B(_12627_),
    .Y(_12645_));
 sky130_fd_sc_hd__xnor2_1 _22625_ (.A(_12624_),
    .B(_12645_),
    .Y(_12646_));
 sky130_fd_sc_hd__nand3_1 _22626_ (.A(_12551_),
    .B(_12553_),
    .C(_12646_),
    .Y(_12647_));
 sky130_fd_sc_hd__nand2_1 _22627_ (.A(_12643_),
    .B(_12647_),
    .Y(_12648_));
 sky130_fd_sc_hd__nand2_1 _22628_ (.A(_12648_),
    .B(_11494_),
    .Y(_12649_));
 sky130_fd_sc_hd__nand3_1 _22629_ (.A(_12643_),
    .B(_11496_),
    .C(_12647_),
    .Y(_12650_));
 sky130_fd_sc_hd__nand2_2 _22630_ (.A(_12649_),
    .B(_12650_),
    .Y(_12651_));
 sky130_fd_sc_hd__inv_2 _22631_ (.A(_12651_),
    .Y(_12652_));
 sky130_fd_sc_hd__nand2_1 _22632_ (.A(_12642_),
    .B(_12652_),
    .Y(_12653_));
 sky130_fd_sc_hd__inv_2 _22633_ (.A(_12606_),
    .Y(_12654_));
 sky130_fd_sc_hd__nand2_1 _22634_ (.A(_12554_),
    .B(_12654_),
    .Y(_12656_));
 sky130_fd_sc_hd__or2_1 _22635_ (.A(_12621_),
    .B(_12610_),
    .X(_12657_));
 sky130_fd_sc_hd__nand2_1 _22636_ (.A(_12657_),
    .B(_12623_),
    .Y(_12658_));
 sky130_fd_sc_hd__clkinvlp_2 _22637_ (.A(_12658_),
    .Y(_12659_));
 sky130_fd_sc_hd__nand3_1 _22638_ (.A(_12551_),
    .B(_12553_),
    .C(_12659_),
    .Y(_12660_));
 sky130_fd_sc_hd__nand2_1 _22639_ (.A(_12656_),
    .B(_12660_),
    .Y(_12661_));
 sky130_fd_sc_hd__nand2_1 _22640_ (.A(_12661_),
    .B(_11105_),
    .Y(_12662_));
 sky130_fd_sc_hd__nand3_1 _22641_ (.A(_12656_),
    .B(_12261_),
    .C(_12660_),
    .Y(_12663_));
 sky130_fd_sc_hd__nand2_2 _22642_ (.A(_12662_),
    .B(_12663_),
    .Y(_12664_));
 sky130_fd_sc_hd__inv_2 _22643_ (.A(_12664_),
    .Y(_12665_));
 sky130_fd_sc_hd__nand2_1 _22644_ (.A(_12554_),
    .B(_12619_),
    .Y(_12667_));
 sky130_fd_sc_hd__nand2_1 _22645_ (.A(_12620_),
    .B(_12617_),
    .Y(_12668_));
 sky130_fd_sc_hd__xnor2_1 _22646_ (.A(_12613_),
    .B(_12668_),
    .Y(_12669_));
 sky130_fd_sc_hd__nand3_1 _22647_ (.A(_12551_),
    .B(_12553_),
    .C(_12669_),
    .Y(_12670_));
 sky130_fd_sc_hd__nand2_1 _22648_ (.A(_12667_),
    .B(_12670_),
    .Y(_12671_));
 sky130_fd_sc_hd__nand2_1 _22649_ (.A(_12671_),
    .B(_12270_),
    .Y(_12672_));
 sky130_fd_sc_hd__nand3_1 _22650_ (.A(_12667_),
    .B(_11117_),
    .C(_12670_),
    .Y(_12673_));
 sky130_fd_sc_hd__nand2_1 _22651_ (.A(_12672_),
    .B(_12673_),
    .Y(_12674_));
 sky130_fd_sc_hd__inv_2 _22652_ (.A(_12674_),
    .Y(_12675_));
 sky130_fd_sc_hd__nand2_1 _22653_ (.A(_12665_),
    .B(_12675_),
    .Y(_12676_));
 sky130_fd_sc_hd__nor2_1 _22654_ (.A(_12653_),
    .B(_12676_),
    .Y(_12678_));
 sky130_fd_sc_hd__nand2_1 _22655_ (.A(_12588_),
    .B(_12678_),
    .Y(_12679_));
 sky130_fd_sc_hd__inv_2 _22656_ (.A(_12663_),
    .Y(_12680_));
 sky130_fd_sc_hd__o21ai_2 _22657_ (.A1(_12672_),
    .A2(_12680_),
    .B1(_12662_),
    .Y(_12681_));
 sky130_fd_sc_hd__nor2_1 _22658_ (.A(_12641_),
    .B(_12651_),
    .Y(_12682_));
 sky130_fd_sc_hd__inv_2 _22659_ (.A(_12640_),
    .Y(_12683_));
 sky130_fd_sc_hd__o21ai_1 _22660_ (.A1(_12649_),
    .A2(_12683_),
    .B1(_12639_),
    .Y(_12684_));
 sky130_fd_sc_hd__a21oi_1 _22661_ (.A1(_12681_),
    .A2(_12682_),
    .B1(_12684_),
    .Y(_12685_));
 sky130_fd_sc_hd__nand2_2 _22662_ (.A(_12679_),
    .B(_12685_),
    .Y(_12686_));
 sky130_fd_sc_hd__inv_2 _22663_ (.A(_12308_),
    .Y(_12687_));
 sky130_fd_sc_hd__nand2_1 _22664_ (.A(_12286_),
    .B(_12687_),
    .Y(_12689_));
 sky130_fd_sc_hd__inv_2 _22665_ (.A(_12332_),
    .Y(_12690_));
 sky130_fd_sc_hd__nand2_1 _22666_ (.A(_12689_),
    .B(_12690_),
    .Y(_12691_));
 sky130_fd_sc_hd__inv_2 _22667_ (.A(_12319_),
    .Y(_12692_));
 sky130_fd_sc_hd__nand2_1 _22668_ (.A(_12691_),
    .B(_12692_),
    .Y(_12693_));
 sky130_fd_sc_hd__nand3_1 _22669_ (.A(_12689_),
    .B(_12319_),
    .C(_12690_),
    .Y(_12694_));
 sky130_fd_sc_hd__nand2_1 _22670_ (.A(_12693_),
    .B(_12694_),
    .Y(_12695_));
 sky130_fd_sc_hd__inv_2 _22671_ (.A(_12695_),
    .Y(_12696_));
 sky130_fd_sc_hd__nand2_1 _22672_ (.A(_12696_),
    .B(_11986_),
    .Y(_12697_));
 sky130_fd_sc_hd__nand2_1 _22673_ (.A(_12695_),
    .B(_12017_),
    .Y(_12698_));
 sky130_fd_sc_hd__nand2_1 _22674_ (.A(_12697_),
    .B(_12698_),
    .Y(_12700_));
 sky130_fd_sc_hd__inv_2 _22675_ (.A(_12700_),
    .Y(_12701_));
 sky130_fd_sc_hd__nand2_1 _22676_ (.A(_12595_),
    .B(_12247_),
    .Y(_12702_));
 sky130_fd_sc_hd__or2_1 _22677_ (.A(_12240_),
    .B(_12702_),
    .X(_12703_));
 sky130_fd_sc_hd__nand2_1 _22678_ (.A(_12702_),
    .B(_12240_),
    .Y(_12704_));
 sky130_fd_sc_hd__nand3_1 _22679_ (.A(_12703_),
    .B(_10939_),
    .C(_12704_),
    .Y(_12705_));
 sky130_fd_sc_hd__nand2_1 _22680_ (.A(_12705_),
    .B(_12599_),
    .Y(_12706_));
 sky130_fd_sc_hd__inv_2 _22681_ (.A(_12706_),
    .Y(_12707_));
 sky130_fd_sc_hd__nand2_2 _22682_ (.A(_12634_),
    .B(_12707_),
    .Y(_12708_));
 sky130_fd_sc_hd__nand2_2 _22683_ (.A(_12286_),
    .B(_12307_),
    .Y(_12709_));
 sky130_fd_sc_hd__nand2_2 _22684_ (.A(_12709_),
    .B(_12305_),
    .Y(_12711_));
 sky130_fd_sc_hd__xor2_1 _22685_ (.A(_12295_),
    .B(_12711_),
    .X(_12712_));
 sky130_fd_sc_hd__nand2_2 _22686_ (.A(_12712_),
    .B(_12002_),
    .Y(_12713_));
 sky130_fd_sc_hd__or2_1 _22687_ (.A(_12296_),
    .B(_12711_),
    .X(_12714_));
 sky130_fd_sc_hd__nand2_1 _22688_ (.A(_12711_),
    .B(_12296_),
    .Y(_12715_));
 sky130_fd_sc_hd__nand3_1 _22689_ (.A(_12714_),
    .B(_12012_),
    .C(_12715_),
    .Y(_12716_));
 sky130_fd_sc_hd__or2_1 _22690_ (.A(_12307_),
    .B(_12286_),
    .X(_12717_));
 sky130_fd_sc_hd__nand2_1 _22691_ (.A(_12717_),
    .B(_12709_),
    .Y(_12718_));
 sky130_fd_sc_hd__nand2_1 _22692_ (.A(_12718_),
    .B(_12101_),
    .Y(_12719_));
 sky130_fd_sc_hd__nand3_2 _22693_ (.A(_12717_),
    .B(_12008_),
    .C(_12709_),
    .Y(_12720_));
 sky130_fd_sc_hd__nand2_1 _22694_ (.A(_12719_),
    .B(_12720_),
    .Y(_12722_));
 sky130_fd_sc_hd__inv_2 _22695_ (.A(_12722_),
    .Y(_12723_));
 sky130_fd_sc_hd__nand3_1 _22696_ (.A(_12713_),
    .B(_12716_),
    .C(_12723_),
    .Y(_12724_));
 sky130_fd_sc_hd__inv_2 _22697_ (.A(_12724_),
    .Y(_12725_));
 sky130_fd_sc_hd__nand2_1 _22698_ (.A(_12703_),
    .B(_12704_),
    .Y(_12726_));
 sky130_fd_sc_hd__nand2_1 _22699_ (.A(_12726_),
    .B(_08738_),
    .Y(_12727_));
 sky130_fd_sc_hd__nand3_2 _22700_ (.A(_12708_),
    .B(_12725_),
    .C(_12727_),
    .Y(_12728_));
 sky130_fd_sc_hd__inv_2 _22701_ (.A(_12720_),
    .Y(_12729_));
 sky130_fd_sc_hd__a21boi_2 _22702_ (.A1(_12713_),
    .A2(_12729_),
    .B1_N(_12716_),
    .Y(_12730_));
 sky130_fd_sc_hd__nand2_1 _22703_ (.A(_12728_),
    .B(_12730_),
    .Y(_12731_));
 sky130_fd_sc_hd__or2_1 _22704_ (.A(_12701_),
    .B(_12731_),
    .X(_12733_));
 sky130_fd_sc_hd__inv_6 _22705_ (.A(_12554_),
    .Y(_12734_));
 sky130_fd_sc_hd__nand2_1 _22706_ (.A(_12731_),
    .B(_12701_),
    .Y(_12735_));
 sky130_fd_sc_hd__nand3_1 _22707_ (.A(_12733_),
    .B(_12734_),
    .C(_12735_),
    .Y(_12736_));
 sky130_fd_sc_hd__nand2_1 _22708_ (.A(net223),
    .B(_12696_),
    .Y(_12737_));
 sky130_fd_sc_hd__nand2_1 _22709_ (.A(_12736_),
    .B(_12737_),
    .Y(_12738_));
 sky130_fd_sc_hd__nand2_1 _22710_ (.A(_12738_),
    .B(_11586_),
    .Y(_12739_));
 sky130_fd_sc_hd__nand3_1 _22711_ (.A(_12736_),
    .B(_11588_),
    .C(_12737_),
    .Y(_12740_));
 sky130_fd_sc_hd__nand2_2 _22712_ (.A(_12739_),
    .B(_12740_),
    .Y(_12741_));
 sky130_fd_sc_hd__nand3_1 _22713_ (.A(_12708_),
    .B(_12727_),
    .C(_12723_),
    .Y(_12742_));
 sky130_fd_sc_hd__nand2_1 _22714_ (.A(_12742_),
    .B(_12720_),
    .Y(_12744_));
 sky130_fd_sc_hd__nand3_1 _22715_ (.A(_12744_),
    .B(_12716_),
    .C(_12713_),
    .Y(_12745_));
 sky130_fd_sc_hd__nand2_1 _22716_ (.A(_12713_),
    .B(_12716_),
    .Y(_12746_));
 sky130_fd_sc_hd__nand3_1 _22717_ (.A(_12742_),
    .B(_12746_),
    .C(_12720_),
    .Y(_12747_));
 sky130_fd_sc_hd__a21o_1 _22718_ (.A1(_12745_),
    .A2(_12747_),
    .B1(_12555_),
    .X(_12748_));
 sky130_fd_sc_hd__nand2_2 _22719_ (.A(net223),
    .B(_12712_),
    .Y(_12749_));
 sky130_fd_sc_hd__nand2_1 _22720_ (.A(_12748_),
    .B(_12749_),
    .Y(_12750_));
 sky130_fd_sc_hd__nand2_1 _22721_ (.A(_12750_),
    .B(_11600_),
    .Y(_12751_));
 sky130_fd_sc_hd__nand3_2 _22722_ (.A(_12748_),
    .B(_11603_),
    .C(_12749_),
    .Y(_12752_));
 sky130_fd_sc_hd__nand2_2 _22723_ (.A(_12751_),
    .B(_12752_),
    .Y(_12753_));
 sky130_fd_sc_hd__nor2_2 _22724_ (.A(_12741_),
    .B(_12753_),
    .Y(_12755_));
 sky130_fd_sc_hd__a21o_1 _22725_ (.A1(_12708_),
    .A2(_12727_),
    .B1(_12723_),
    .X(_12756_));
 sky130_fd_sc_hd__nand3_1 _22726_ (.A(_12734_),
    .B(_12742_),
    .C(_12756_),
    .Y(_12757_));
 sky130_fd_sc_hd__a21o_1 _22727_ (.A1(_12551_),
    .A2(_12553_),
    .B1(_12718_),
    .X(_12758_));
 sky130_fd_sc_hd__nand2_1 _22728_ (.A(_12757_),
    .B(_12758_),
    .Y(_12759_));
 sky130_fd_sc_hd__nand2_1 _22729_ (.A(_12759_),
    .B(_11614_),
    .Y(_12760_));
 sky130_fd_sc_hd__nand3_1 _22730_ (.A(_12757_),
    .B(_11616_),
    .C(_12758_),
    .Y(_12761_));
 sky130_fd_sc_hd__nand2_1 _22731_ (.A(_12760_),
    .B(_12761_),
    .Y(_12762_));
 sky130_fd_sc_hd__nand2_1 _22732_ (.A(_12727_),
    .B(_12705_),
    .Y(_12763_));
 sky130_fd_sc_hd__nand2_1 _22733_ (.A(_12634_),
    .B(_12599_),
    .Y(_12764_));
 sky130_fd_sc_hd__xor2_1 _22734_ (.A(_12763_),
    .B(_12764_),
    .X(_12766_));
 sky130_fd_sc_hd__nand2_1 _22735_ (.A(_12734_),
    .B(_12766_),
    .Y(_12767_));
 sky130_fd_sc_hd__nand2_1 _22736_ (.A(_12555_),
    .B(_12726_),
    .Y(_12768_));
 sky130_fd_sc_hd__nand2_1 _22737_ (.A(_12767_),
    .B(_12768_),
    .Y(_12769_));
 sky130_fd_sc_hd__or2_4 _22738_ (.A(_09410_),
    .B(_12769_),
    .X(_12770_));
 sky130_fd_sc_hd__buf_4 _22739_ (.A(_09410_),
    .X(_12771_));
 sky130_fd_sc_hd__nand2_1 _22740_ (.A(_12769_),
    .B(_12771_),
    .Y(_12772_));
 sky130_fd_sc_hd__nand2_1 _22741_ (.A(_12770_),
    .B(_12772_),
    .Y(_12773_));
 sky130_fd_sc_hd__nor2_1 _22742_ (.A(_12762_),
    .B(_12773_),
    .Y(_12774_));
 sky130_fd_sc_hd__nand2_1 _22743_ (.A(_12755_),
    .B(_12774_),
    .Y(_12775_));
 sky130_fd_sc_hd__inv_2 _22744_ (.A(_12775_),
    .Y(_12777_));
 sky130_fd_sc_hd__nand2_1 _22745_ (.A(_12686_),
    .B(_12777_),
    .Y(_12778_));
 sky130_fd_sc_hd__o21ai_1 _22746_ (.A1(_12770_),
    .A2(_12762_),
    .B1(_12760_),
    .Y(_12779_));
 sky130_fd_sc_hd__o21ai_1 _22747_ (.A1(_12752_),
    .A2(_12741_),
    .B1(_12739_),
    .Y(_12780_));
 sky130_fd_sc_hd__a21oi_1 _22748_ (.A1(_12779_),
    .A2(_12755_),
    .B1(_12780_),
    .Y(_12781_));
 sky130_fd_sc_hd__nand2_2 _22749_ (.A(_12781_),
    .B(_12778_),
    .Y(_12782_));
 sky130_fd_sc_hd__inv_2 _22750_ (.A(_12728_),
    .Y(_12783_));
 sky130_fd_sc_hd__nand2_1 _22751_ (.A(_12693_),
    .B(_12318_),
    .Y(_12784_));
 sky130_fd_sc_hd__inv_2 _22752_ (.A(_12327_),
    .Y(_12785_));
 sky130_fd_sc_hd__nand2_1 _22753_ (.A(_12784_),
    .B(_12785_),
    .Y(_12786_));
 sky130_fd_sc_hd__nand3_1 _22754_ (.A(_12693_),
    .B(_12327_),
    .C(_12318_),
    .Y(_12788_));
 sky130_fd_sc_hd__nand2_1 _22755_ (.A(_12786_),
    .B(_12788_),
    .Y(_12789_));
 sky130_fd_sc_hd__nand2_1 _22756_ (.A(_12789_),
    .B(_11983_),
    .Y(_12790_));
 sky130_fd_sc_hd__nand3_1 _22757_ (.A(_12786_),
    .B(_11990_),
    .C(_12788_),
    .Y(_12791_));
 sky130_fd_sc_hd__nand3_1 _22758_ (.A(_12701_),
    .B(_12790_),
    .C(_12791_),
    .Y(_12792_));
 sky130_fd_sc_hd__inv_2 _22759_ (.A(_12792_),
    .Y(_12793_));
 sky130_fd_sc_hd__nand2_1 _22760_ (.A(_12783_),
    .B(_12793_),
    .Y(_12794_));
 sky130_fd_sc_hd__nor2_1 _22761_ (.A(_12730_),
    .B(_12792_),
    .Y(_12795_));
 sky130_fd_sc_hd__nand2_1 _22762_ (.A(_12790_),
    .B(_12791_),
    .Y(_12796_));
 sky130_fd_sc_hd__o21ai_1 _22763_ (.A1(_12697_),
    .A2(_12796_),
    .B1(_12791_),
    .Y(_12797_));
 sky130_fd_sc_hd__nor2_1 _22764_ (.A(_12795_),
    .B(_12797_),
    .Y(_12799_));
 sky130_fd_sc_hd__nand2_1 _22765_ (.A(_12794_),
    .B(_12799_),
    .Y(_12800_));
 sky130_fd_sc_hd__inv_2 _22766_ (.A(_12341_),
    .Y(_12801_));
 sky130_fd_sc_hd__inv_2 _22767_ (.A(_12340_),
    .Y(_12802_));
 sky130_fd_sc_hd__nand2_1 _22768_ (.A(_12336_),
    .B(_12802_),
    .Y(_12803_));
 sky130_fd_sc_hd__nand2_1 _22769_ (.A(_12803_),
    .B(_12189_),
    .Y(_12804_));
 sky130_fd_sc_hd__or2_1 _22770_ (.A(_12801_),
    .B(_12804_),
    .X(_12805_));
 sky130_fd_sc_hd__nand2_1 _22771_ (.A(_12804_),
    .B(_12801_),
    .Y(_12806_));
 sky130_fd_sc_hd__nand2_1 _22772_ (.A(_12805_),
    .B(_12806_),
    .Y(_12807_));
 sky130_fd_sc_hd__nand2_1 _22773_ (.A(_12807_),
    .B(_12118_),
    .Y(_12808_));
 sky130_fd_sc_hd__nand3_1 _22774_ (.A(_12805_),
    .B(_12120_),
    .C(_12806_),
    .Y(_12810_));
 sky130_fd_sc_hd__nand2_1 _22775_ (.A(_12808_),
    .B(_12810_),
    .Y(_12811_));
 sky130_fd_sc_hd__inv_2 _22776_ (.A(_12811_),
    .Y(_12812_));
 sky130_fd_sc_hd__or2_1 _22777_ (.A(_12802_),
    .B(_12336_),
    .X(_12813_));
 sky130_fd_sc_hd__nand2_1 _22778_ (.A(_12813_),
    .B(_12803_),
    .Y(_12814_));
 sky130_fd_sc_hd__inv_2 _22779_ (.A(_12814_),
    .Y(_12815_));
 sky130_fd_sc_hd__nand2_1 _22780_ (.A(_12815_),
    .B(_11671_),
    .Y(_12816_));
 sky130_fd_sc_hd__buf_6 _22781_ (.A(_07677_),
    .X(_12817_));
 sky130_fd_sc_hd__nand2_1 _22782_ (.A(_12814_),
    .B(_12817_),
    .Y(_12818_));
 sky130_fd_sc_hd__nand2_1 _22783_ (.A(_12816_),
    .B(_12818_),
    .Y(_12819_));
 sky130_fd_sc_hd__inv_4 _22784_ (.A(_12819_),
    .Y(_12821_));
 sky130_fd_sc_hd__nand2_1 _22785_ (.A(_12812_),
    .B(_12821_),
    .Y(_12822_));
 sky130_fd_sc_hd__inv_2 _22786_ (.A(_12822_),
    .Y(_12823_));
 sky130_fd_sc_hd__nand2_1 _22787_ (.A(_12800_),
    .B(_12823_),
    .Y(_12824_));
 sky130_fd_sc_hd__inv_2 _22788_ (.A(_12816_),
    .Y(_12825_));
 sky130_fd_sc_hd__a21boi_2 _22789_ (.A1(_12808_),
    .A2(_12825_),
    .B1_N(_12810_),
    .Y(_12826_));
 sky130_fd_sc_hd__nand2_1 _22790_ (.A(_12824_),
    .B(_12826_),
    .Y(_12827_));
 sky130_fd_sc_hd__nand2_1 _22791_ (.A(_12336_),
    .B(_12342_),
    .Y(_12828_));
 sky130_fd_sc_hd__inv_2 _22792_ (.A(_12197_),
    .Y(_12829_));
 sky130_fd_sc_hd__nand2_1 _22793_ (.A(_12828_),
    .B(_12829_),
    .Y(_12830_));
 sky130_fd_sc_hd__inv_2 _22794_ (.A(_12175_),
    .Y(_12832_));
 sky130_fd_sc_hd__nand2_1 _22795_ (.A(_12830_),
    .B(_12832_),
    .Y(_12833_));
 sky130_fd_sc_hd__nand3_1 _22796_ (.A(_12828_),
    .B(_12829_),
    .C(_12175_),
    .Y(_12834_));
 sky130_fd_sc_hd__nand2_1 _22797_ (.A(_12833_),
    .B(_12834_),
    .Y(_12835_));
 sky130_fd_sc_hd__nand2_1 _22798_ (.A(_12835_),
    .B(_12149_),
    .Y(_12836_));
 sky130_fd_sc_hd__nand3_1 _22799_ (.A(_12833_),
    .B(_12834_),
    .C(_12147_),
    .Y(_12837_));
 sky130_fd_sc_hd__nand2_1 _22800_ (.A(_12836_),
    .B(_12837_),
    .Y(_12838_));
 sky130_fd_sc_hd__inv_2 _22801_ (.A(_12838_),
    .Y(_12839_));
 sky130_fd_sc_hd__nand2_1 _22802_ (.A(_12827_),
    .B(_12839_),
    .Y(_12840_));
 sky130_fd_sc_hd__nand3_1 _22803_ (.A(_12824_),
    .B(_12838_),
    .C(_12826_),
    .Y(_12841_));
 sky130_fd_sc_hd__nand3_1 _22804_ (.A(_12840_),
    .B(_12734_),
    .C(_12841_),
    .Y(_12843_));
 sky130_fd_sc_hd__or2_1 _22805_ (.A(_12835_),
    .B(_12734_),
    .X(_12844_));
 sky130_fd_sc_hd__nand2_1 _22806_ (.A(_12843_),
    .B(_12844_),
    .Y(_12845_));
 sky130_fd_sc_hd__nand2_1 _22807_ (.A(_12845_),
    .B(_11701_),
    .Y(_12846_));
 sky130_fd_sc_hd__nand3_1 _22808_ (.A(_12843_),
    .B(_11703_),
    .C(_12844_),
    .Y(_12847_));
 sky130_fd_sc_hd__nand2_1 _22809_ (.A(_12846_),
    .B(_12847_),
    .Y(_12848_));
 sky130_fd_sc_hd__nand2_1 _22810_ (.A(_12800_),
    .B(_12821_),
    .Y(_12849_));
 sky130_fd_sc_hd__nand2_1 _22811_ (.A(_12849_),
    .B(_12816_),
    .Y(_12850_));
 sky130_fd_sc_hd__nand2_1 _22812_ (.A(_12850_),
    .B(_12812_),
    .Y(_12851_));
 sky130_fd_sc_hd__nand3_1 _22813_ (.A(_12849_),
    .B(_12811_),
    .C(_12816_),
    .Y(_12852_));
 sky130_fd_sc_hd__nand2_1 _22814_ (.A(_12851_),
    .B(_12852_),
    .Y(_12854_));
 sky130_fd_sc_hd__nand2_1 _22815_ (.A(_12854_),
    .B(_12734_),
    .Y(_12855_));
 sky130_fd_sc_hd__nand2_1 _22816_ (.A(\div1i.quot[7] ),
    .B(_12807_),
    .Y(_12856_));
 sky130_fd_sc_hd__nand2_1 _22817_ (.A(_12855_),
    .B(_12856_),
    .Y(_12857_));
 sky130_fd_sc_hd__nand2_1 _22818_ (.A(_12857_),
    .B(_11715_),
    .Y(_12858_));
 sky130_fd_sc_hd__nand3_2 _22819_ (.A(_12855_),
    .B(_11717_),
    .C(_12856_),
    .Y(_12859_));
 sky130_fd_sc_hd__nand2_2 _22820_ (.A(_12858_),
    .B(_12859_),
    .Y(_12860_));
 sky130_fd_sc_hd__nor2_2 _22821_ (.A(_12848_),
    .B(_12860_),
    .Y(_12861_));
 sky130_fd_sc_hd__or2_1 _22822_ (.A(_12821_),
    .B(_12800_),
    .X(_12862_));
 sky130_fd_sc_hd__nand3_1 _22823_ (.A(_12862_),
    .B(_12734_),
    .C(_12849_),
    .Y(_12863_));
 sky130_fd_sc_hd__nand2_1 _22824_ (.A(net223),
    .B(_12815_),
    .Y(_12865_));
 sky130_fd_sc_hd__nand2_1 _22825_ (.A(_12863_),
    .B(_12865_),
    .Y(_12866_));
 sky130_fd_sc_hd__nand2_1 _22826_ (.A(_12866_),
    .B(_06149_),
    .Y(_12867_));
 sky130_fd_sc_hd__nand3_1 _22827_ (.A(_12863_),
    .B(_09944_),
    .C(_12865_),
    .Y(_12868_));
 sky130_fd_sc_hd__nand2_1 _22828_ (.A(_12867_),
    .B(_12868_),
    .Y(_12869_));
 sky130_fd_sc_hd__nand2_1 _22829_ (.A(_12735_),
    .B(_12697_),
    .Y(_12870_));
 sky130_fd_sc_hd__xor2_1 _22830_ (.A(_12796_),
    .B(_12870_),
    .X(_12871_));
 sky130_fd_sc_hd__buf_6 _22831_ (.A(_12734_),
    .X(_12872_));
 sky130_fd_sc_hd__nand2_1 _22832_ (.A(_12871_),
    .B(_12872_),
    .Y(_12873_));
 sky130_fd_sc_hd__nand2_1 _22833_ (.A(\div1i.quot[7] ),
    .B(_12789_),
    .Y(_12874_));
 sky130_fd_sc_hd__nand2_1 _22834_ (.A(_12873_),
    .B(_12874_),
    .Y(_12876_));
 sky130_fd_sc_hd__nand2_1 _22835_ (.A(_12876_),
    .B(_11185_),
    .Y(_12877_));
 sky130_fd_sc_hd__nand3_1 _22836_ (.A(_12873_),
    .B(_12187_),
    .C(_12874_),
    .Y(_12878_));
 sky130_fd_sc_hd__nand2_1 _22837_ (.A(_12877_),
    .B(_12878_),
    .Y(_12879_));
 sky130_fd_sc_hd__nor2_2 _22838_ (.A(_12869_),
    .B(_12879_),
    .Y(_12880_));
 sky130_fd_sc_hd__nand2_1 _22839_ (.A(_12861_),
    .B(_12880_),
    .Y(_12881_));
 sky130_fd_sc_hd__inv_2 _22840_ (.A(_12881_),
    .Y(_12882_));
 sky130_fd_sc_hd__nand2_1 _22841_ (.A(_12782_),
    .B(_12882_),
    .Y(_12883_));
 sky130_fd_sc_hd__o21ai_1 _22842_ (.A1(_12878_),
    .A2(_12869_),
    .B1(_12867_),
    .Y(_12884_));
 sky130_fd_sc_hd__o21ai_1 _22843_ (.A1(_12859_),
    .A2(_12848_),
    .B1(_12846_),
    .Y(_12885_));
 sky130_fd_sc_hd__a21oi_1 _22844_ (.A1(_12861_),
    .A2(_12884_),
    .B1(_12885_),
    .Y(_12887_));
 sky130_fd_sc_hd__nand2_2 _22845_ (.A(_12883_),
    .B(_12887_),
    .Y(_12888_));
 sky130_fd_sc_hd__nand2_1 _22846_ (.A(_12833_),
    .B(_12174_),
    .Y(_12889_));
 sky130_fd_sc_hd__inv_2 _22847_ (.A(_12163_),
    .Y(_12890_));
 sky130_fd_sc_hd__nand2_1 _22848_ (.A(_12889_),
    .B(_12890_),
    .Y(_12891_));
 sky130_fd_sc_hd__nand3_1 _22849_ (.A(_12833_),
    .B(_12163_),
    .C(_12174_),
    .Y(_12892_));
 sky130_fd_sc_hd__nand2_1 _22850_ (.A(_12891_),
    .B(_12892_),
    .Y(_12893_));
 sky130_fd_sc_hd__buf_6 _22851_ (.A(_07905_),
    .X(_12894_));
 sky130_fd_sc_hd__nand2_1 _22852_ (.A(_12893_),
    .B(_12894_),
    .Y(_12895_));
 sky130_fd_sc_hd__nand3_1 _22853_ (.A(_12891_),
    .B(_11754_),
    .C(_12892_),
    .Y(_12896_));
 sky130_fd_sc_hd__nand3_1 _22854_ (.A(_12895_),
    .B(_12896_),
    .C(_12839_),
    .Y(_12898_));
 sky130_fd_sc_hd__nor2_1 _22855_ (.A(_12898_),
    .B(_12822_),
    .Y(_12899_));
 sky130_fd_sc_hd__nand2_1 _22856_ (.A(_12800_),
    .B(_12899_),
    .Y(_12900_));
 sky130_fd_sc_hd__nor2_1 _22857_ (.A(_12898_),
    .B(_12826_),
    .Y(_12901_));
 sky130_fd_sc_hd__nand2_1 _22858_ (.A(_12895_),
    .B(_12896_),
    .Y(_12902_));
 sky130_fd_sc_hd__o21ai_1 _22859_ (.A1(_12837_),
    .A2(_12902_),
    .B1(_12896_),
    .Y(_12903_));
 sky130_fd_sc_hd__nor2_1 _22860_ (.A(_12901_),
    .B(_12903_),
    .Y(_12904_));
 sky130_fd_sc_hd__nand2_1 _22861_ (.A(_12900_),
    .B(_12904_),
    .Y(_12905_));
 sky130_fd_sc_hd__clkinvlp_2 _22862_ (.A(_12379_),
    .Y(_12906_));
 sky130_fd_sc_hd__inv_2 _22863_ (.A(_12389_),
    .Y(_12907_));
 sky130_fd_sc_hd__nand2_1 _22864_ (.A(_12344_),
    .B(_12907_),
    .Y(_12909_));
 sky130_fd_sc_hd__nand2_1 _22865_ (.A(_12909_),
    .B(_12388_),
    .Y(_12910_));
 sky130_fd_sc_hd__or2_1 _22866_ (.A(_12906_),
    .B(_12910_),
    .X(_12911_));
 sky130_fd_sc_hd__nand2_1 _22867_ (.A(_12910_),
    .B(_12906_),
    .Y(_12912_));
 sky130_fd_sc_hd__nand2_1 _22868_ (.A(_12911_),
    .B(_12912_),
    .Y(_12913_));
 sky130_fd_sc_hd__buf_6 _22869_ (.A(_07957_),
    .X(_12914_));
 sky130_fd_sc_hd__nand2_1 _22870_ (.A(_12913_),
    .B(_12914_),
    .Y(_12915_));
 sky130_fd_sc_hd__nand3_1 _22871_ (.A(_12911_),
    .B(_11774_),
    .C(_12912_),
    .Y(_12916_));
 sky130_fd_sc_hd__nand2_1 _22872_ (.A(_12915_),
    .B(_12916_),
    .Y(_12917_));
 sky130_fd_sc_hd__or2_1 _22873_ (.A(_12907_),
    .B(_12344_),
    .X(_12918_));
 sky130_fd_sc_hd__nand2_1 _22874_ (.A(_12918_),
    .B(_12909_),
    .Y(_12920_));
 sky130_fd_sc_hd__inv_2 _22875_ (.A(_12920_),
    .Y(_12921_));
 sky130_fd_sc_hd__nand2_1 _22876_ (.A(_12921_),
    .B(_11199_),
    .Y(_12922_));
 sky130_fd_sc_hd__nand2_1 _22877_ (.A(_12920_),
    .B(_08465_),
    .Y(_12923_));
 sky130_fd_sc_hd__nand2_1 _22878_ (.A(_12922_),
    .B(_12923_),
    .Y(_12924_));
 sky130_fd_sc_hd__inv_2 _22879_ (.A(_12924_),
    .Y(_12925_));
 sky130_fd_sc_hd__nand2b_1 _22880_ (.A_N(_12917_),
    .B(_12925_),
    .Y(_12926_));
 sky130_fd_sc_hd__inv_4 _22881_ (.A(_12926_),
    .Y(_12927_));
 sky130_fd_sc_hd__nand2_1 _22882_ (.A(_12905_),
    .B(_12927_),
    .Y(_12928_));
 sky130_fd_sc_hd__inv_2 _22883_ (.A(_12922_),
    .Y(_12929_));
 sky130_fd_sc_hd__a21boi_2 _22884_ (.A1(_12915_),
    .A2(_12929_),
    .B1_N(_12916_),
    .Y(_12931_));
 sky130_fd_sc_hd__nand2_1 _22885_ (.A(_12928_),
    .B(_12931_),
    .Y(_12932_));
 sky130_fd_sc_hd__inv_2 _22886_ (.A(_12434_),
    .Y(_12933_));
 sky130_fd_sc_hd__nand2_1 _22887_ (.A(_12395_),
    .B(_12933_),
    .Y(_12934_));
 sky130_fd_sc_hd__nand3_1 _22888_ (.A(_12391_),
    .B(_12394_),
    .C(_12434_),
    .Y(_12935_));
 sky130_fd_sc_hd__nand2_1 _22889_ (.A(_12934_),
    .B(_12935_),
    .Y(_12936_));
 sky130_fd_sc_hd__inv_2 _22890_ (.A(_12936_),
    .Y(_12937_));
 sky130_fd_sc_hd__nand2_1 _22891_ (.A(_12937_),
    .B(_11797_),
    .Y(_12938_));
 sky130_fd_sc_hd__buf_6 _22892_ (.A(_07948_),
    .X(_12939_));
 sky130_fd_sc_hd__nand2_1 _22893_ (.A(_12936_),
    .B(_12939_),
    .Y(_12940_));
 sky130_fd_sc_hd__nand2_1 _22894_ (.A(_12938_),
    .B(_12940_),
    .Y(_12942_));
 sky130_fd_sc_hd__inv_2 _22895_ (.A(_12942_),
    .Y(_12943_));
 sky130_fd_sc_hd__nand2_1 _22896_ (.A(_12932_),
    .B(_12943_),
    .Y(_12944_));
 sky130_fd_sc_hd__nand3_1 _22897_ (.A(_12928_),
    .B(_12942_),
    .C(_12931_),
    .Y(_12945_));
 sky130_fd_sc_hd__nand3_1 _22898_ (.A(_12944_),
    .B(_12872_),
    .C(_12945_),
    .Y(_12946_));
 sky130_fd_sc_hd__nand2_1 _22899_ (.A(\div1i.quot[7] ),
    .B(_12937_),
    .Y(_12947_));
 sky130_fd_sc_hd__nand2_1 _22900_ (.A(_12946_),
    .B(_12947_),
    .Y(_12948_));
 sky130_fd_sc_hd__nand2_1 _22901_ (.A(_12948_),
    .B(_11808_),
    .Y(_12949_));
 sky130_fd_sc_hd__nand3_1 _22902_ (.A(_12946_),
    .B(_11811_),
    .C(_12947_),
    .Y(_12950_));
 sky130_fd_sc_hd__nand2_1 _22903_ (.A(_12949_),
    .B(_12950_),
    .Y(_12951_));
 sky130_fd_sc_hd__nand2_1 _22904_ (.A(_12905_),
    .B(_12925_),
    .Y(_12953_));
 sky130_fd_sc_hd__nand2_1 _22905_ (.A(_12953_),
    .B(_12922_),
    .Y(_12954_));
 sky130_fd_sc_hd__xor2_1 _22906_ (.A(_12917_),
    .B(_12954_),
    .X(_12955_));
 sky130_fd_sc_hd__nand2_1 _22907_ (.A(_12955_),
    .B(_12872_),
    .Y(_12956_));
 sky130_fd_sc_hd__nand2_1 _22908_ (.A(\div1i.quot[7] ),
    .B(_12913_),
    .Y(_12957_));
 sky130_fd_sc_hd__nand2_1 _22909_ (.A(_12956_),
    .B(_12957_),
    .Y(_12958_));
 sky130_fd_sc_hd__nand2_1 _22910_ (.A(_12958_),
    .B(_10173_),
    .Y(_12959_));
 sky130_fd_sc_hd__nand3_2 _22911_ (.A(_12956_),
    .B(_07400_),
    .C(_12957_),
    .Y(_12960_));
 sky130_fd_sc_hd__nand2_1 _22912_ (.A(_12959_),
    .B(_12960_),
    .Y(_12961_));
 sky130_fd_sc_hd__nor2_1 _22913_ (.A(_12951_),
    .B(_12961_),
    .Y(_12962_));
 sky130_fd_sc_hd__nand3_1 _22914_ (.A(_12900_),
    .B(_12924_),
    .C(_12904_),
    .Y(_12964_));
 sky130_fd_sc_hd__nand3_1 _22915_ (.A(_12953_),
    .B(_12734_),
    .C(_12964_),
    .Y(_12965_));
 sky130_fd_sc_hd__nand2_1 _22916_ (.A(net223),
    .B(_12921_),
    .Y(_12966_));
 sky130_fd_sc_hd__nand2_1 _22917_ (.A(_12965_),
    .B(_12966_),
    .Y(_12967_));
 sky130_fd_sc_hd__or2_1 _22918_ (.A(_10138_),
    .B(_12967_),
    .X(_12968_));
 sky130_fd_sc_hd__nand2_1 _22919_ (.A(_12967_),
    .B(_10138_),
    .Y(_12969_));
 sky130_fd_sc_hd__nand2_2 _22920_ (.A(_12968_),
    .B(_12969_),
    .Y(_12970_));
 sky130_fd_sc_hd__nand2_1 _22921_ (.A(_12840_),
    .B(_12837_),
    .Y(_12971_));
 sky130_fd_sc_hd__xor2_1 _22922_ (.A(_12902_),
    .B(_12971_),
    .X(_12972_));
 sky130_fd_sc_hd__nand2_1 _22923_ (.A(_12972_),
    .B(_12872_),
    .Y(_12973_));
 sky130_fd_sc_hd__nand2_1 _22924_ (.A(\div1i.quot[7] ),
    .B(_12893_),
    .Y(_12975_));
 sky130_fd_sc_hd__nand2_1 _22925_ (.A(_12973_),
    .B(_12975_),
    .Y(_12976_));
 sky130_fd_sc_hd__nand2_1 _22926_ (.A(_12976_),
    .B(_11838_),
    .Y(_12977_));
 sky130_fd_sc_hd__nand3_2 _22927_ (.A(_12973_),
    .B(_11840_),
    .C(_12975_),
    .Y(_12978_));
 sky130_fd_sc_hd__nand3b_1 _22928_ (.A_N(_12970_),
    .B(_12977_),
    .C(_12978_),
    .Y(_12979_));
 sky130_fd_sc_hd__inv_2 _22929_ (.A(_12979_),
    .Y(_12980_));
 sky130_fd_sc_hd__nand3_1 _22930_ (.A(_12888_),
    .B(_12962_),
    .C(_12980_),
    .Y(_12981_));
 sky130_fd_sc_hd__inv_2 _22931_ (.A(_12969_),
    .Y(_12982_));
 sky130_fd_sc_hd__o21bai_1 _22932_ (.A1(_12970_),
    .A2(_12978_),
    .B1_N(_12982_),
    .Y(_12983_));
 sky130_fd_sc_hd__o21ai_1 _22933_ (.A1(_12951_),
    .A2(_12960_),
    .B1(_12949_),
    .Y(_12984_));
 sky130_fd_sc_hd__a21oi_1 _22934_ (.A1(_12962_),
    .A2(_12983_),
    .B1(_12984_),
    .Y(_12985_));
 sky130_fd_sc_hd__nand2_2 _22935_ (.A(_12981_),
    .B(_12985_),
    .Y(_12986_));
 sky130_fd_sc_hd__nand2_1 _22936_ (.A(_12934_),
    .B(_12432_),
    .Y(_12987_));
 sky130_fd_sc_hd__inv_2 _22937_ (.A(_12426_),
    .Y(_12988_));
 sky130_fd_sc_hd__nand2_1 _22938_ (.A(_12987_),
    .B(_12988_),
    .Y(_12989_));
 sky130_fd_sc_hd__nand3_1 _22939_ (.A(_12934_),
    .B(_12426_),
    .C(_12432_),
    .Y(_12990_));
 sky130_fd_sc_hd__nand2_1 _22940_ (.A(_12989_),
    .B(_12990_),
    .Y(_12991_));
 sky130_fd_sc_hd__buf_6 _22941_ (.A(_08001_),
    .X(_12992_));
 sky130_fd_sc_hd__nand2_1 _22942_ (.A(_12991_),
    .B(_12992_),
    .Y(_12993_));
 sky130_fd_sc_hd__nand3_1 _22943_ (.A(_12989_),
    .B(_11858_),
    .C(_12990_),
    .Y(_12994_));
 sky130_fd_sc_hd__nand3_1 _22944_ (.A(_12943_),
    .B(_12993_),
    .C(_12994_),
    .Y(_12996_));
 sky130_fd_sc_hd__inv_2 _22945_ (.A(_12996_),
    .Y(_12997_));
 sky130_fd_sc_hd__nand3_2 _22946_ (.A(_12905_),
    .B(_12927_),
    .C(_12997_),
    .Y(_12998_));
 sky130_fd_sc_hd__inv_2 _22947_ (.A(_12993_),
    .Y(_12999_));
 sky130_fd_sc_hd__o21ai_1 _22948_ (.A1(_12938_),
    .A2(_12999_),
    .B1(_12994_),
    .Y(_13000_));
 sky130_fd_sc_hd__nor2_1 _22949_ (.A(_12931_),
    .B(_12996_),
    .Y(_13001_));
 sky130_fd_sc_hd__nor2_1 _22950_ (.A(_13000_),
    .B(_13001_),
    .Y(_13002_));
 sky130_fd_sc_hd__nand2_1 _22951_ (.A(_12998_),
    .B(_13002_),
    .Y(_13003_));
 sky130_fd_sc_hd__inv_2 _22952_ (.A(_12440_),
    .Y(_13004_));
 sky130_fd_sc_hd__nand2_1 _22953_ (.A(_12485_),
    .B(_12486_),
    .Y(_13005_));
 sky130_fd_sc_hd__nand2_1 _22954_ (.A(_13004_),
    .B(_13005_),
    .Y(_13007_));
 sky130_fd_sc_hd__inv_2 _22955_ (.A(_13005_),
    .Y(_13008_));
 sky130_fd_sc_hd__nand2_1 _22956_ (.A(_12440_),
    .B(_13008_),
    .Y(_13009_));
 sky130_fd_sc_hd__nand2_1 _22957_ (.A(_13007_),
    .B(_13009_),
    .Y(_13010_));
 sky130_fd_sc_hd__nand2_1 _22958_ (.A(_13010_),
    .B(_10749_),
    .Y(_13011_));
 sky130_fd_sc_hd__nand3_2 _22959_ (.A(_13007_),
    .B(_08554_),
    .C(_13009_),
    .Y(_13012_));
 sky130_fd_sc_hd__nand2_1 _22960_ (.A(_13011_),
    .B(_13012_),
    .Y(_13013_));
 sky130_fd_sc_hd__inv_2 _22961_ (.A(_13013_),
    .Y(_13014_));
 sky130_fd_sc_hd__nand2_1 _22962_ (.A(_13003_),
    .B(_13014_),
    .Y(_13015_));
 sky130_fd_sc_hd__nand3_1 _22963_ (.A(_12998_),
    .B(_13002_),
    .C(_13013_),
    .Y(_13016_));
 sky130_fd_sc_hd__nand3_1 _22964_ (.A(_13015_),
    .B(_12872_),
    .C(_13016_),
    .Y(_13018_));
 sky130_fd_sc_hd__or2_1 _22965_ (.A(_13010_),
    .B(_12734_),
    .X(_13019_));
 sky130_fd_sc_hd__nand2_1 _22966_ (.A(_13018_),
    .B(_13019_),
    .Y(_13020_));
 sky130_fd_sc_hd__or2_1 _22967_ (.A(_09664_),
    .B(_13020_),
    .X(_13021_));
 sky130_fd_sc_hd__buf_6 _22968_ (.A(_09664_),
    .X(_13022_));
 sky130_fd_sc_hd__nand2_1 _22969_ (.A(_13020_),
    .B(_13022_),
    .Y(_13023_));
 sky130_fd_sc_hd__nand2_1 _22970_ (.A(_13021_),
    .B(_13023_),
    .Y(_13024_));
 sky130_fd_sc_hd__inv_2 _22971_ (.A(_13024_),
    .Y(_13025_));
 sky130_fd_sc_hd__nand2_1 _22972_ (.A(_12993_),
    .B(_12994_),
    .Y(_13026_));
 sky130_fd_sc_hd__nand2_1 _22973_ (.A(_12944_),
    .B(_12938_),
    .Y(_13027_));
 sky130_fd_sc_hd__xor2_1 _22974_ (.A(_13026_),
    .B(_13027_),
    .X(_13029_));
 sky130_fd_sc_hd__nand2_1 _22975_ (.A(_13029_),
    .B(_12872_),
    .Y(_13030_));
 sky130_fd_sc_hd__nand2_1 _22976_ (.A(\div1i.quot[7] ),
    .B(_12991_),
    .Y(_13031_));
 sky130_fd_sc_hd__nand2_1 _22977_ (.A(_13030_),
    .B(_13031_),
    .Y(_13032_));
 sky130_fd_sc_hd__nand2_1 _22978_ (.A(_13032_),
    .B(_11896_),
    .Y(_13033_));
 sky130_fd_sc_hd__nand3_2 _22979_ (.A(_13030_),
    .B(_11899_),
    .C(_13031_),
    .Y(_13034_));
 sky130_fd_sc_hd__nand3_1 _22980_ (.A(_13025_),
    .B(_13033_),
    .C(_13034_),
    .Y(_13035_));
 sky130_fd_sc_hd__nand2_1 _22981_ (.A(_13015_),
    .B(_13012_),
    .Y(_13036_));
 sky130_fd_sc_hd__nand2_1 _22982_ (.A(_13009_),
    .B(_12486_),
    .Y(_13037_));
 sky130_fd_sc_hd__xor2_2 _22983_ (.A(_12476_),
    .B(_13037_),
    .X(_13038_));
 sky130_fd_sc_hd__inv_2 _22984_ (.A(_13038_),
    .Y(_13040_));
 sky130_fd_sc_hd__nand2_1 _22985_ (.A(_13040_),
    .B(_12495_),
    .Y(_13041_));
 sky130_fd_sc_hd__buf_6 _22986_ (.A(_08041_),
    .X(_13042_));
 sky130_fd_sc_hd__nand2_1 _22987_ (.A(_13038_),
    .B(_13042_),
    .Y(_13043_));
 sky130_fd_sc_hd__nand2_1 _22988_ (.A(_13041_),
    .B(_13043_),
    .Y(_13044_));
 sky130_fd_sc_hd__inv_2 _22989_ (.A(_13044_),
    .Y(_13045_));
 sky130_fd_sc_hd__nand2_1 _22990_ (.A(_13036_),
    .B(_13045_),
    .Y(_13046_));
 sky130_fd_sc_hd__nand3_1 _22991_ (.A(_13015_),
    .B(_13044_),
    .C(_13012_),
    .Y(_13047_));
 sky130_fd_sc_hd__nand2_1 _22992_ (.A(_13046_),
    .B(_13047_),
    .Y(_13048_));
 sky130_fd_sc_hd__nand2_1 _22993_ (.A(_13048_),
    .B(_12872_),
    .Y(_13049_));
 sky130_fd_sc_hd__nand2_1 _22994_ (.A(_13038_),
    .B(\div1i.quot[7] ),
    .Y(_13051_));
 sky130_fd_sc_hd__nand2_1 _22995_ (.A(_13049_),
    .B(_13051_),
    .Y(_13052_));
 sky130_fd_sc_hd__nand2_1 _22996_ (.A(_13052_),
    .B(_12506_),
    .Y(_13053_));
 sky130_fd_sc_hd__nand3_1 _22997_ (.A(_13049_),
    .B(_11376_),
    .C(_13051_),
    .Y(_13054_));
 sky130_fd_sc_hd__nand2_1 _22998_ (.A(_13053_),
    .B(_13054_),
    .Y(_13055_));
 sky130_fd_sc_hd__inv_2 _22999_ (.A(_13055_),
    .Y(_13056_));
 sky130_fd_sc_hd__nand3_1 _23000_ (.A(_13041_),
    .B(_13043_),
    .C(_13014_),
    .Y(_13057_));
 sky130_fd_sc_hd__inv_2 _23001_ (.A(_13057_),
    .Y(_13058_));
 sky130_fd_sc_hd__nand2_1 _23002_ (.A(_13058_),
    .B(_13003_),
    .Y(_13059_));
 sky130_fd_sc_hd__inv_2 _23003_ (.A(_13043_),
    .Y(_13060_));
 sky130_fd_sc_hd__o21a_1 _23004_ (.A1(_13012_),
    .A2(_13060_),
    .B1(_13041_),
    .X(_13062_));
 sky130_fd_sc_hd__nand2_1 _23005_ (.A(_13059_),
    .B(_13062_),
    .Y(_13063_));
 sky130_fd_sc_hd__o21bai_1 _23006_ (.A1(_12487_),
    .A2(_13004_),
    .B1_N(_12541_),
    .Y(_13064_));
 sky130_fd_sc_hd__or2_1 _23007_ (.A(_12510_),
    .B(_13064_),
    .X(_13065_));
 sky130_fd_sc_hd__nand2_1 _23008_ (.A(_13064_),
    .B(_12510_),
    .Y(_13066_));
 sky130_fd_sc_hd__nand2_1 _23009_ (.A(_13065_),
    .B(_13066_),
    .Y(_13067_));
 sky130_fd_sc_hd__inv_2 _23010_ (.A(_13067_),
    .Y(_13068_));
 sky130_fd_sc_hd__nand2_1 _23011_ (.A(_13068_),
    .B(_11935_),
    .Y(_13069_));
 sky130_fd_sc_hd__nand2_1 _23012_ (.A(_13067_),
    .B(_08611_),
    .Y(_13070_));
 sky130_fd_sc_hd__nand2_1 _23013_ (.A(_13069_),
    .B(_13070_),
    .Y(_13071_));
 sky130_fd_sc_hd__inv_2 _23014_ (.A(_13071_),
    .Y(_13073_));
 sky130_fd_sc_hd__nand2_1 _23015_ (.A(_13063_),
    .B(_13073_),
    .Y(_13074_));
 sky130_fd_sc_hd__nand3_1 _23016_ (.A(_13059_),
    .B(_13062_),
    .C(_13071_),
    .Y(_13075_));
 sky130_fd_sc_hd__nand3_1 _23017_ (.A(_13074_),
    .B(_13075_),
    .C(_12872_),
    .Y(_13076_));
 sky130_fd_sc_hd__nand2_1 _23018_ (.A(_13068_),
    .B(\div1i.quot[7] ),
    .Y(_13077_));
 sky130_fd_sc_hd__nand2_1 _23019_ (.A(_13076_),
    .B(_13077_),
    .Y(_13078_));
 sky130_fd_sc_hd__nand2_1 _23020_ (.A(_13078_),
    .B(_11946_),
    .Y(_13079_));
 sky130_fd_sc_hd__nand3_1 _23021_ (.A(_13076_),
    .B(_11948_),
    .C(_13077_),
    .Y(_13080_));
 sky130_fd_sc_hd__nand2_2 _23022_ (.A(_13079_),
    .B(_13080_),
    .Y(_13081_));
 sky130_fd_sc_hd__inv_2 _23023_ (.A(_13081_),
    .Y(_13082_));
 sky130_fd_sc_hd__nand2_1 _23024_ (.A(_13056_),
    .B(_13082_),
    .Y(_13084_));
 sky130_fd_sc_hd__nor2_1 _23025_ (.A(_13035_),
    .B(_13084_),
    .Y(_13085_));
 sky130_fd_sc_hd__nand2_4 _23026_ (.A(_12986_),
    .B(_13085_),
    .Y(_13086_));
 sky130_fd_sc_hd__o21ai_1 _23027_ (.A1(_13024_),
    .A2(_13034_),
    .B1(_13023_),
    .Y(_13087_));
 sky130_fd_sc_hd__nor2_1 _23028_ (.A(_13081_),
    .B(_13055_),
    .Y(_13088_));
 sky130_fd_sc_hd__inv_2 _23029_ (.A(_13080_),
    .Y(_13089_));
 sky130_fd_sc_hd__o21ai_1 _23030_ (.A1(_13054_),
    .A2(_13089_),
    .B1(_13079_),
    .Y(_13090_));
 sky130_fd_sc_hd__a21oi_2 _23031_ (.A1(_13087_),
    .A2(_13088_),
    .B1(_13090_),
    .Y(_13091_));
 sky130_fd_sc_hd__nand2_2 _23032_ (.A(_13086_),
    .B(_13091_),
    .Y(_13092_));
 sky130_fd_sc_hd__nand2_1 _23033_ (.A(_13066_),
    .B(_12508_),
    .Y(_13093_));
 sky130_fd_sc_hd__xor2_2 _23034_ (.A(_12536_),
    .B(_13093_),
    .X(_13095_));
 sky130_fd_sc_hd__nand3_2 _23035_ (.A(_13074_),
    .B(_12872_),
    .C(_13069_),
    .Y(_13096_));
 sky130_fd_sc_hd__xnor2_4 _23036_ (.A(_13095_),
    .B(_13096_),
    .Y(_13097_));
 sky130_fd_sc_hd__nand2_4 _23037_ (.A(_13092_),
    .B(_13097_),
    .Y(_13098_));
 sky130_fd_sc_hd__clkinvlp_2 _23038_ (.A(_13097_),
    .Y(_13099_));
 sky130_fd_sc_hd__nand3_4 _23039_ (.A(_13086_),
    .B(_13091_),
    .C(_13099_),
    .Y(_13100_));
 sky130_fd_sc_hd__nand2_8 _23040_ (.A(_13100_),
    .B(_13098_),
    .Y(_13101_));
 sky130_fd_sc_hd__buf_8 _23041_ (.A(_13101_),
    .X(_13102_));
 sky130_fd_sc_hd__buf_6 _23042_ (.A(net236),
    .X(\div1i.quot[6] ));
 sky130_fd_sc_hd__nand2_1 _23043_ (.A(_12686_),
    .B(_12774_),
    .Y(_13103_));
 sky130_fd_sc_hd__inv_2 _23044_ (.A(_12779_),
    .Y(_13105_));
 sky130_fd_sc_hd__nand2_1 _23045_ (.A(_13103_),
    .B(_13105_),
    .Y(_13106_));
 sky130_fd_sc_hd__inv_2 _23046_ (.A(_12753_),
    .Y(_13107_));
 sky130_fd_sc_hd__nand2_2 _23047_ (.A(_13106_),
    .B(_13107_),
    .Y(_13108_));
 sky130_fd_sc_hd__nand2_1 _23048_ (.A(_13108_),
    .B(_12752_),
    .Y(_13109_));
 sky130_fd_sc_hd__inv_2 _23049_ (.A(_12741_),
    .Y(_13110_));
 sky130_fd_sc_hd__nand2_1 _23050_ (.A(_13109_),
    .B(_13110_),
    .Y(_13111_));
 sky130_fd_sc_hd__nand3_1 _23051_ (.A(_13108_),
    .B(_12741_),
    .C(_12752_),
    .Y(_13112_));
 sky130_fd_sc_hd__nand2_1 _23052_ (.A(_13111_),
    .B(_13112_),
    .Y(_13113_));
 sky130_fd_sc_hd__nand2_1 _23053_ (.A(_13113_),
    .B(_11983_),
    .Y(_13114_));
 sky130_fd_sc_hd__nand3_1 _23054_ (.A(_13103_),
    .B(_12753_),
    .C(_13105_),
    .Y(_13116_));
 sky130_fd_sc_hd__nand3_2 _23055_ (.A(_13108_),
    .B(_11986_),
    .C(_13116_),
    .Y(_13117_));
 sky130_fd_sc_hd__inv_2 _23056_ (.A(_13117_),
    .Y(_13118_));
 sky130_fd_sc_hd__nand3_2 _23057_ (.A(_13111_),
    .B(_11990_),
    .C(_13112_),
    .Y(_13119_));
 sky130_fd_sc_hd__nand3_1 _23058_ (.A(_13114_),
    .B(_13118_),
    .C(_13119_),
    .Y(_13120_));
 sky130_fd_sc_hd__nand2_1 _23059_ (.A(_13120_),
    .B(_13119_),
    .Y(_13121_));
 sky130_fd_sc_hd__inv_2 _23060_ (.A(_12773_),
    .Y(_13122_));
 sky130_fd_sc_hd__nand2_1 _23061_ (.A(_12686_),
    .B(_13122_),
    .Y(_13123_));
 sky130_fd_sc_hd__nand2_1 _23062_ (.A(_13123_),
    .B(_12770_),
    .Y(_13124_));
 sky130_fd_sc_hd__inv_2 _23063_ (.A(_12762_),
    .Y(_13125_));
 sky130_fd_sc_hd__nand2_1 _23064_ (.A(_13124_),
    .B(_13125_),
    .Y(_13127_));
 sky130_fd_sc_hd__nand3_1 _23065_ (.A(_13123_),
    .B(_12762_),
    .C(_12770_),
    .Y(_13128_));
 sky130_fd_sc_hd__nand2_1 _23066_ (.A(_13127_),
    .B(_13128_),
    .Y(_13129_));
 sky130_fd_sc_hd__nand2_1 _23067_ (.A(_13129_),
    .B(_12002_),
    .Y(_13130_));
 sky130_fd_sc_hd__or2_1 _23068_ (.A(_13122_),
    .B(_12686_),
    .X(_13131_));
 sky130_fd_sc_hd__nand2_1 _23069_ (.A(_13131_),
    .B(_13123_),
    .Y(_13132_));
 sky130_fd_sc_hd__inv_2 _23070_ (.A(_13132_),
    .Y(_13133_));
 sky130_fd_sc_hd__nand2_1 _23071_ (.A(_13133_),
    .B(_12008_),
    .Y(_13134_));
 sky130_fd_sc_hd__inv_2 _23072_ (.A(_13134_),
    .Y(_13135_));
 sky130_fd_sc_hd__inv_2 _23073_ (.A(_13129_),
    .Y(_13136_));
 sky130_fd_sc_hd__nand2_1 _23074_ (.A(_13136_),
    .B(_12012_),
    .Y(_13138_));
 sky130_fd_sc_hd__inv_2 _23075_ (.A(_13138_),
    .Y(_13139_));
 sky130_fd_sc_hd__a21oi_1 _23076_ (.A1(_13130_),
    .A2(_13135_),
    .B1(_13139_),
    .Y(_13140_));
 sky130_fd_sc_hd__nand2_1 _23077_ (.A(_13108_),
    .B(_13116_),
    .Y(_13141_));
 sky130_fd_sc_hd__nand2_1 _23078_ (.A(_13141_),
    .B(_12017_),
    .Y(_13142_));
 sky130_fd_sc_hd__nand2_1 _23079_ (.A(_13142_),
    .B(_13117_),
    .Y(_13143_));
 sky130_fd_sc_hd__inv_2 _23080_ (.A(_13143_),
    .Y(_13144_));
 sky130_fd_sc_hd__nand3_1 _23081_ (.A(_13114_),
    .B(_13144_),
    .C(_13119_),
    .Y(_13145_));
 sky130_fd_sc_hd__nor2_1 _23082_ (.A(_13140_),
    .B(_13145_),
    .Y(_13146_));
 sky130_fd_sc_hd__nor2_1 _23083_ (.A(_13121_),
    .B(_13146_),
    .Y(_13147_));
 sky130_fd_sc_hd__inv_2 _23084_ (.A(_13145_),
    .Y(_13149_));
 sky130_fd_sc_hd__nand2_1 _23085_ (.A(_12579_),
    .B(_12582_),
    .Y(_13150_));
 sky130_fd_sc_hd__nand2_1 _23086_ (.A(_13150_),
    .B(_12583_),
    .Y(_13151_));
 sky130_fd_sc_hd__nand2_1 _23087_ (.A(_13151_),
    .B(_12585_),
    .Y(_13152_));
 sky130_fd_sc_hd__nand2_1 _23088_ (.A(_13152_),
    .B(_12030_),
    .Y(_13153_));
 sky130_fd_sc_hd__o21ai_1 _23089_ (.A1(_12032_),
    .A2(\div1i.quot[7] ),
    .B1(_12033_),
    .Y(_13154_));
 sky130_fd_sc_hd__nand3_1 _23090_ (.A(_13151_),
    .B(_12035_),
    .C(_12585_),
    .Y(_13155_));
 sky130_fd_sc_hd__inv_2 _23091_ (.A(_13155_),
    .Y(_13156_));
 sky130_fd_sc_hd__a21o_1 _23092_ (.A1(_13153_),
    .A2(_13154_),
    .B1(_13156_),
    .X(_13157_));
 sky130_fd_sc_hd__nand2_1 _23093_ (.A(_12586_),
    .B(_12570_),
    .Y(_13158_));
 sky130_fd_sc_hd__nand2_1 _23094_ (.A(_12585_),
    .B(_12579_),
    .Y(_13160_));
 sky130_fd_sc_hd__xor2_1 _23095_ (.A(_13158_),
    .B(_13160_),
    .X(_13161_));
 sky130_fd_sc_hd__nand2_1 _23096_ (.A(_13161_),
    .B(_12043_),
    .Y(_13162_));
 sky130_fd_sc_hd__nand2_1 _23097_ (.A(_13157_),
    .B(_13162_),
    .Y(_13163_));
 sky130_fd_sc_hd__inv_2 _23098_ (.A(_13161_),
    .Y(_13164_));
 sky130_fd_sc_hd__nand2_1 _23099_ (.A(_13164_),
    .B(_12047_),
    .Y(_13165_));
 sky130_fd_sc_hd__nand2_1 _23100_ (.A(_13163_),
    .B(_13165_),
    .Y(_13166_));
 sky130_fd_sc_hd__nand2_1 _23101_ (.A(_12581_),
    .B(_12585_),
    .Y(_13167_));
 sky130_fd_sc_hd__nand2_1 _23102_ (.A(_13167_),
    .B(_12586_),
    .Y(_13168_));
 sky130_fd_sc_hd__nand2_1 _23103_ (.A(_13168_),
    .B(_12674_),
    .Y(_13169_));
 sky130_fd_sc_hd__nand3_1 _23104_ (.A(_13167_),
    .B(_12586_),
    .C(_12675_),
    .Y(_13171_));
 sky130_fd_sc_hd__nand2_1 _23105_ (.A(_13169_),
    .B(_13171_),
    .Y(_13172_));
 sky130_fd_sc_hd__nand2_1 _23106_ (.A(_13172_),
    .B(_12056_),
    .Y(_13173_));
 sky130_fd_sc_hd__nand3_1 _23107_ (.A(_13169_),
    .B(_12058_),
    .C(_13171_),
    .Y(_13174_));
 sky130_fd_sc_hd__nand2_1 _23108_ (.A(_13173_),
    .B(_13174_),
    .Y(_13175_));
 sky130_fd_sc_hd__inv_2 _23109_ (.A(_13175_),
    .Y(_13176_));
 sky130_fd_sc_hd__nand2_1 _23110_ (.A(_13166_),
    .B(_13176_),
    .Y(_13177_));
 sky130_fd_sc_hd__nand2_1 _23111_ (.A(_13177_),
    .B(_13174_),
    .Y(_13178_));
 sky130_fd_sc_hd__nand2_1 _23112_ (.A(_13171_),
    .B(_12672_),
    .Y(_13179_));
 sky130_fd_sc_hd__xor2_2 _23113_ (.A(_12664_),
    .B(_13179_),
    .X(_13180_));
 sky130_fd_sc_hd__buf_6 _23114_ (.A(_09823_),
    .X(_13182_));
 sky130_fd_sc_hd__nand2_1 _23115_ (.A(_13180_),
    .B(_13182_),
    .Y(_13183_));
 sky130_fd_sc_hd__nand2_1 _23116_ (.A(_13178_),
    .B(_13183_),
    .Y(_13184_));
 sky130_fd_sc_hd__or2_1 _23117_ (.A(_09823_),
    .B(_13180_),
    .X(_13185_));
 sky130_fd_sc_hd__nand2_1 _23118_ (.A(_13184_),
    .B(_13185_),
    .Y(_13186_));
 sky130_fd_sc_hd__nor2_1 _23119_ (.A(_12664_),
    .B(_12674_),
    .Y(_13187_));
 sky130_fd_sc_hd__nand3_1 _23120_ (.A(_13167_),
    .B(_13187_),
    .C(_12586_),
    .Y(_13188_));
 sky130_fd_sc_hd__inv_2 _23121_ (.A(_12681_),
    .Y(_13189_));
 sky130_fd_sc_hd__nand2_1 _23122_ (.A(_13188_),
    .B(_13189_),
    .Y(_13190_));
 sky130_fd_sc_hd__nand2_1 _23123_ (.A(_13190_),
    .B(_12652_),
    .Y(_13191_));
 sky130_fd_sc_hd__nand2_1 _23124_ (.A(_13191_),
    .B(_12649_),
    .Y(_13193_));
 sky130_fd_sc_hd__nand2_1 _23125_ (.A(_13193_),
    .B(_12642_),
    .Y(_13194_));
 sky130_fd_sc_hd__nand3_1 _23126_ (.A(_13191_),
    .B(_12641_),
    .C(_12649_),
    .Y(_13195_));
 sky130_fd_sc_hd__nand2_1 _23127_ (.A(_13194_),
    .B(_13195_),
    .Y(_13196_));
 sky130_fd_sc_hd__buf_6 _23128_ (.A(_08738_),
    .X(_13197_));
 sky130_fd_sc_hd__nand2_1 _23129_ (.A(_13196_),
    .B(_13197_),
    .Y(_13198_));
 sky130_fd_sc_hd__nand3_1 _23130_ (.A(_13188_),
    .B(_12651_),
    .C(_13189_),
    .Y(_13199_));
 sky130_fd_sc_hd__nand2_1 _23131_ (.A(_13191_),
    .B(_13199_),
    .Y(_13200_));
 sky130_fd_sc_hd__nand2_1 _23132_ (.A(_13200_),
    .B(_12085_),
    .Y(_13201_));
 sky130_fd_sc_hd__nand3_2 _23133_ (.A(_13191_),
    .B(_12087_),
    .C(_13199_),
    .Y(_13202_));
 sky130_fd_sc_hd__nand2_1 _23134_ (.A(_13201_),
    .B(_13202_),
    .Y(_13204_));
 sky130_fd_sc_hd__inv_2 _23135_ (.A(_13204_),
    .Y(_13205_));
 sky130_fd_sc_hd__nand3_1 _23136_ (.A(_13194_),
    .B(_10939_),
    .C(_13195_),
    .Y(_13206_));
 sky130_fd_sc_hd__nand3_1 _23137_ (.A(_13198_),
    .B(_13205_),
    .C(_13206_),
    .Y(_13207_));
 sky130_fd_sc_hd__inv_2 _23138_ (.A(_13207_),
    .Y(_13208_));
 sky130_fd_sc_hd__nand2_1 _23139_ (.A(_13186_),
    .B(_13208_),
    .Y(_13209_));
 sky130_fd_sc_hd__inv_2 _23140_ (.A(_13202_),
    .Y(_13210_));
 sky130_fd_sc_hd__a21boi_1 _23141_ (.A1(_13198_),
    .A2(_13210_),
    .B1_N(_13206_),
    .Y(_13211_));
 sky130_fd_sc_hd__nand2_1 _23142_ (.A(_13209_),
    .B(_13211_),
    .Y(_13212_));
 sky130_fd_sc_hd__nand2_1 _23143_ (.A(_13138_),
    .B(_13130_),
    .Y(_13213_));
 sky130_fd_sc_hd__inv_2 _23144_ (.A(_13213_),
    .Y(_13215_));
 sky130_fd_sc_hd__nand2_1 _23145_ (.A(_13132_),
    .B(_12101_),
    .Y(_13216_));
 sky130_fd_sc_hd__nand2_1 _23146_ (.A(_13134_),
    .B(_13216_),
    .Y(_13217_));
 sky130_fd_sc_hd__inv_4 _23147_ (.A(_13217_),
    .Y(_13218_));
 sky130_fd_sc_hd__nand2_1 _23148_ (.A(_13215_),
    .B(_13218_),
    .Y(_13219_));
 sky130_fd_sc_hd__inv_2 _23149_ (.A(_13219_),
    .Y(_13220_));
 sky130_fd_sc_hd__nand3_1 _23150_ (.A(_13149_),
    .B(_13212_),
    .C(_13220_),
    .Y(_13221_));
 sky130_fd_sc_hd__nand2_2 _23151_ (.A(_13147_),
    .B(_13221_),
    .Y(_13222_));
 sky130_fd_sc_hd__inv_2 _23152_ (.A(_12869_),
    .Y(_13223_));
 sky130_fd_sc_hd__inv_2 _23153_ (.A(_12879_),
    .Y(_13224_));
 sky130_fd_sc_hd__nand2_1 _23154_ (.A(_12782_),
    .B(_13224_),
    .Y(_13226_));
 sky130_fd_sc_hd__nand2_1 _23155_ (.A(_13226_),
    .B(_12878_),
    .Y(_13227_));
 sky130_fd_sc_hd__or2_1 _23156_ (.A(_13223_),
    .B(_13227_),
    .X(_13228_));
 sky130_fd_sc_hd__nand2_1 _23157_ (.A(_13227_),
    .B(_13223_),
    .Y(_13229_));
 sky130_fd_sc_hd__nand2_1 _23158_ (.A(_13228_),
    .B(_13229_),
    .Y(_13230_));
 sky130_fd_sc_hd__nand2_1 _23159_ (.A(_13230_),
    .B(_12118_),
    .Y(_13231_));
 sky130_fd_sc_hd__nand3_1 _23160_ (.A(_13228_),
    .B(_12120_),
    .C(_13229_),
    .Y(_13232_));
 sky130_fd_sc_hd__nand2_1 _23161_ (.A(_13231_),
    .B(_13232_),
    .Y(_13233_));
 sky130_fd_sc_hd__inv_2 _23162_ (.A(_13233_),
    .Y(_13234_));
 sky130_fd_sc_hd__or2_1 _23163_ (.A(_13224_),
    .B(_12782_),
    .X(_13235_));
 sky130_fd_sc_hd__nand2_1 _23164_ (.A(_13235_),
    .B(_13226_),
    .Y(_13237_));
 sky130_fd_sc_hd__inv_2 _23165_ (.A(_13237_),
    .Y(_13238_));
 sky130_fd_sc_hd__nand2_1 _23166_ (.A(_13238_),
    .B(_11671_),
    .Y(_13239_));
 sky130_fd_sc_hd__nand2_1 _23167_ (.A(_13237_),
    .B(_12817_),
    .Y(_13240_));
 sky130_fd_sc_hd__nand2_1 _23168_ (.A(_13239_),
    .B(_13240_),
    .Y(_13241_));
 sky130_fd_sc_hd__inv_2 _23169_ (.A(_13241_),
    .Y(_13242_));
 sky130_fd_sc_hd__nand2_1 _23170_ (.A(_13234_),
    .B(_13242_),
    .Y(_13243_));
 sky130_fd_sc_hd__inv_2 _23171_ (.A(_13243_),
    .Y(_13244_));
 sky130_fd_sc_hd__nand2_1 _23172_ (.A(_13222_),
    .B(_13244_),
    .Y(_13245_));
 sky130_fd_sc_hd__inv_2 _23173_ (.A(_13239_),
    .Y(_13246_));
 sky130_fd_sc_hd__a21boi_2 _23174_ (.A1(_13231_),
    .A2(_13246_),
    .B1_N(_13232_),
    .Y(_13248_));
 sky130_fd_sc_hd__nand2_1 _23175_ (.A(_13245_),
    .B(_13248_),
    .Y(_13249_));
 sky130_fd_sc_hd__nand2_1 _23176_ (.A(_12782_),
    .B(_12880_),
    .Y(_13250_));
 sky130_fd_sc_hd__inv_2 _23177_ (.A(_12884_),
    .Y(_13251_));
 sky130_fd_sc_hd__nand2_1 _23178_ (.A(_13250_),
    .B(_13251_),
    .Y(_13252_));
 sky130_fd_sc_hd__inv_2 _23179_ (.A(_12860_),
    .Y(_13253_));
 sky130_fd_sc_hd__nand2_1 _23180_ (.A(_13252_),
    .B(_13253_),
    .Y(_13254_));
 sky130_fd_sc_hd__nand3_1 _23181_ (.A(_13250_),
    .B(_12860_),
    .C(_13251_),
    .Y(_13255_));
 sky130_fd_sc_hd__nand2_1 _23182_ (.A(_13254_),
    .B(_13255_),
    .Y(_13256_));
 sky130_fd_sc_hd__inv_2 _23183_ (.A(_13256_),
    .Y(_13257_));
 sky130_fd_sc_hd__nand2_1 _23184_ (.A(_13257_),
    .B(_12147_),
    .Y(_13259_));
 sky130_fd_sc_hd__nand2_1 _23185_ (.A(_13256_),
    .B(_12149_),
    .Y(_13260_));
 sky130_fd_sc_hd__nand2_1 _23186_ (.A(_13259_),
    .B(_13260_),
    .Y(_13261_));
 sky130_fd_sc_hd__inv_2 _23187_ (.A(_13261_),
    .Y(_13262_));
 sky130_fd_sc_hd__nand2_1 _23188_ (.A(_13249_),
    .B(_13262_),
    .Y(_13263_));
 sky130_fd_sc_hd__inv_6 _23189_ (.A(_13101_),
    .Y(_13264_));
 sky130_fd_sc_hd__nand3_1 _23190_ (.A(_13245_),
    .B(_13261_),
    .C(_13248_),
    .Y(_13265_));
 sky130_fd_sc_hd__nand3_1 _23191_ (.A(_13263_),
    .B(_13264_),
    .C(_13265_),
    .Y(_13266_));
 sky130_fd_sc_hd__nand2_1 _23192_ (.A(net236),
    .B(_13257_),
    .Y(_13267_));
 sky130_fd_sc_hd__nand2_1 _23193_ (.A(_13266_),
    .B(_13267_),
    .Y(_13268_));
 sky130_fd_sc_hd__nand2_1 _23194_ (.A(_13268_),
    .B(_11701_),
    .Y(_13270_));
 sky130_fd_sc_hd__nand3_1 _23195_ (.A(_13266_),
    .B(_11703_),
    .C(_13267_),
    .Y(_13271_));
 sky130_fd_sc_hd__nand2_1 _23196_ (.A(_13270_),
    .B(_13271_),
    .Y(_13272_));
 sky130_fd_sc_hd__nand2_1 _23197_ (.A(_13222_),
    .B(_13242_),
    .Y(_13273_));
 sky130_fd_sc_hd__nand2_1 _23198_ (.A(_13273_),
    .B(_13239_),
    .Y(_13274_));
 sky130_fd_sc_hd__nand2_1 _23199_ (.A(_13274_),
    .B(_13234_),
    .Y(_13275_));
 sky130_fd_sc_hd__nand3_1 _23200_ (.A(_13273_),
    .B(_13233_),
    .C(_13239_),
    .Y(_13276_));
 sky130_fd_sc_hd__nand2_1 _23201_ (.A(_13275_),
    .B(_13276_),
    .Y(_13277_));
 sky130_fd_sc_hd__nand2_1 _23202_ (.A(_13277_),
    .B(_13264_),
    .Y(_13278_));
 sky130_fd_sc_hd__nand2_1 _23203_ (.A(net236),
    .B(_13230_),
    .Y(_13279_));
 sky130_fd_sc_hd__nand2_1 _23204_ (.A(_13278_),
    .B(_13279_),
    .Y(_13281_));
 sky130_fd_sc_hd__nand2_1 _23205_ (.A(_13281_),
    .B(_11715_),
    .Y(_13282_));
 sky130_fd_sc_hd__nand3_2 _23206_ (.A(_13278_),
    .B(_11717_),
    .C(_13279_),
    .Y(_13283_));
 sky130_fd_sc_hd__nand2_1 _23207_ (.A(_13282_),
    .B(_13283_),
    .Y(_13284_));
 sky130_fd_sc_hd__nor2_1 _23208_ (.A(_13272_),
    .B(_13284_),
    .Y(_13285_));
 sky130_fd_sc_hd__nand2_1 _23209_ (.A(_13220_),
    .B(_13212_),
    .Y(_13286_));
 sky130_fd_sc_hd__nand2_1 _23210_ (.A(_13286_),
    .B(_13140_),
    .Y(_13287_));
 sky130_fd_sc_hd__nand2_1 _23211_ (.A(_13287_),
    .B(_13144_),
    .Y(_13288_));
 sky130_fd_sc_hd__nand2_1 _23212_ (.A(_13288_),
    .B(_13117_),
    .Y(_13289_));
 sky130_fd_sc_hd__nand3_1 _23213_ (.A(_13289_),
    .B(_13119_),
    .C(_13114_),
    .Y(_13290_));
 sky130_fd_sc_hd__nand2_1 _23214_ (.A(_13114_),
    .B(_13119_),
    .Y(_13292_));
 sky130_fd_sc_hd__nand3_1 _23215_ (.A(_13288_),
    .B(_13117_),
    .C(_13292_),
    .Y(_13293_));
 sky130_fd_sc_hd__nand2_1 _23216_ (.A(_13290_),
    .B(_13293_),
    .Y(_13294_));
 sky130_fd_sc_hd__nand2_1 _23217_ (.A(_13294_),
    .B(_13264_),
    .Y(_13295_));
 sky130_fd_sc_hd__nand2_1 _23218_ (.A(net236),
    .B(_13113_),
    .Y(_13296_));
 sky130_fd_sc_hd__nand3_1 _23219_ (.A(_13295_),
    .B(_12187_),
    .C(_13296_),
    .Y(_13297_));
 sky130_fd_sc_hd__or2_1 _23220_ (.A(_13242_),
    .B(_13222_),
    .X(_13298_));
 sky130_fd_sc_hd__nand3_1 _23221_ (.A(_13298_),
    .B(_13264_),
    .C(_13273_),
    .Y(_13299_));
 sky130_fd_sc_hd__nand2_1 _23222_ (.A(net236),
    .B(_13238_),
    .Y(_13300_));
 sky130_fd_sc_hd__nand3_1 _23223_ (.A(_13299_),
    .B(_09944_),
    .C(_13300_),
    .Y(_13301_));
 sky130_fd_sc_hd__inv_2 _23224_ (.A(_13301_),
    .Y(_13303_));
 sky130_fd_sc_hd__buf_6 _23225_ (.A(_09944_),
    .X(_13304_));
 sky130_fd_sc_hd__a21o_1 _23226_ (.A1(_13299_),
    .A2(_13300_),
    .B1(_13304_),
    .X(_13305_));
 sky130_fd_sc_hd__o21ai_1 _23227_ (.A1(_13297_),
    .A2(_13303_),
    .B1(_13305_),
    .Y(_13306_));
 sky130_fd_sc_hd__inv_2 _23228_ (.A(_13271_),
    .Y(_13307_));
 sky130_fd_sc_hd__o21ai_1 _23229_ (.A1(_13283_),
    .A2(_13307_),
    .B1(_13270_),
    .Y(_13308_));
 sky130_fd_sc_hd__a21oi_1 _23230_ (.A1(_13285_),
    .A2(_13306_),
    .B1(_13308_),
    .Y(_13309_));
 sky130_fd_sc_hd__inv_2 _23231_ (.A(_13152_),
    .Y(_13310_));
 sky130_fd_sc_hd__nand2_1 _23232_ (.A(_13101_),
    .B(_13310_),
    .Y(_13311_));
 sky130_fd_sc_hd__nand2_1 _23233_ (.A(_13153_),
    .B(_13155_),
    .Y(_13312_));
 sky130_fd_sc_hd__xor2_1 _23234_ (.A(_13154_),
    .B(_13312_),
    .X(_13314_));
 sky130_fd_sc_hd__nand3b_1 _23235_ (.A_N(_13314_),
    .B(_13098_),
    .C(_13100_),
    .Y(_13315_));
 sky130_fd_sc_hd__nand2_1 _23236_ (.A(_13311_),
    .B(_13315_),
    .Y(_13316_));
 sky130_fd_sc_hd__nand2_1 _23237_ (.A(_13316_),
    .B(_11069_),
    .Y(_13317_));
 sky130_fd_sc_hd__nor2_1 _23238_ (.A(_12032_),
    .B(_12872_),
    .Y(_13318_));
 sky130_fd_sc_hd__or2_1 _23239_ (.A(_11412_),
    .B(_13318_),
    .X(_13319_));
 sky130_fd_sc_hd__nand2_1 _23240_ (.A(_13319_),
    .B(_12583_),
    .Y(_13320_));
 sky130_fd_sc_hd__inv_2 _23241_ (.A(_13320_),
    .Y(_13321_));
 sky130_fd_sc_hd__nand2_1 _23242_ (.A(_13101_),
    .B(_13321_),
    .Y(_13322_));
 sky130_fd_sc_hd__nand3_1 _23243_ (.A(_13098_),
    .B(_13100_),
    .C(_13318_),
    .Y(_13323_));
 sky130_fd_sc_hd__nand2_1 _23244_ (.A(_13322_),
    .B(_13323_),
    .Y(_13325_));
 sky130_fd_sc_hd__nand2_2 _23245_ (.A(_13325_),
    .B(_11421_),
    .Y(_13326_));
 sky130_fd_sc_hd__nand2_1 _23246_ (.A(_13317_),
    .B(_13326_),
    .Y(_13327_));
 sky130_fd_sc_hd__inv_2 _23247_ (.A(_13327_),
    .Y(_13328_));
 sky130_fd_sc_hd__nand3_1 _23248_ (.A(_13322_),
    .B(_11426_),
    .C(_13323_),
    .Y(_13329_));
 sky130_fd_sc_hd__nand3_2 _23249_ (.A(_13101_),
    .B(_12033_),
    .C(_12221_),
    .Y(_13330_));
 sky130_fd_sc_hd__inv_2 _23250_ (.A(_13330_),
    .Y(_13331_));
 sky130_fd_sc_hd__nand3_2 _23251_ (.A(_13326_),
    .B(_13329_),
    .C(_13331_),
    .Y(_13332_));
 sky130_fd_sc_hd__nand2_1 _23252_ (.A(_13328_),
    .B(_13332_),
    .Y(_13333_));
 sky130_fd_sc_hd__or2_1 _23253_ (.A(_11069_),
    .B(_13316_),
    .X(_13334_));
 sky130_fd_sc_hd__nand2_1 _23254_ (.A(_13333_),
    .B(_13334_),
    .Y(_13336_));
 sky130_fd_sc_hd__inv_2 _23255_ (.A(_13336_),
    .Y(_13337_));
 sky130_fd_sc_hd__clkinvlp_2 _23256_ (.A(_13200_),
    .Y(_13338_));
 sky130_fd_sc_hd__nand2_1 _23257_ (.A(_13102_),
    .B(_13338_),
    .Y(_13339_));
 sky130_fd_sc_hd__nand2_1 _23258_ (.A(_13186_),
    .B(_13205_),
    .Y(_13340_));
 sky130_fd_sc_hd__nand3_1 _23259_ (.A(_13184_),
    .B(_13204_),
    .C(_13185_),
    .Y(_13341_));
 sky130_fd_sc_hd__nand2_1 _23260_ (.A(_13340_),
    .B(_13341_),
    .Y(_13342_));
 sky130_fd_sc_hd__inv_2 _23261_ (.A(_13342_),
    .Y(_13343_));
 sky130_fd_sc_hd__nand3_1 _23262_ (.A(_13098_),
    .B(_13100_),
    .C(_13343_),
    .Y(_13344_));
 sky130_fd_sc_hd__nand2_1 _23263_ (.A(_13339_),
    .B(_13344_),
    .Y(_13345_));
 sky130_fd_sc_hd__nand2_1 _23264_ (.A(_13345_),
    .B(_11482_),
    .Y(_13347_));
 sky130_fd_sc_hd__nand3_1 _23265_ (.A(_13339_),
    .B(_11484_),
    .C(_13344_),
    .Y(_13348_));
 sky130_fd_sc_hd__nand2_1 _23266_ (.A(_13347_),
    .B(_13348_),
    .Y(_13349_));
 sky130_fd_sc_hd__inv_2 _23267_ (.A(_13349_),
    .Y(_13350_));
 sky130_fd_sc_hd__nand2_1 _23268_ (.A(_13102_),
    .B(_13180_),
    .Y(_13351_));
 sky130_fd_sc_hd__nand2_1 _23269_ (.A(_13185_),
    .B(_13183_),
    .Y(_13352_));
 sky130_fd_sc_hd__xor2_1 _23270_ (.A(_13178_),
    .B(_13352_),
    .X(_13353_));
 sky130_fd_sc_hd__nand3_1 _23271_ (.A(_13098_),
    .B(_13100_),
    .C(_13353_),
    .Y(_13354_));
 sky130_fd_sc_hd__nand2_1 _23272_ (.A(_13351_),
    .B(_13354_),
    .Y(_13355_));
 sky130_fd_sc_hd__nand2_1 _23273_ (.A(_13355_),
    .B(_11496_),
    .Y(_13356_));
 sky130_fd_sc_hd__nand3_2 _23274_ (.A(_13351_),
    .B(_11494_),
    .C(_13354_),
    .Y(_13358_));
 sky130_fd_sc_hd__nand2_1 _23275_ (.A(_13358_),
    .B(_13356_),
    .Y(_13359_));
 sky130_fd_sc_hd__inv_2 _23276_ (.A(_13359_),
    .Y(_13360_));
 sky130_fd_sc_hd__nand2_1 _23277_ (.A(_13350_),
    .B(_13360_),
    .Y(_13361_));
 sky130_fd_sc_hd__inv_2 _23278_ (.A(_13172_),
    .Y(_13362_));
 sky130_fd_sc_hd__nand2_1 _23279_ (.A(_13102_),
    .B(_13362_),
    .Y(_13363_));
 sky130_fd_sc_hd__or2_1 _23280_ (.A(_13176_),
    .B(_13166_),
    .X(_13364_));
 sky130_fd_sc_hd__nand2_1 _23281_ (.A(_13364_),
    .B(_13177_),
    .Y(_13365_));
 sky130_fd_sc_hd__inv_2 _23282_ (.A(_13365_),
    .Y(_13366_));
 sky130_fd_sc_hd__nand3_1 _23283_ (.A(_13098_),
    .B(_13100_),
    .C(_13366_),
    .Y(_13367_));
 sky130_fd_sc_hd__nand2_1 _23284_ (.A(_13363_),
    .B(_13367_),
    .Y(_13369_));
 sky130_fd_sc_hd__nand2_2 _23285_ (.A(_13369_),
    .B(_11105_),
    .Y(_13370_));
 sky130_fd_sc_hd__nand3_2 _23286_ (.A(_13363_),
    .B(_12261_),
    .C(_13367_),
    .Y(_13371_));
 sky130_fd_sc_hd__nand2_4 _23287_ (.A(_13371_),
    .B(_13370_),
    .Y(_13372_));
 sky130_fd_sc_hd__inv_2 _23288_ (.A(_13372_),
    .Y(_13373_));
 sky130_fd_sc_hd__nand2_1 _23289_ (.A(_13101_),
    .B(_13164_),
    .Y(_13374_));
 sky130_fd_sc_hd__nand2_1 _23290_ (.A(_13165_),
    .B(_13162_),
    .Y(_13375_));
 sky130_fd_sc_hd__xnor2_1 _23291_ (.A(_13157_),
    .B(_13375_),
    .Y(_13376_));
 sky130_fd_sc_hd__nand3_1 _23292_ (.A(_13098_),
    .B(_13100_),
    .C(_13376_),
    .Y(_13377_));
 sky130_fd_sc_hd__nand2_1 _23293_ (.A(_13374_),
    .B(_13377_),
    .Y(_13378_));
 sky130_fd_sc_hd__nand2_1 _23294_ (.A(_13378_),
    .B(_12270_),
    .Y(_13380_));
 sky130_fd_sc_hd__nand3_1 _23295_ (.A(_13374_),
    .B(_11117_),
    .C(_13377_),
    .Y(_13381_));
 sky130_fd_sc_hd__nand2_1 _23296_ (.A(_13380_),
    .B(_13381_),
    .Y(_13382_));
 sky130_fd_sc_hd__inv_4 _23297_ (.A(_13382_),
    .Y(_13383_));
 sky130_fd_sc_hd__nand2_1 _23298_ (.A(_13373_),
    .B(_13383_),
    .Y(_13384_));
 sky130_fd_sc_hd__nor2_1 _23299_ (.A(_13361_),
    .B(_13384_),
    .Y(_13385_));
 sky130_fd_sc_hd__nand2_1 _23300_ (.A(_13337_),
    .B(_13385_),
    .Y(_13386_));
 sky130_fd_sc_hd__inv_2 _23301_ (.A(_13371_),
    .Y(_13387_));
 sky130_fd_sc_hd__o21ai_2 _23302_ (.A1(_13380_),
    .A2(_13387_),
    .B1(_13370_),
    .Y(_13388_));
 sky130_fd_sc_hd__nor2_1 _23303_ (.A(_13349_),
    .B(_13359_),
    .Y(_13389_));
 sky130_fd_sc_hd__inv_2 _23304_ (.A(_13348_),
    .Y(_13391_));
 sky130_fd_sc_hd__o21ai_1 _23305_ (.A1(_13358_),
    .A2(_13391_),
    .B1(_13347_),
    .Y(_13392_));
 sky130_fd_sc_hd__a21oi_1 _23306_ (.A1(_13388_),
    .A2(_13389_),
    .B1(_13392_),
    .Y(_13393_));
 sky130_fd_sc_hd__nand2_2 _23307_ (.A(_13386_),
    .B(_13393_),
    .Y(_13394_));
 sky130_fd_sc_hd__nand2_1 _23308_ (.A(_13212_),
    .B(_13218_),
    .Y(_13395_));
 sky130_fd_sc_hd__or2_1 _23309_ (.A(_13218_),
    .B(_13212_),
    .X(_13396_));
 sky130_fd_sc_hd__nand3_1 _23310_ (.A(_13264_),
    .B(_13395_),
    .C(_13396_),
    .Y(_13397_));
 sky130_fd_sc_hd__nand2_1 _23311_ (.A(_13101_),
    .B(_13133_),
    .Y(_13398_));
 sky130_fd_sc_hd__nand2_1 _23312_ (.A(_13397_),
    .B(_13398_),
    .Y(_13399_));
 sky130_fd_sc_hd__nand2_1 _23313_ (.A(_13399_),
    .B(_11614_),
    .Y(_13400_));
 sky130_fd_sc_hd__nand3_1 _23314_ (.A(_13397_),
    .B(_11616_),
    .C(_13398_),
    .Y(_13402_));
 sky130_fd_sc_hd__nand2_1 _23315_ (.A(_13400_),
    .B(_13402_),
    .Y(_13403_));
 sky130_fd_sc_hd__inv_2 _23316_ (.A(_13403_),
    .Y(_13404_));
 sky130_fd_sc_hd__nand2_1 _23317_ (.A(_13198_),
    .B(_13206_),
    .Y(_13405_));
 sky130_fd_sc_hd__nand2_1 _23318_ (.A(_13340_),
    .B(_13202_),
    .Y(_13406_));
 sky130_fd_sc_hd__xor2_1 _23319_ (.A(_13405_),
    .B(_13406_),
    .X(_13407_));
 sky130_fd_sc_hd__nand2_1 _23320_ (.A(_13407_),
    .B(_13264_),
    .Y(_13408_));
 sky130_fd_sc_hd__nand2_1 _23321_ (.A(_13102_),
    .B(_13196_),
    .Y(_13409_));
 sky130_fd_sc_hd__nand2_1 _23322_ (.A(_13408_),
    .B(_13409_),
    .Y(_13410_));
 sky130_fd_sc_hd__nand2_1 _23323_ (.A(_13410_),
    .B(_12771_),
    .Y(_13411_));
 sky130_fd_sc_hd__nand3_2 _23324_ (.A(_13408_),
    .B(_08951_),
    .C(_13409_),
    .Y(_13413_));
 sky130_fd_sc_hd__nand2_1 _23325_ (.A(_13411_),
    .B(_13413_),
    .Y(_13414_));
 sky130_fd_sc_hd__inv_2 _23326_ (.A(_13414_),
    .Y(_13415_));
 sky130_fd_sc_hd__nand2_1 _23327_ (.A(_13404_),
    .B(_13415_),
    .Y(_13416_));
 sky130_fd_sc_hd__nand2_1 _23328_ (.A(_13395_),
    .B(_13134_),
    .Y(_13417_));
 sky130_fd_sc_hd__nand2_1 _23329_ (.A(_13417_),
    .B(_13215_),
    .Y(_13418_));
 sky130_fd_sc_hd__nand3_1 _23330_ (.A(_13395_),
    .B(_13213_),
    .C(_13134_),
    .Y(_13419_));
 sky130_fd_sc_hd__nand2_1 _23331_ (.A(_13418_),
    .B(_13419_),
    .Y(_13420_));
 sky130_fd_sc_hd__nand2_1 _23332_ (.A(_13420_),
    .B(_13264_),
    .Y(_13421_));
 sky130_fd_sc_hd__nand2_1 _23333_ (.A(_13102_),
    .B(_13129_),
    .Y(_13422_));
 sky130_fd_sc_hd__nand2_1 _23334_ (.A(_13421_),
    .B(_13422_),
    .Y(_13424_));
 sky130_fd_sc_hd__nand2_1 _23335_ (.A(_13424_),
    .B(_11600_),
    .Y(_13425_));
 sky130_fd_sc_hd__nand3_2 _23336_ (.A(_13421_),
    .B(_11603_),
    .C(_13422_),
    .Y(_13426_));
 sky130_fd_sc_hd__nand2_1 _23337_ (.A(_13425_),
    .B(_13426_),
    .Y(_13427_));
 sky130_fd_sc_hd__or2_1 _23338_ (.A(_13141_),
    .B(_13264_),
    .X(_13428_));
 sky130_fd_sc_hd__nand3_1 _23339_ (.A(_13286_),
    .B(_13143_),
    .C(_13140_),
    .Y(_13429_));
 sky130_fd_sc_hd__nand3_1 _23340_ (.A(_13288_),
    .B(_13264_),
    .C(_13429_),
    .Y(_13430_));
 sky130_fd_sc_hd__nand2_1 _23341_ (.A(_13428_),
    .B(_13430_),
    .Y(_13431_));
 sky130_fd_sc_hd__nand2_1 _23342_ (.A(_13431_),
    .B(_11586_),
    .Y(_13432_));
 sky130_fd_sc_hd__nand3_2 _23343_ (.A(_13428_),
    .B(_13430_),
    .C(_11588_),
    .Y(_13433_));
 sky130_fd_sc_hd__nand2_2 _23344_ (.A(_13432_),
    .B(_13433_),
    .Y(_13435_));
 sky130_fd_sc_hd__nor2_1 _23345_ (.A(_13427_),
    .B(_13435_),
    .Y(_13436_));
 sky130_fd_sc_hd__nor2b_1 _23346_ (.A(_13416_),
    .B_N(_13436_),
    .Y(_13437_));
 sky130_fd_sc_hd__nand2_1 _23347_ (.A(_13394_),
    .B(_13437_),
    .Y(_13438_));
 sky130_fd_sc_hd__clkinvlp_2 _23348_ (.A(_13402_),
    .Y(_13439_));
 sky130_fd_sc_hd__o21ai_2 _23349_ (.A1(_13413_),
    .A2(_13439_),
    .B1(_13400_),
    .Y(_13440_));
 sky130_fd_sc_hd__inv_2 _23350_ (.A(_13433_),
    .Y(_13441_));
 sky130_fd_sc_hd__o21ai_1 _23351_ (.A1(_13426_),
    .A2(_13441_),
    .B1(_13432_),
    .Y(_13442_));
 sky130_fd_sc_hd__a21oi_1 _23352_ (.A1(_13436_),
    .A2(_13440_),
    .B1(_13442_),
    .Y(_13443_));
 sky130_fd_sc_hd__nand2_2 _23353_ (.A(_13438_),
    .B(_13443_),
    .Y(_13444_));
 sky130_fd_sc_hd__nand2_1 _23354_ (.A(_13295_),
    .B(_13296_),
    .Y(_13446_));
 sky130_fd_sc_hd__nand2_1 _23355_ (.A(_13446_),
    .B(_11185_),
    .Y(_13447_));
 sky130_fd_sc_hd__nand2_1 _23356_ (.A(_13447_),
    .B(_13297_),
    .Y(_13448_));
 sky130_fd_sc_hd__nand2_1 _23357_ (.A(_13305_),
    .B(_13301_),
    .Y(_13449_));
 sky130_fd_sc_hd__nor2_1 _23358_ (.A(_13448_),
    .B(_13449_),
    .Y(_13450_));
 sky130_fd_sc_hd__nand3_1 _23359_ (.A(_13444_),
    .B(_13285_),
    .C(_13450_),
    .Y(_13451_));
 sky130_fd_sc_hd__nand2_2 _23360_ (.A(_13309_),
    .B(_13451_),
    .Y(_13452_));
 sky130_fd_sc_hd__nand2_1 _23361_ (.A(_12977_),
    .B(_12978_),
    .Y(_13453_));
 sky130_fd_sc_hd__inv_4 _23362_ (.A(_13453_),
    .Y(_13454_));
 sky130_fd_sc_hd__or2_1 _23363_ (.A(_13454_),
    .B(_12888_),
    .X(_13455_));
 sky130_fd_sc_hd__nand2_1 _23364_ (.A(_12888_),
    .B(_13454_),
    .Y(_13457_));
 sky130_fd_sc_hd__nand2_1 _23365_ (.A(_13455_),
    .B(_13457_),
    .Y(_13458_));
 sky130_fd_sc_hd__inv_2 _23366_ (.A(_13458_),
    .Y(_13459_));
 sky130_fd_sc_hd__nand2_1 _23367_ (.A(_13459_),
    .B(_11199_),
    .Y(_13460_));
 sky130_fd_sc_hd__buf_6 _23368_ (.A(_08465_),
    .X(_13461_));
 sky130_fd_sc_hd__nand2_1 _23369_ (.A(_13458_),
    .B(_13461_),
    .Y(_13462_));
 sky130_fd_sc_hd__nand2_1 _23370_ (.A(_13460_),
    .B(_13462_),
    .Y(_13463_));
 sky130_fd_sc_hd__inv_2 _23371_ (.A(_13463_),
    .Y(_13464_));
 sky130_fd_sc_hd__nand2_1 _23372_ (.A(_13254_),
    .B(_12859_),
    .Y(_13465_));
 sky130_fd_sc_hd__inv_2 _23373_ (.A(_12848_),
    .Y(_13466_));
 sky130_fd_sc_hd__nand2_1 _23374_ (.A(_13465_),
    .B(_13466_),
    .Y(_13468_));
 sky130_fd_sc_hd__nand3_1 _23375_ (.A(_13254_),
    .B(_12848_),
    .C(_12859_),
    .Y(_13469_));
 sky130_fd_sc_hd__nand2_1 _23376_ (.A(_13468_),
    .B(_13469_),
    .Y(_13470_));
 sky130_fd_sc_hd__nand2_1 _23377_ (.A(_13470_),
    .B(_12894_),
    .Y(_13471_));
 sky130_fd_sc_hd__nand3_1 _23378_ (.A(_13468_),
    .B(_11754_),
    .C(_13469_),
    .Y(_13472_));
 sky130_fd_sc_hd__nand3_1 _23379_ (.A(_13262_),
    .B(_13471_),
    .C(_13472_),
    .Y(_13473_));
 sky130_fd_sc_hd__inv_2 _23380_ (.A(_13473_),
    .Y(_13474_));
 sky130_fd_sc_hd__nand3_1 _23381_ (.A(_13222_),
    .B(_13244_),
    .C(_13474_),
    .Y(_13475_));
 sky130_fd_sc_hd__inv_2 _23382_ (.A(_13471_),
    .Y(_13476_));
 sky130_fd_sc_hd__o21ai_1 _23383_ (.A1(_13259_),
    .A2(_13476_),
    .B1(_13472_),
    .Y(_13477_));
 sky130_fd_sc_hd__nor2_1 _23384_ (.A(_13248_),
    .B(_13473_),
    .Y(_13479_));
 sky130_fd_sc_hd__nor2_1 _23385_ (.A(_13477_),
    .B(_13479_),
    .Y(_13480_));
 sky130_fd_sc_hd__nand2_1 _23386_ (.A(_13475_),
    .B(_13480_),
    .Y(_13481_));
 sky130_fd_sc_hd__or2_1 _23387_ (.A(_13464_),
    .B(_13481_),
    .X(_13482_));
 sky130_fd_sc_hd__buf_6 _23388_ (.A(_13264_),
    .X(_13483_));
 sky130_fd_sc_hd__nand2_1 _23389_ (.A(_13481_),
    .B(_13464_),
    .Y(_13484_));
 sky130_fd_sc_hd__nand3_1 _23390_ (.A(_13482_),
    .B(_13483_),
    .C(_13484_),
    .Y(_13485_));
 sky130_fd_sc_hd__nand2_1 _23391_ (.A(\div1i.quot[6] ),
    .B(_13459_),
    .Y(_13486_));
 sky130_fd_sc_hd__nand2_1 _23392_ (.A(_13485_),
    .B(_13486_),
    .Y(_13487_));
 sky130_fd_sc_hd__xor2_2 _23393_ (.A(_06754_),
    .B(_13487_),
    .X(_13488_));
 sky130_fd_sc_hd__nand2_1 _23394_ (.A(_13471_),
    .B(_13472_),
    .Y(_13490_));
 sky130_fd_sc_hd__nand2_1 _23395_ (.A(_13263_),
    .B(_13259_),
    .Y(_13491_));
 sky130_fd_sc_hd__xor2_1 _23396_ (.A(_13490_),
    .B(_13491_),
    .X(_13492_));
 sky130_fd_sc_hd__nand2_1 _23397_ (.A(_13492_),
    .B(_13483_),
    .Y(_13493_));
 sky130_fd_sc_hd__nand2_1 _23398_ (.A(\div1i.quot[6] ),
    .B(_13470_),
    .Y(_13494_));
 sky130_fd_sc_hd__nand2_1 _23399_ (.A(_13493_),
    .B(_13494_),
    .Y(_13495_));
 sky130_fd_sc_hd__nand2_1 _23400_ (.A(_13495_),
    .B(_11838_),
    .Y(_13496_));
 sky130_fd_sc_hd__nand3_1 _23401_ (.A(_13493_),
    .B(_11840_),
    .C(_13494_),
    .Y(_13497_));
 sky130_fd_sc_hd__nand2_1 _23402_ (.A(_13496_),
    .B(_13497_),
    .Y(_13498_));
 sky130_fd_sc_hd__nor2_1 _23403_ (.A(_13488_),
    .B(_13498_),
    .Y(_13499_));
 sky130_fd_sc_hd__nand2_1 _23404_ (.A(_13452_),
    .B(_13499_),
    .Y(_13501_));
 sky130_fd_sc_hd__buf_6 _23405_ (.A(_10138_),
    .X(_13502_));
 sky130_fd_sc_hd__nand2_1 _23406_ (.A(_13487_),
    .B(_13502_),
    .Y(_13503_));
 sky130_fd_sc_hd__o21a_1 _23407_ (.A1(_13497_),
    .A2(_13488_),
    .B1(_13503_),
    .X(_13504_));
 sky130_fd_sc_hd__nand2_1 _23408_ (.A(_13501_),
    .B(_13504_),
    .Y(_13505_));
 sky130_fd_sc_hd__nand2_1 _23409_ (.A(_12888_),
    .B(_12980_),
    .Y(_13506_));
 sky130_fd_sc_hd__inv_2 _23410_ (.A(_12983_),
    .Y(_13507_));
 sky130_fd_sc_hd__a21o_1 _23411_ (.A1(_13506_),
    .A2(_13507_),
    .B1(_12961_),
    .X(_13508_));
 sky130_fd_sc_hd__nand3_1 _23412_ (.A(_13506_),
    .B(_12961_),
    .C(_13507_),
    .Y(_13509_));
 sky130_fd_sc_hd__nand2_1 _23413_ (.A(_13508_),
    .B(_13509_),
    .Y(_13510_));
 sky130_fd_sc_hd__inv_2 _23414_ (.A(_13510_),
    .Y(_13512_));
 sky130_fd_sc_hd__nand2_1 _23415_ (.A(_13512_),
    .B(_11797_),
    .Y(_13513_));
 sky130_fd_sc_hd__nand2_1 _23416_ (.A(_13510_),
    .B(_12939_),
    .Y(_13514_));
 sky130_fd_sc_hd__nand2_1 _23417_ (.A(_13513_),
    .B(_13514_),
    .Y(_13515_));
 sky130_fd_sc_hd__inv_4 _23418_ (.A(_13515_),
    .Y(_13516_));
 sky130_fd_sc_hd__nand2_1 _23419_ (.A(_13457_),
    .B(_12978_),
    .Y(_13517_));
 sky130_fd_sc_hd__xor2_2 _23420_ (.A(_12970_),
    .B(_13517_),
    .X(_13518_));
 sky130_fd_sc_hd__inv_2 _23421_ (.A(_13518_),
    .Y(_13519_));
 sky130_fd_sc_hd__nand2_1 _23422_ (.A(_13519_),
    .B(_11774_),
    .Y(_13520_));
 sky130_fd_sc_hd__nand2_1 _23423_ (.A(_13518_),
    .B(_12914_),
    .Y(_13521_));
 sky130_fd_sc_hd__nand2_1 _23424_ (.A(_13520_),
    .B(_13521_),
    .Y(_13523_));
 sky130_fd_sc_hd__or2_1 _23425_ (.A(_13463_),
    .B(_13523_),
    .X(_13524_));
 sky130_fd_sc_hd__inv_4 _23426_ (.A(_13524_),
    .Y(_13525_));
 sky130_fd_sc_hd__nand2_1 _23427_ (.A(_13481_),
    .B(_13525_),
    .Y(_13526_));
 sky130_fd_sc_hd__inv_2 _23428_ (.A(_13460_),
    .Y(_13527_));
 sky130_fd_sc_hd__a21boi_1 _23429_ (.A1(_13527_),
    .A2(_13521_),
    .B1_N(_13520_),
    .Y(_13528_));
 sky130_fd_sc_hd__nand2_1 _23430_ (.A(_13526_),
    .B(_13528_),
    .Y(_13529_));
 sky130_fd_sc_hd__or2_1 _23431_ (.A(_13516_),
    .B(_13529_),
    .X(_13530_));
 sky130_fd_sc_hd__nand2_1 _23432_ (.A(_13529_),
    .B(_13516_),
    .Y(_13531_));
 sky130_fd_sc_hd__nand3_1 _23433_ (.A(_13530_),
    .B(_13483_),
    .C(_13531_),
    .Y(_13532_));
 sky130_fd_sc_hd__nand2_1 _23434_ (.A(\div1i.quot[6] ),
    .B(_13512_),
    .Y(_13534_));
 sky130_fd_sc_hd__nand2_1 _23435_ (.A(_13532_),
    .B(_13534_),
    .Y(_13535_));
 sky130_fd_sc_hd__xor2_2 _23436_ (.A(_11811_),
    .B(_13535_),
    .X(_13536_));
 sky130_fd_sc_hd__buf_4 _23437_ (.A(_10173_),
    .X(_13537_));
 sky130_fd_sc_hd__nand2_1 _23438_ (.A(_13484_),
    .B(_13460_),
    .Y(_13538_));
 sky130_fd_sc_hd__xor2_1 _23439_ (.A(_13523_),
    .B(_13538_),
    .X(_13539_));
 sky130_fd_sc_hd__nand2_1 _23440_ (.A(_13539_),
    .B(_13483_),
    .Y(_13540_));
 sky130_fd_sc_hd__nand2_1 _23441_ (.A(\div1i.quot[6] ),
    .B(_13518_),
    .Y(_13541_));
 sky130_fd_sc_hd__nand2_1 _23442_ (.A(_13540_),
    .B(_13541_),
    .Y(_13542_));
 sky130_fd_sc_hd__or2_1 _23443_ (.A(_13537_),
    .B(_13542_),
    .X(_13543_));
 sky130_fd_sc_hd__nand2_1 _23444_ (.A(_13542_),
    .B(_13537_),
    .Y(_13545_));
 sky130_fd_sc_hd__nand2_1 _23445_ (.A(_13543_),
    .B(_13545_),
    .Y(_13546_));
 sky130_fd_sc_hd__nor2_1 _23446_ (.A(_13536_),
    .B(_13546_),
    .Y(_13547_));
 sky130_fd_sc_hd__nand2_1 _23447_ (.A(_13505_),
    .B(_13547_),
    .Y(_13548_));
 sky130_fd_sc_hd__nand2_1 _23448_ (.A(_13535_),
    .B(_11808_),
    .Y(_13549_));
 sky130_fd_sc_hd__o21a_1 _23449_ (.A1(_13543_),
    .A2(_13536_),
    .B1(_13549_),
    .X(_13550_));
 sky130_fd_sc_hd__nand2_2 _23450_ (.A(_13548_),
    .B(_13550_),
    .Y(_13551_));
 sky130_fd_sc_hd__nand2_1 _23451_ (.A(_13033_),
    .B(_13034_),
    .Y(_13552_));
 sky130_fd_sc_hd__nand2b_1 _23452_ (.A_N(_12986_),
    .B(_13552_),
    .Y(_13553_));
 sky130_fd_sc_hd__nand2b_1 _23453_ (.A_N(_13552_),
    .B(_12986_),
    .Y(_13554_));
 sky130_fd_sc_hd__nand2_1 _23454_ (.A(_13553_),
    .B(_13554_),
    .Y(_13556_));
 sky130_fd_sc_hd__or2_1 _23455_ (.A(_10749_),
    .B(_13556_),
    .X(_13557_));
 sky130_fd_sc_hd__nand2_1 _23456_ (.A(_13556_),
    .B(_10749_),
    .Y(_13558_));
 sky130_fd_sc_hd__nand2_1 _23457_ (.A(_13557_),
    .B(_13558_),
    .Y(_13559_));
 sky130_fd_sc_hd__inv_4 _23458_ (.A(_13559_),
    .Y(_13560_));
 sky130_fd_sc_hd__nand2_1 _23459_ (.A(_13508_),
    .B(_12960_),
    .Y(_13561_));
 sky130_fd_sc_hd__inv_2 _23460_ (.A(_12951_),
    .Y(_13562_));
 sky130_fd_sc_hd__nand2_1 _23461_ (.A(_13561_),
    .B(_13562_),
    .Y(_13563_));
 sky130_fd_sc_hd__nand3_1 _23462_ (.A(_13508_),
    .B(_12960_),
    .C(_12951_),
    .Y(_13564_));
 sky130_fd_sc_hd__nand2_1 _23463_ (.A(_13563_),
    .B(_13564_),
    .Y(_13565_));
 sky130_fd_sc_hd__nand2_1 _23464_ (.A(_13565_),
    .B(_12992_),
    .Y(_13567_));
 sky130_fd_sc_hd__nand3_2 _23465_ (.A(_13563_),
    .B(_11858_),
    .C(_13564_),
    .Y(_13568_));
 sky130_fd_sc_hd__nand3_1 _23466_ (.A(_13516_),
    .B(_13567_),
    .C(_13568_),
    .Y(_13569_));
 sky130_fd_sc_hd__inv_2 _23467_ (.A(_13569_),
    .Y(_13570_));
 sky130_fd_sc_hd__nand3_1 _23468_ (.A(_13481_),
    .B(_13525_),
    .C(_13570_),
    .Y(_13571_));
 sky130_fd_sc_hd__inv_2 _23469_ (.A(_13513_),
    .Y(_13572_));
 sky130_fd_sc_hd__inv_2 _23470_ (.A(_13568_),
    .Y(_13573_));
 sky130_fd_sc_hd__a21o_1 _23471_ (.A1(_13567_),
    .A2(_13572_),
    .B1(_13573_),
    .X(_13574_));
 sky130_fd_sc_hd__nor2_1 _23472_ (.A(_13528_),
    .B(_13569_),
    .Y(_13575_));
 sky130_fd_sc_hd__nor2_1 _23473_ (.A(_13574_),
    .B(_13575_),
    .Y(_13576_));
 sky130_fd_sc_hd__nand2_1 _23474_ (.A(_13571_),
    .B(_13576_),
    .Y(_13578_));
 sky130_fd_sc_hd__or2_1 _23475_ (.A(_13560_),
    .B(_13578_),
    .X(_13579_));
 sky130_fd_sc_hd__nand2_1 _23476_ (.A(_13578_),
    .B(_13560_),
    .Y(_13580_));
 sky130_fd_sc_hd__nand2_1 _23477_ (.A(_13579_),
    .B(_13580_),
    .Y(_13581_));
 sky130_fd_sc_hd__nand2_1 _23478_ (.A(_13581_),
    .B(_13483_),
    .Y(_13582_));
 sky130_fd_sc_hd__nand2_1 _23479_ (.A(\div1i.quot[6] ),
    .B(_13556_),
    .Y(_13583_));
 sky130_fd_sc_hd__nand2_1 _23480_ (.A(_13582_),
    .B(_13583_),
    .Y(_13584_));
 sky130_fd_sc_hd__nand2_1 _23481_ (.A(_13584_),
    .B(_08020_),
    .Y(_13585_));
 sky130_fd_sc_hd__nand3_1 _23482_ (.A(_13582_),
    .B(_13022_),
    .C(_13583_),
    .Y(_13586_));
 sky130_fd_sc_hd__nand2_2 _23483_ (.A(_13585_),
    .B(_13586_),
    .Y(_13587_));
 sky130_fd_sc_hd__inv_2 _23484_ (.A(_13587_),
    .Y(_13589_));
 sky130_fd_sc_hd__nand2_1 _23485_ (.A(_13567_),
    .B(_13568_),
    .Y(_13590_));
 sky130_fd_sc_hd__nand2_1 _23486_ (.A(_13531_),
    .B(_13513_),
    .Y(_13591_));
 sky130_fd_sc_hd__xor2_1 _23487_ (.A(_13590_),
    .B(_13591_),
    .X(_13592_));
 sky130_fd_sc_hd__nand2_1 _23488_ (.A(_13592_),
    .B(_13483_),
    .Y(_13593_));
 sky130_fd_sc_hd__nand2_1 _23489_ (.A(_13565_),
    .B(\div1i.quot[6] ),
    .Y(_13594_));
 sky130_fd_sc_hd__nand2_1 _23490_ (.A(_13593_),
    .B(_13594_),
    .Y(_13595_));
 sky130_fd_sc_hd__nand2_1 _23491_ (.A(_13595_),
    .B(_11896_),
    .Y(_13596_));
 sky130_fd_sc_hd__nand3_2 _23492_ (.A(_13593_),
    .B(_11899_),
    .C(_13594_),
    .Y(_13597_));
 sky130_fd_sc_hd__nand3_1 _23493_ (.A(_13589_),
    .B(_13596_),
    .C(_13597_),
    .Y(_13598_));
 sky130_fd_sc_hd__nand2_1 _23494_ (.A(_13580_),
    .B(_13557_),
    .Y(_13600_));
 sky130_fd_sc_hd__nand2_1 _23495_ (.A(_13554_),
    .B(_13034_),
    .Y(_13601_));
 sky130_fd_sc_hd__or2_1 _23496_ (.A(_13025_),
    .B(_13601_),
    .X(_13602_));
 sky130_fd_sc_hd__nand2_1 _23497_ (.A(_13601_),
    .B(_13025_),
    .Y(_13603_));
 sky130_fd_sc_hd__nand2_1 _23498_ (.A(_13602_),
    .B(_13603_),
    .Y(_13604_));
 sky130_fd_sc_hd__nand2_1 _23499_ (.A(_13604_),
    .B(_13042_),
    .Y(_13605_));
 sky130_fd_sc_hd__nand3_1 _23500_ (.A(_13602_),
    .B(_12495_),
    .C(_13603_),
    .Y(_13606_));
 sky130_fd_sc_hd__nand2_1 _23501_ (.A(_13605_),
    .B(_13606_),
    .Y(_13607_));
 sky130_fd_sc_hd__inv_2 _23502_ (.A(_13607_),
    .Y(_13608_));
 sky130_fd_sc_hd__nand2_1 _23503_ (.A(_13600_),
    .B(_13608_),
    .Y(_13609_));
 sky130_fd_sc_hd__nand3_1 _23504_ (.A(_13580_),
    .B(_13607_),
    .C(_13557_),
    .Y(_13611_));
 sky130_fd_sc_hd__nand2_1 _23505_ (.A(_13609_),
    .B(_13611_),
    .Y(_13612_));
 sky130_fd_sc_hd__nand2_1 _23506_ (.A(_13612_),
    .B(_13483_),
    .Y(_13613_));
 sky130_fd_sc_hd__nand2_1 _23507_ (.A(_13604_),
    .B(\div1i.quot[6] ),
    .Y(_13614_));
 sky130_fd_sc_hd__nand2_1 _23508_ (.A(_13613_),
    .B(_13614_),
    .Y(_13615_));
 sky130_fd_sc_hd__nand2_1 _23509_ (.A(_13615_),
    .B(_12506_),
    .Y(_13616_));
 sky130_fd_sc_hd__nand3_1 _23510_ (.A(_13613_),
    .B(_11376_),
    .C(_13614_),
    .Y(_13617_));
 sky130_fd_sc_hd__nand2_1 _23511_ (.A(_13616_),
    .B(_13617_),
    .Y(_13618_));
 sky130_fd_sc_hd__inv_2 _23512_ (.A(_13618_),
    .Y(_13619_));
 sky130_fd_sc_hd__nand2_1 _23513_ (.A(_13608_),
    .B(_13560_),
    .Y(_13620_));
 sky130_fd_sc_hd__inv_2 _23514_ (.A(_13620_),
    .Y(_13622_));
 sky130_fd_sc_hd__nand2_1 _23515_ (.A(_13578_),
    .B(_13622_),
    .Y(_13623_));
 sky130_fd_sc_hd__o21a_1 _23516_ (.A1(_13557_),
    .A2(_13607_),
    .B1(_13606_),
    .X(_13624_));
 sky130_fd_sc_hd__nand2_1 _23517_ (.A(_13623_),
    .B(_13624_),
    .Y(_13625_));
 sky130_fd_sc_hd__a41o_1 _23518_ (.A1(_12986_),
    .A2(_13025_),
    .A3(_13034_),
    .A4(_13033_),
    .B1(_13087_),
    .X(_13626_));
 sky130_fd_sc_hd__or2_1 _23519_ (.A(_13056_),
    .B(_13626_),
    .X(_13627_));
 sky130_fd_sc_hd__nand2_1 _23520_ (.A(_13626_),
    .B(_13056_),
    .Y(_13628_));
 sky130_fd_sc_hd__nand2_1 _23521_ (.A(_13627_),
    .B(_13628_),
    .Y(_13629_));
 sky130_fd_sc_hd__inv_2 _23522_ (.A(_13629_),
    .Y(_13630_));
 sky130_fd_sc_hd__nand2_1 _23523_ (.A(_13630_),
    .B(_11935_),
    .Y(_13631_));
 sky130_fd_sc_hd__buf_6 _23524_ (.A(_08611_),
    .X(_13633_));
 sky130_fd_sc_hd__nand2_1 _23525_ (.A(_13629_),
    .B(_13633_),
    .Y(_13634_));
 sky130_fd_sc_hd__nand2_1 _23526_ (.A(_13631_),
    .B(_13634_),
    .Y(_13635_));
 sky130_fd_sc_hd__inv_2 _23527_ (.A(_13635_),
    .Y(_13636_));
 sky130_fd_sc_hd__nand2_1 _23528_ (.A(_13625_),
    .B(_13636_),
    .Y(_13637_));
 sky130_fd_sc_hd__nand3_1 _23529_ (.A(_13623_),
    .B(_13635_),
    .C(_13624_),
    .Y(_13638_));
 sky130_fd_sc_hd__nand3_1 _23530_ (.A(_13637_),
    .B(_13638_),
    .C(_13483_),
    .Y(_13639_));
 sky130_fd_sc_hd__nand2_1 _23531_ (.A(_13630_),
    .B(\div1i.quot[6] ),
    .Y(_13640_));
 sky130_fd_sc_hd__nand2_1 _23532_ (.A(_13639_),
    .B(_13640_),
    .Y(_13641_));
 sky130_fd_sc_hd__nand2_1 _23533_ (.A(_13641_),
    .B(_11946_),
    .Y(_13642_));
 sky130_fd_sc_hd__nand3_1 _23534_ (.A(_13639_),
    .B(_11948_),
    .C(_13640_),
    .Y(_13644_));
 sky130_fd_sc_hd__nand2_2 _23535_ (.A(_13642_),
    .B(_13644_),
    .Y(_13645_));
 sky130_fd_sc_hd__inv_2 _23536_ (.A(_13645_),
    .Y(_13646_));
 sky130_fd_sc_hd__nand2_1 _23537_ (.A(_13619_),
    .B(_13646_),
    .Y(_13647_));
 sky130_fd_sc_hd__nor2_1 _23538_ (.A(_13598_),
    .B(_13647_),
    .Y(_13648_));
 sky130_fd_sc_hd__nand2_4 _23539_ (.A(_13551_),
    .B(_13648_),
    .Y(_13649_));
 sky130_fd_sc_hd__o21ai_1 _23540_ (.A1(_13597_),
    .A2(_13587_),
    .B1(_13586_),
    .Y(_13650_));
 sky130_fd_sc_hd__nor2_1 _23541_ (.A(_13645_),
    .B(_13618_),
    .Y(_13651_));
 sky130_fd_sc_hd__o21ai_1 _23542_ (.A1(_13617_),
    .A2(_13645_),
    .B1(_13642_),
    .Y(_13652_));
 sky130_fd_sc_hd__a21oi_2 _23543_ (.A1(_13650_),
    .A2(_13651_),
    .B1(_13652_),
    .Y(_13653_));
 sky130_fd_sc_hd__nand2_4 _23544_ (.A(_13649_),
    .B(_13653_),
    .Y(_13655_));
 sky130_fd_sc_hd__nand2_1 _23545_ (.A(_13628_),
    .B(_13054_),
    .Y(_13656_));
 sky130_fd_sc_hd__xor2_2 _23546_ (.A(_13081_),
    .B(_13656_),
    .X(_13657_));
 sky130_fd_sc_hd__nand3_1 _23547_ (.A(_13637_),
    .B(_13483_),
    .C(_13631_),
    .Y(_13658_));
 sky130_fd_sc_hd__xnor2_2 _23548_ (.A(_13657_),
    .B(_13658_),
    .Y(_13659_));
 sky130_fd_sc_hd__nand2_8 _23549_ (.A(_13655_),
    .B(_13659_),
    .Y(_13660_));
 sky130_fd_sc_hd__clkinvlp_2 _23550_ (.A(_13659_),
    .Y(_13661_));
 sky130_fd_sc_hd__nand3_4 _23551_ (.A(_13649_),
    .B(_13653_),
    .C(_13661_),
    .Y(_13662_));
 sky130_fd_sc_hd__nand2_8 _23552_ (.A(_13660_),
    .B(_13662_),
    .Y(_13663_));
 sky130_fd_sc_hd__buf_8 _23553_ (.A(_13663_),
    .X(_13664_));
 sky130_fd_sc_hd__buf_8 _23554_ (.A(net226),
    .X(\div1i.quot[5] ));
 sky130_fd_sc_hd__nand2_1 _23555_ (.A(_13326_),
    .B(_13329_),
    .Y(_13666_));
 sky130_fd_sc_hd__nand2_1 _23556_ (.A(_13666_),
    .B(_13330_),
    .Y(_13667_));
 sky130_fd_sc_hd__nand2_1 _23557_ (.A(_13667_),
    .B(_13332_),
    .Y(_13668_));
 sky130_fd_sc_hd__inv_2 _23558_ (.A(_13668_),
    .Y(_13669_));
 sky130_fd_sc_hd__nand2_1 _23559_ (.A(_13664_),
    .B(_13669_),
    .Y(_13670_));
 sky130_fd_sc_hd__o21ai_1 _23560_ (.A1(_12032_),
    .A2(\div1i.quot[6] ),
    .B1(_12033_),
    .Y(_13671_));
 sky130_fd_sc_hd__nand2_1 _23561_ (.A(_13668_),
    .B(_12030_),
    .Y(_13672_));
 sky130_fd_sc_hd__nand3_1 _23562_ (.A(_13667_),
    .B(_12035_),
    .C(_13332_),
    .Y(_13673_));
 sky130_fd_sc_hd__nand2_1 _23563_ (.A(_13672_),
    .B(_13673_),
    .Y(_13674_));
 sky130_fd_sc_hd__xor2_1 _23564_ (.A(_13671_),
    .B(_13674_),
    .X(_13676_));
 sky130_fd_sc_hd__nand3b_1 _23565_ (.A_N(_13676_),
    .B(_13660_),
    .C(_13662_),
    .Y(_13677_));
 sky130_fd_sc_hd__nand2_1 _23566_ (.A(_13670_),
    .B(_13677_),
    .Y(_13678_));
 sky130_fd_sc_hd__buf_6 _23567_ (.A(_11069_),
    .X(_13679_));
 sky130_fd_sc_hd__nand2_1 _23568_ (.A(_13678_),
    .B(_13679_),
    .Y(_13680_));
 sky130_fd_sc_hd__nor2_1 _23569_ (.A(_12032_),
    .B(_13483_),
    .Y(_13681_));
 sky130_fd_sc_hd__or2_1 _23570_ (.A(_11412_),
    .B(_13681_),
    .X(_13682_));
 sky130_fd_sc_hd__nand2_1 _23571_ (.A(_13682_),
    .B(_13330_),
    .Y(_13683_));
 sky130_fd_sc_hd__clkinvlp_2 _23572_ (.A(_13683_),
    .Y(_13684_));
 sky130_fd_sc_hd__nand2_2 _23573_ (.A(_13664_),
    .B(_13684_),
    .Y(_13685_));
 sky130_fd_sc_hd__nand3_1 _23574_ (.A(_13660_),
    .B(_13662_),
    .C(_13681_),
    .Y(_13687_));
 sky130_fd_sc_hd__nand2_2 _23575_ (.A(_13685_),
    .B(_13687_),
    .Y(_13688_));
 sky130_fd_sc_hd__nand2_4 _23576_ (.A(_13688_),
    .B(_11421_),
    .Y(_13689_));
 sky130_fd_sc_hd__nand2_2 _23577_ (.A(_13680_),
    .B(_13689_),
    .Y(_13690_));
 sky130_fd_sc_hd__inv_2 _23578_ (.A(_13690_),
    .Y(_13691_));
 sky130_fd_sc_hd__nand3_2 _23579_ (.A(_13685_),
    .B(_11426_),
    .C(_13687_),
    .Y(_13692_));
 sky130_fd_sc_hd__nand3_2 _23580_ (.A(_13664_),
    .B(_12033_),
    .C(_12221_),
    .Y(_13693_));
 sky130_fd_sc_hd__inv_2 _23581_ (.A(_13693_),
    .Y(_13694_));
 sky130_fd_sc_hd__nand3_4 _23582_ (.A(_13689_),
    .B(_13692_),
    .C(_13694_),
    .Y(_13695_));
 sky130_fd_sc_hd__or2_4 _23583_ (.A(_13679_),
    .B(_13678_),
    .X(_13696_));
 sky130_fd_sc_hd__inv_2 _23584_ (.A(_13696_),
    .Y(_13698_));
 sky130_fd_sc_hd__a21oi_2 _23585_ (.A1(_13691_),
    .A2(_13695_),
    .B1(_13698_),
    .Y(_13699_));
 sky130_fd_sc_hd__inv_2 _23586_ (.A(_13388_),
    .Y(_13700_));
 sky130_fd_sc_hd__o21ai_1 _23587_ (.A1(_13384_),
    .A2(_13336_),
    .B1(_13700_),
    .Y(_13701_));
 sky130_fd_sc_hd__or2_1 _23588_ (.A(_13360_),
    .B(_13701_),
    .X(_13702_));
 sky130_fd_sc_hd__nand2_1 _23589_ (.A(_13701_),
    .B(_13360_),
    .Y(_13703_));
 sky130_fd_sc_hd__nand2_1 _23590_ (.A(_13702_),
    .B(_13703_),
    .Y(_13704_));
 sky130_fd_sc_hd__inv_2 _23591_ (.A(_13704_),
    .Y(_13705_));
 sky130_fd_sc_hd__nand2_1 _23592_ (.A(_13663_),
    .B(_13705_),
    .Y(_13706_));
 sky130_fd_sc_hd__nand2_1 _23593_ (.A(_13705_),
    .B(_12087_),
    .Y(_13707_));
 sky130_fd_sc_hd__nand2_1 _23594_ (.A(_13704_),
    .B(_12085_),
    .Y(_13709_));
 sky130_fd_sc_hd__nand2_1 _23595_ (.A(_13707_),
    .B(_13709_),
    .Y(_13710_));
 sky130_fd_sc_hd__inv_2 _23596_ (.A(_13710_),
    .Y(_13711_));
 sky130_fd_sc_hd__nand2_1 _23597_ (.A(_13337_),
    .B(_13383_),
    .Y(_13712_));
 sky130_fd_sc_hd__nand2_1 _23598_ (.A(_13336_),
    .B(_13382_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand2_1 _23599_ (.A(_13712_),
    .B(_13713_),
    .Y(_13714_));
 sky130_fd_sc_hd__nand2_1 _23600_ (.A(_13714_),
    .B(_12056_),
    .Y(_13715_));
 sky130_fd_sc_hd__nand3_1 _23601_ (.A(_13712_),
    .B(_12058_),
    .C(_13713_),
    .Y(_13716_));
 sky130_fd_sc_hd__nand2_1 _23602_ (.A(_13715_),
    .B(_13716_),
    .Y(_13717_));
 sky130_fd_sc_hd__inv_2 _23603_ (.A(_13717_),
    .Y(_13718_));
 sky130_fd_sc_hd__inv_2 _23604_ (.A(_13673_),
    .Y(_13720_));
 sky130_fd_sc_hd__a21o_1 _23605_ (.A1(_13672_),
    .A2(_13671_),
    .B1(_13720_),
    .X(_13721_));
 sky130_fd_sc_hd__nand2_1 _23606_ (.A(_13334_),
    .B(_13317_),
    .Y(_13722_));
 sky130_fd_sc_hd__nand2_1 _23607_ (.A(_13332_),
    .B(_13326_),
    .Y(_13723_));
 sky130_fd_sc_hd__xor2_1 _23608_ (.A(_13722_),
    .B(_13723_),
    .X(_13724_));
 sky130_fd_sc_hd__nand2_1 _23609_ (.A(_13724_),
    .B(_12043_),
    .Y(_13725_));
 sky130_fd_sc_hd__nand2_1 _23610_ (.A(_13721_),
    .B(_13725_),
    .Y(_13726_));
 sky130_fd_sc_hd__inv_2 _23611_ (.A(_13724_),
    .Y(_13727_));
 sky130_fd_sc_hd__nand2_1 _23612_ (.A(_13727_),
    .B(_12047_),
    .Y(_13728_));
 sky130_fd_sc_hd__nand2_1 _23613_ (.A(_13726_),
    .B(_13728_),
    .Y(_13729_));
 sky130_fd_sc_hd__nand2_1 _23614_ (.A(_13718_),
    .B(_13729_),
    .Y(_13731_));
 sky130_fd_sc_hd__nand2_1 _23615_ (.A(_13731_),
    .B(_13716_),
    .Y(_13732_));
 sky130_fd_sc_hd__nand2_1 _23616_ (.A(_13712_),
    .B(_13380_),
    .Y(_13733_));
 sky130_fd_sc_hd__xor2_2 _23617_ (.A(_13372_),
    .B(_13733_),
    .X(_13734_));
 sky130_fd_sc_hd__nand2_1 _23618_ (.A(_13734_),
    .B(_13182_),
    .Y(_13735_));
 sky130_fd_sc_hd__nand2_1 _23619_ (.A(_13732_),
    .B(_13735_),
    .Y(_13736_));
 sky130_fd_sc_hd__inv_4 _23620_ (.A(_13734_),
    .Y(_13737_));
 sky130_fd_sc_hd__nand2_1 _23621_ (.A(_13737_),
    .B(_08176_),
    .Y(_13738_));
 sky130_fd_sc_hd__nand2_1 _23622_ (.A(_13736_),
    .B(_13738_),
    .Y(_13739_));
 sky130_fd_sc_hd__or2_1 _23623_ (.A(_13711_),
    .B(_13739_),
    .X(_13740_));
 sky130_fd_sc_hd__nand2_1 _23624_ (.A(_13739_),
    .B(_13711_),
    .Y(_13742_));
 sky130_fd_sc_hd__nand2_1 _23625_ (.A(_13740_),
    .B(_13742_),
    .Y(_13743_));
 sky130_fd_sc_hd__inv_2 _23626_ (.A(_13743_),
    .Y(_13744_));
 sky130_fd_sc_hd__nand3_1 _23627_ (.A(_13660_),
    .B(_13662_),
    .C(_13744_),
    .Y(_13745_));
 sky130_fd_sc_hd__nand2_1 _23628_ (.A(_13706_),
    .B(_13745_),
    .Y(_13746_));
 sky130_fd_sc_hd__nand2_1 _23629_ (.A(_13746_),
    .B(_11482_),
    .Y(_13747_));
 sky130_fd_sc_hd__nand3_1 _23630_ (.A(_13706_),
    .B(_11484_),
    .C(_13745_),
    .Y(_13748_));
 sky130_fd_sc_hd__nand2_1 _23631_ (.A(_13747_),
    .B(_13748_),
    .Y(_13749_));
 sky130_fd_sc_hd__inv_2 _23632_ (.A(_13749_),
    .Y(_13750_));
 sky130_fd_sc_hd__nand2_1 _23633_ (.A(_13663_),
    .B(_13737_),
    .Y(_13751_));
 sky130_fd_sc_hd__nand2_1 _23634_ (.A(_13738_),
    .B(_13735_),
    .Y(_13753_));
 sky130_fd_sc_hd__xnor2_1 _23635_ (.A(_13732_),
    .B(_13753_),
    .Y(_13754_));
 sky130_fd_sc_hd__nand3_1 _23636_ (.A(_13660_),
    .B(_13662_),
    .C(_13754_),
    .Y(_13755_));
 sky130_fd_sc_hd__nand2_1 _23637_ (.A(_13751_),
    .B(_13755_),
    .Y(_13756_));
 sky130_fd_sc_hd__nand2_1 _23638_ (.A(_13756_),
    .B(_11494_),
    .Y(_13757_));
 sky130_fd_sc_hd__nand3_1 _23639_ (.A(_13751_),
    .B(_11496_),
    .C(_13755_),
    .Y(_13758_));
 sky130_fd_sc_hd__nand2_2 _23640_ (.A(_13757_),
    .B(_13758_),
    .Y(_13759_));
 sky130_fd_sc_hd__inv_2 _23641_ (.A(_13759_),
    .Y(_13760_));
 sky130_fd_sc_hd__nand2_1 _23642_ (.A(_13750_),
    .B(_13760_),
    .Y(_13761_));
 sky130_fd_sc_hd__inv_2 _23643_ (.A(_13714_),
    .Y(_13762_));
 sky130_fd_sc_hd__nand2_1 _23644_ (.A(_13663_),
    .B(_13762_),
    .Y(_13764_));
 sky130_fd_sc_hd__or2_1 _23645_ (.A(_13729_),
    .B(_13718_),
    .X(_13765_));
 sky130_fd_sc_hd__nand2_1 _23646_ (.A(_13765_),
    .B(_13731_),
    .Y(_13766_));
 sky130_fd_sc_hd__inv_2 _23647_ (.A(_13766_),
    .Y(_13767_));
 sky130_fd_sc_hd__nand3_1 _23648_ (.A(_13660_),
    .B(_13662_),
    .C(_13767_),
    .Y(_13768_));
 sky130_fd_sc_hd__nand2_1 _23649_ (.A(_13764_),
    .B(_13768_),
    .Y(_13769_));
 sky130_fd_sc_hd__nand2_1 _23650_ (.A(_13769_),
    .B(_11105_),
    .Y(_13770_));
 sky130_fd_sc_hd__nand3_1 _23651_ (.A(_13764_),
    .B(_12261_),
    .C(_13768_),
    .Y(_13771_));
 sky130_fd_sc_hd__nand2_2 _23652_ (.A(_13770_),
    .B(_13771_),
    .Y(_13772_));
 sky130_fd_sc_hd__inv_2 _23653_ (.A(_13772_),
    .Y(_13773_));
 sky130_fd_sc_hd__nand2_1 _23654_ (.A(_13663_),
    .B(_13727_),
    .Y(_13775_));
 sky130_fd_sc_hd__nand2_1 _23655_ (.A(_13728_),
    .B(_13725_),
    .Y(_13776_));
 sky130_fd_sc_hd__xnor2_1 _23656_ (.A(_13721_),
    .B(_13776_),
    .Y(_13777_));
 sky130_fd_sc_hd__nand3_1 _23657_ (.A(_13660_),
    .B(_13662_),
    .C(_13777_),
    .Y(_13778_));
 sky130_fd_sc_hd__nand2_1 _23658_ (.A(_13775_),
    .B(_13778_),
    .Y(_13779_));
 sky130_fd_sc_hd__nand2_1 _23659_ (.A(_13779_),
    .B(_12270_),
    .Y(_13780_));
 sky130_fd_sc_hd__nand3_1 _23660_ (.A(_13775_),
    .B(_11117_),
    .C(_13778_),
    .Y(_13781_));
 sky130_fd_sc_hd__nand2_1 _23661_ (.A(_13780_),
    .B(_13781_),
    .Y(_13782_));
 sky130_fd_sc_hd__inv_2 _23662_ (.A(_13782_),
    .Y(_13783_));
 sky130_fd_sc_hd__nand2_1 _23663_ (.A(_13773_),
    .B(_13783_),
    .Y(_13784_));
 sky130_fd_sc_hd__nor2_1 _23664_ (.A(_13761_),
    .B(_13784_),
    .Y(_13786_));
 sky130_fd_sc_hd__nand2_1 _23665_ (.A(_13699_),
    .B(_13786_),
    .Y(_13787_));
 sky130_fd_sc_hd__inv_2 _23666_ (.A(_13771_),
    .Y(_13788_));
 sky130_fd_sc_hd__o21ai_2 _23667_ (.A1(_13780_),
    .A2(_13788_),
    .B1(_13770_),
    .Y(_13789_));
 sky130_fd_sc_hd__nor2_1 _23668_ (.A(_13749_),
    .B(_13759_),
    .Y(_13790_));
 sky130_fd_sc_hd__inv_2 _23669_ (.A(_13748_),
    .Y(_13791_));
 sky130_fd_sc_hd__o21ai_1 _23670_ (.A1(_13757_),
    .A2(_13791_),
    .B1(_13747_),
    .Y(_13792_));
 sky130_fd_sc_hd__a21oi_1 _23671_ (.A1(_13789_),
    .A2(_13790_),
    .B1(_13792_),
    .Y(_13793_));
 sky130_fd_sc_hd__nand2_2 _23672_ (.A(_13787_),
    .B(_13793_),
    .Y(_13794_));
 sky130_fd_sc_hd__inv_2 _23673_ (.A(_13416_),
    .Y(_13795_));
 sky130_fd_sc_hd__nand2_1 _23674_ (.A(_13394_),
    .B(_13795_),
    .Y(_13797_));
 sky130_fd_sc_hd__inv_2 _23675_ (.A(_13440_),
    .Y(_13798_));
 sky130_fd_sc_hd__nand2_1 _23676_ (.A(_13797_),
    .B(_13798_),
    .Y(_13799_));
 sky130_fd_sc_hd__inv_2 _23677_ (.A(_13427_),
    .Y(_13800_));
 sky130_fd_sc_hd__nand2_1 _23678_ (.A(_13799_),
    .B(_13800_),
    .Y(_13801_));
 sky130_fd_sc_hd__nand3_1 _23679_ (.A(_13797_),
    .B(_13427_),
    .C(_13798_),
    .Y(_13802_));
 sky130_fd_sc_hd__nand2_1 _23680_ (.A(_13801_),
    .B(_13802_),
    .Y(_13803_));
 sky130_fd_sc_hd__inv_2 _23681_ (.A(_13803_),
    .Y(_13804_));
 sky130_fd_sc_hd__nand2_1 _23682_ (.A(_13804_),
    .B(_11986_),
    .Y(_13805_));
 sky130_fd_sc_hd__nand2_1 _23683_ (.A(_13803_),
    .B(_12017_),
    .Y(_13806_));
 sky130_fd_sc_hd__nand2_1 _23684_ (.A(_13805_),
    .B(_13806_),
    .Y(_13808_));
 sky130_fd_sc_hd__inv_2 _23685_ (.A(_13808_),
    .Y(_13809_));
 sky130_fd_sc_hd__nand2_1 _23686_ (.A(_13703_),
    .B(_13358_),
    .Y(_13810_));
 sky130_fd_sc_hd__or2_1 _23687_ (.A(_13350_),
    .B(_13810_),
    .X(_13811_));
 sky130_fd_sc_hd__nand2_1 _23688_ (.A(_13810_),
    .B(_13350_),
    .Y(_13812_));
 sky130_fd_sc_hd__nand3_1 _23689_ (.A(_13811_),
    .B(_10939_),
    .C(_13812_),
    .Y(_13813_));
 sky130_fd_sc_hd__nand2_1 _23690_ (.A(_13813_),
    .B(_13707_),
    .Y(_13814_));
 sky130_fd_sc_hd__inv_2 _23691_ (.A(_13814_),
    .Y(_13815_));
 sky130_fd_sc_hd__nand2_1 _23692_ (.A(_13742_),
    .B(_13815_),
    .Y(_13816_));
 sky130_fd_sc_hd__nand2_2 _23693_ (.A(_13394_),
    .B(_13415_),
    .Y(_13817_));
 sky130_fd_sc_hd__nand2_2 _23694_ (.A(_13817_),
    .B(_13413_),
    .Y(_13819_));
 sky130_fd_sc_hd__xor2_1 _23695_ (.A(_13403_),
    .B(_13819_),
    .X(_13820_));
 sky130_fd_sc_hd__nand2_2 _23696_ (.A(_13820_),
    .B(_12002_),
    .Y(_13821_));
 sky130_fd_sc_hd__or2_1 _23697_ (.A(_13404_),
    .B(_13819_),
    .X(_13822_));
 sky130_fd_sc_hd__nand2_1 _23698_ (.A(_13819_),
    .B(_13404_),
    .Y(_13823_));
 sky130_fd_sc_hd__nand3_1 _23699_ (.A(_13822_),
    .B(_12012_),
    .C(_13823_),
    .Y(_13824_));
 sky130_fd_sc_hd__or2_1 _23700_ (.A(_13415_),
    .B(_13394_),
    .X(_13825_));
 sky130_fd_sc_hd__nand2_1 _23701_ (.A(_13825_),
    .B(_13817_),
    .Y(_13826_));
 sky130_fd_sc_hd__nand2_1 _23702_ (.A(_13826_),
    .B(_12101_),
    .Y(_13827_));
 sky130_fd_sc_hd__nand3_2 _23703_ (.A(_13825_),
    .B(_12008_),
    .C(_13817_),
    .Y(_13828_));
 sky130_fd_sc_hd__nand2_1 _23704_ (.A(_13827_),
    .B(_13828_),
    .Y(_13830_));
 sky130_fd_sc_hd__inv_2 _23705_ (.A(_13830_),
    .Y(_13831_));
 sky130_fd_sc_hd__nand3_1 _23706_ (.A(_13821_),
    .B(_13824_),
    .C(_13831_),
    .Y(_13832_));
 sky130_fd_sc_hd__inv_2 _23707_ (.A(_13832_),
    .Y(_13833_));
 sky130_fd_sc_hd__nand2_1 _23708_ (.A(_13811_),
    .B(_13812_),
    .Y(_13834_));
 sky130_fd_sc_hd__nand2_1 _23709_ (.A(_13834_),
    .B(_13197_),
    .Y(_13835_));
 sky130_fd_sc_hd__nand3_2 _23710_ (.A(_13816_),
    .B(_13833_),
    .C(_13835_),
    .Y(_13836_));
 sky130_fd_sc_hd__clkinvlp_2 _23711_ (.A(_13828_),
    .Y(_13837_));
 sky130_fd_sc_hd__a21boi_2 _23712_ (.A1(_13821_),
    .A2(_13837_),
    .B1_N(_13824_),
    .Y(_13838_));
 sky130_fd_sc_hd__nand2_1 _23713_ (.A(_13836_),
    .B(_13838_),
    .Y(_13839_));
 sky130_fd_sc_hd__or2_1 _23714_ (.A(_13809_),
    .B(_13839_),
    .X(_13841_));
 sky130_fd_sc_hd__inv_6 _23715_ (.A(_13663_),
    .Y(_13842_));
 sky130_fd_sc_hd__nand2_1 _23716_ (.A(_13839_),
    .B(_13809_),
    .Y(_13843_));
 sky130_fd_sc_hd__nand3_1 _23717_ (.A(_13841_),
    .B(_13842_),
    .C(_13843_),
    .Y(_13844_));
 sky130_fd_sc_hd__nand2_1 _23718_ (.A(net226),
    .B(_13804_),
    .Y(_13845_));
 sky130_fd_sc_hd__nand2_1 _23719_ (.A(_13844_),
    .B(_13845_),
    .Y(_13846_));
 sky130_fd_sc_hd__nand2_1 _23720_ (.A(_13846_),
    .B(_11586_),
    .Y(_13847_));
 sky130_fd_sc_hd__nand3_1 _23721_ (.A(_13844_),
    .B(_11588_),
    .C(_13845_),
    .Y(_13848_));
 sky130_fd_sc_hd__nand2_2 _23722_ (.A(_13847_),
    .B(_13848_),
    .Y(_13849_));
 sky130_fd_sc_hd__nand3_1 _23723_ (.A(_13816_),
    .B(_13835_),
    .C(_13831_),
    .Y(_13850_));
 sky130_fd_sc_hd__nand2_1 _23724_ (.A(_13850_),
    .B(_13828_),
    .Y(_13852_));
 sky130_fd_sc_hd__nand3_1 _23725_ (.A(_13852_),
    .B(_13824_),
    .C(_13821_),
    .Y(_13853_));
 sky130_fd_sc_hd__nand2_1 _23726_ (.A(_13821_),
    .B(_13824_),
    .Y(_13854_));
 sky130_fd_sc_hd__nand3_1 _23727_ (.A(_13850_),
    .B(_13854_),
    .C(_13828_),
    .Y(_13855_));
 sky130_fd_sc_hd__a21o_1 _23728_ (.A1(_13853_),
    .A2(_13855_),
    .B1(_13664_),
    .X(_13856_));
 sky130_fd_sc_hd__nand2_2 _23729_ (.A(net226),
    .B(_13820_),
    .Y(_13857_));
 sky130_fd_sc_hd__nand2_1 _23730_ (.A(_13856_),
    .B(_13857_),
    .Y(_13858_));
 sky130_fd_sc_hd__nand2_1 _23731_ (.A(_13858_),
    .B(_11600_),
    .Y(_13859_));
 sky130_fd_sc_hd__nand3_4 _23732_ (.A(_13856_),
    .B(_11603_),
    .C(_13857_),
    .Y(_13860_));
 sky130_fd_sc_hd__nand2_2 _23733_ (.A(_13859_),
    .B(_13860_),
    .Y(_13861_));
 sky130_fd_sc_hd__nor2_2 _23734_ (.A(_13861_),
    .B(_13849_),
    .Y(_13863_));
 sky130_fd_sc_hd__a21o_1 _23735_ (.A1(_13816_),
    .A2(_13835_),
    .B1(_13831_),
    .X(_13864_));
 sky130_fd_sc_hd__nand3_1 _23736_ (.A(_13842_),
    .B(_13850_),
    .C(_13864_),
    .Y(_13865_));
 sky130_fd_sc_hd__a21o_1 _23737_ (.A1(_13660_),
    .A2(_13662_),
    .B1(_13826_),
    .X(_13866_));
 sky130_fd_sc_hd__nand2_1 _23738_ (.A(_13865_),
    .B(_13866_),
    .Y(_13867_));
 sky130_fd_sc_hd__nand2_1 _23739_ (.A(_13867_),
    .B(_11614_),
    .Y(_13868_));
 sky130_fd_sc_hd__nand3_1 _23740_ (.A(_13865_),
    .B(_11616_),
    .C(_13866_),
    .Y(_13869_));
 sky130_fd_sc_hd__nand2_1 _23741_ (.A(_13868_),
    .B(_13869_),
    .Y(_13870_));
 sky130_fd_sc_hd__nand2_1 _23742_ (.A(_13835_),
    .B(_13813_),
    .Y(_13871_));
 sky130_fd_sc_hd__nand2_1 _23743_ (.A(_13742_),
    .B(_13707_),
    .Y(_13872_));
 sky130_fd_sc_hd__xor2_1 _23744_ (.A(_13871_),
    .B(_13872_),
    .X(_13874_));
 sky130_fd_sc_hd__nand2_1 _23745_ (.A(_13842_),
    .B(_13874_),
    .Y(_13875_));
 sky130_fd_sc_hd__nand2_1 _23746_ (.A(_13664_),
    .B(_13834_),
    .Y(_13876_));
 sky130_fd_sc_hd__nand2_1 _23747_ (.A(_13875_),
    .B(_13876_),
    .Y(_13877_));
 sky130_fd_sc_hd__or2_4 _23748_ (.A(_12771_),
    .B(_13877_),
    .X(_13878_));
 sky130_fd_sc_hd__nand2_1 _23749_ (.A(_13877_),
    .B(_12771_),
    .Y(_13879_));
 sky130_fd_sc_hd__nand2_1 _23750_ (.A(_13878_),
    .B(_13879_),
    .Y(_13880_));
 sky130_fd_sc_hd__nor2_2 _23751_ (.A(_13870_),
    .B(_13880_),
    .Y(_13881_));
 sky130_fd_sc_hd__nand2_1 _23752_ (.A(_13863_),
    .B(_13881_),
    .Y(_13882_));
 sky130_fd_sc_hd__inv_2 _23753_ (.A(_13882_),
    .Y(_13883_));
 sky130_fd_sc_hd__nand2_1 _23754_ (.A(_13794_),
    .B(_13883_),
    .Y(_13885_));
 sky130_fd_sc_hd__o21ai_2 _23755_ (.A1(_13878_),
    .A2(_13870_),
    .B1(_13868_),
    .Y(_13886_));
 sky130_fd_sc_hd__o21ai_1 _23756_ (.A1(_13860_),
    .A2(_13849_),
    .B1(_13847_),
    .Y(_13887_));
 sky130_fd_sc_hd__a21oi_1 _23757_ (.A1(_13886_),
    .A2(_13863_),
    .B1(_13887_),
    .Y(_13888_));
 sky130_fd_sc_hd__nand2_2 _23758_ (.A(_13885_),
    .B(_13888_),
    .Y(_13889_));
 sky130_fd_sc_hd__inv_2 _23759_ (.A(_13836_),
    .Y(_13890_));
 sky130_fd_sc_hd__nand2_1 _23760_ (.A(_13801_),
    .B(_13426_),
    .Y(_13891_));
 sky130_fd_sc_hd__inv_2 _23761_ (.A(_13435_),
    .Y(_13892_));
 sky130_fd_sc_hd__nand2_1 _23762_ (.A(_13891_),
    .B(_13892_),
    .Y(_13893_));
 sky130_fd_sc_hd__nand3_1 _23763_ (.A(_13801_),
    .B(_13435_),
    .C(_13426_),
    .Y(_13894_));
 sky130_fd_sc_hd__nand2_1 _23764_ (.A(_13893_),
    .B(_13894_),
    .Y(_13896_));
 sky130_fd_sc_hd__nand2_1 _23765_ (.A(_13896_),
    .B(_11983_),
    .Y(_13897_));
 sky130_fd_sc_hd__nand3_1 _23766_ (.A(_13893_),
    .B(_11990_),
    .C(_13894_),
    .Y(_13898_));
 sky130_fd_sc_hd__nand3_1 _23767_ (.A(_13809_),
    .B(_13897_),
    .C(_13898_),
    .Y(_13899_));
 sky130_fd_sc_hd__inv_2 _23768_ (.A(_13899_),
    .Y(_13900_));
 sky130_fd_sc_hd__nand2_1 _23769_ (.A(_13890_),
    .B(_13900_),
    .Y(_13901_));
 sky130_fd_sc_hd__nor2_1 _23770_ (.A(_13838_),
    .B(_13899_),
    .Y(_13902_));
 sky130_fd_sc_hd__nand2_1 _23771_ (.A(_13897_),
    .B(_13898_),
    .Y(_13903_));
 sky130_fd_sc_hd__o21ai_1 _23772_ (.A1(_13805_),
    .A2(_13903_),
    .B1(_13898_),
    .Y(_13904_));
 sky130_fd_sc_hd__nor2_1 _23773_ (.A(_13902_),
    .B(_13904_),
    .Y(_13905_));
 sky130_fd_sc_hd__nand2_1 _23774_ (.A(_13901_),
    .B(_13905_),
    .Y(_13907_));
 sky130_fd_sc_hd__inv_2 _23775_ (.A(_13449_),
    .Y(_13908_));
 sky130_fd_sc_hd__inv_2 _23776_ (.A(_13448_),
    .Y(_13909_));
 sky130_fd_sc_hd__nand2_1 _23777_ (.A(_13444_),
    .B(_13909_),
    .Y(_13910_));
 sky130_fd_sc_hd__nand2_1 _23778_ (.A(_13910_),
    .B(_13297_),
    .Y(_13911_));
 sky130_fd_sc_hd__or2_1 _23779_ (.A(_13908_),
    .B(_13911_),
    .X(_13912_));
 sky130_fd_sc_hd__nand2_1 _23780_ (.A(_13911_),
    .B(_13908_),
    .Y(_13913_));
 sky130_fd_sc_hd__nand2_1 _23781_ (.A(_13912_),
    .B(_13913_),
    .Y(_13914_));
 sky130_fd_sc_hd__nand2_1 _23782_ (.A(_13914_),
    .B(_12118_),
    .Y(_13915_));
 sky130_fd_sc_hd__nand3_1 _23783_ (.A(_13912_),
    .B(_12120_),
    .C(_13913_),
    .Y(_13916_));
 sky130_fd_sc_hd__nand2_1 _23784_ (.A(_13915_),
    .B(_13916_),
    .Y(_13918_));
 sky130_fd_sc_hd__inv_2 _23785_ (.A(_13918_),
    .Y(_13919_));
 sky130_fd_sc_hd__or2_1 _23786_ (.A(_13909_),
    .B(_13444_),
    .X(_13920_));
 sky130_fd_sc_hd__nand2_1 _23787_ (.A(_13920_),
    .B(_13910_),
    .Y(_13921_));
 sky130_fd_sc_hd__inv_2 _23788_ (.A(_13921_),
    .Y(_13922_));
 sky130_fd_sc_hd__nand2_1 _23789_ (.A(_13922_),
    .B(_11671_),
    .Y(_13923_));
 sky130_fd_sc_hd__nand2_1 _23790_ (.A(_13921_),
    .B(_12817_),
    .Y(_13924_));
 sky130_fd_sc_hd__nand2_2 _23791_ (.A(_13923_),
    .B(_13924_),
    .Y(_13925_));
 sky130_fd_sc_hd__inv_4 _23792_ (.A(_13925_),
    .Y(_13926_));
 sky130_fd_sc_hd__nand2_1 _23793_ (.A(_13919_),
    .B(_13926_),
    .Y(_13927_));
 sky130_fd_sc_hd__inv_2 _23794_ (.A(_13927_),
    .Y(_13929_));
 sky130_fd_sc_hd__nand2_1 _23795_ (.A(_13907_),
    .B(_13929_),
    .Y(_13930_));
 sky130_fd_sc_hd__inv_2 _23796_ (.A(_13923_),
    .Y(_13931_));
 sky130_fd_sc_hd__a21boi_2 _23797_ (.A1(_13915_),
    .A2(_13931_),
    .B1_N(_13916_),
    .Y(_13932_));
 sky130_fd_sc_hd__nand2_1 _23798_ (.A(_13930_),
    .B(_13932_),
    .Y(_13933_));
 sky130_fd_sc_hd__nand2_1 _23799_ (.A(_13444_),
    .B(_13450_),
    .Y(_13934_));
 sky130_fd_sc_hd__inv_2 _23800_ (.A(_13306_),
    .Y(_13935_));
 sky130_fd_sc_hd__nand2_1 _23801_ (.A(_13934_),
    .B(_13935_),
    .Y(_13936_));
 sky130_fd_sc_hd__inv_2 _23802_ (.A(_13284_),
    .Y(_13937_));
 sky130_fd_sc_hd__nand2_1 _23803_ (.A(_13936_),
    .B(_13937_),
    .Y(_13938_));
 sky130_fd_sc_hd__nand3_1 _23804_ (.A(_13934_),
    .B(_13935_),
    .C(_13284_),
    .Y(_13940_));
 sky130_fd_sc_hd__nand2_1 _23805_ (.A(_13938_),
    .B(_13940_),
    .Y(_13941_));
 sky130_fd_sc_hd__nand2_1 _23806_ (.A(_13941_),
    .B(_12149_),
    .Y(_13942_));
 sky130_fd_sc_hd__nand3_1 _23807_ (.A(_13938_),
    .B(_13940_),
    .C(_12147_),
    .Y(_13943_));
 sky130_fd_sc_hd__nand2_1 _23808_ (.A(_13942_),
    .B(_13943_),
    .Y(_13944_));
 sky130_fd_sc_hd__inv_2 _23809_ (.A(_13944_),
    .Y(_13945_));
 sky130_fd_sc_hd__nand2_1 _23810_ (.A(_13933_),
    .B(_13945_),
    .Y(_13946_));
 sky130_fd_sc_hd__nand3_1 _23811_ (.A(_13930_),
    .B(_13944_),
    .C(_13932_),
    .Y(_13947_));
 sky130_fd_sc_hd__nand3_1 _23812_ (.A(_13946_),
    .B(_13842_),
    .C(_13947_),
    .Y(_13948_));
 sky130_fd_sc_hd__or2_1 _23813_ (.A(_13941_),
    .B(_13842_),
    .X(_13949_));
 sky130_fd_sc_hd__nand2_1 _23814_ (.A(_13948_),
    .B(_13949_),
    .Y(_13951_));
 sky130_fd_sc_hd__nand2_1 _23815_ (.A(_13951_),
    .B(_11701_),
    .Y(_13952_));
 sky130_fd_sc_hd__nand3_1 _23816_ (.A(_13948_),
    .B(_11703_),
    .C(_13949_),
    .Y(_13953_));
 sky130_fd_sc_hd__nand2_1 _23817_ (.A(_13952_),
    .B(_13953_),
    .Y(_13954_));
 sky130_fd_sc_hd__nand2_1 _23818_ (.A(_13907_),
    .B(_13926_),
    .Y(_13955_));
 sky130_fd_sc_hd__nand2_1 _23819_ (.A(_13955_),
    .B(_13923_),
    .Y(_13956_));
 sky130_fd_sc_hd__nand2_1 _23820_ (.A(_13956_),
    .B(_13919_),
    .Y(_13957_));
 sky130_fd_sc_hd__nand3_1 _23821_ (.A(_13955_),
    .B(_13918_),
    .C(_13923_),
    .Y(_13958_));
 sky130_fd_sc_hd__nand2_1 _23822_ (.A(_13957_),
    .B(_13958_),
    .Y(_13959_));
 sky130_fd_sc_hd__nand2_1 _23823_ (.A(_13959_),
    .B(_13842_),
    .Y(_13960_));
 sky130_fd_sc_hd__nand2_2 _23824_ (.A(\div1i.quot[5] ),
    .B(_13914_),
    .Y(_13962_));
 sky130_fd_sc_hd__nand2_1 _23825_ (.A(_13960_),
    .B(_13962_),
    .Y(_13963_));
 sky130_fd_sc_hd__nand2_1 _23826_ (.A(_13963_),
    .B(_11715_),
    .Y(_13964_));
 sky130_fd_sc_hd__nand3_4 _23827_ (.A(_13960_),
    .B(_11717_),
    .C(_13962_),
    .Y(_13965_));
 sky130_fd_sc_hd__nand2_2 _23828_ (.A(_13964_),
    .B(_13965_),
    .Y(_13966_));
 sky130_fd_sc_hd__nor2_2 _23829_ (.A(_13954_),
    .B(_13966_),
    .Y(_13967_));
 sky130_fd_sc_hd__or2_1 _23830_ (.A(_13926_),
    .B(_13907_),
    .X(_13968_));
 sky130_fd_sc_hd__nand3_1 _23831_ (.A(_13968_),
    .B(_13842_),
    .C(_13955_),
    .Y(_13969_));
 sky130_fd_sc_hd__nand2_1 _23832_ (.A(net226),
    .B(_13922_),
    .Y(_13970_));
 sky130_fd_sc_hd__nand2_1 _23833_ (.A(_13969_),
    .B(_13970_),
    .Y(_13971_));
 sky130_fd_sc_hd__nand2_1 _23834_ (.A(_13971_),
    .B(_06149_),
    .Y(_13973_));
 sky130_fd_sc_hd__nand3_1 _23835_ (.A(_13969_),
    .B(_13304_),
    .C(_13970_),
    .Y(_13974_));
 sky130_fd_sc_hd__nand2_1 _23836_ (.A(_13973_),
    .B(_13974_),
    .Y(_13975_));
 sky130_fd_sc_hd__nand2_1 _23837_ (.A(_13843_),
    .B(_13805_),
    .Y(_13976_));
 sky130_fd_sc_hd__xor2_1 _23838_ (.A(_13903_),
    .B(_13976_),
    .X(_13977_));
 sky130_fd_sc_hd__nand2_1 _23839_ (.A(_13977_),
    .B(_13842_),
    .Y(_13978_));
 sky130_fd_sc_hd__nand2_1 _23840_ (.A(\div1i.quot[5] ),
    .B(_13896_),
    .Y(_13979_));
 sky130_fd_sc_hd__nand2_1 _23841_ (.A(_13978_),
    .B(_13979_),
    .Y(_13980_));
 sky130_fd_sc_hd__nand2_1 _23842_ (.A(_13980_),
    .B(_11185_),
    .Y(_13981_));
 sky130_fd_sc_hd__nand3_2 _23843_ (.A(_13978_),
    .B(_12187_),
    .C(_13979_),
    .Y(_13982_));
 sky130_fd_sc_hd__nand2_2 _23844_ (.A(_13981_),
    .B(_13982_),
    .Y(_13984_));
 sky130_fd_sc_hd__nor2_2 _23845_ (.A(_13975_),
    .B(_13984_),
    .Y(_13985_));
 sky130_fd_sc_hd__nand2_1 _23846_ (.A(_13967_),
    .B(_13985_),
    .Y(_13986_));
 sky130_fd_sc_hd__inv_2 _23847_ (.A(_13986_),
    .Y(_13987_));
 sky130_fd_sc_hd__nand2_2 _23848_ (.A(_13889_),
    .B(_13987_),
    .Y(_13988_));
 sky130_fd_sc_hd__o21ai_1 _23849_ (.A1(_13982_),
    .A2(_13975_),
    .B1(_13973_),
    .Y(_13989_));
 sky130_fd_sc_hd__o21ai_1 _23850_ (.A1(_13965_),
    .A2(_13954_),
    .B1(_13952_),
    .Y(_13990_));
 sky130_fd_sc_hd__a21oi_2 _23851_ (.A1(_13967_),
    .A2(_13989_),
    .B1(_13990_),
    .Y(_13991_));
 sky130_fd_sc_hd__nand2_4 _23852_ (.A(_13988_),
    .B(_13991_),
    .Y(_13992_));
 sky130_fd_sc_hd__nand2_1 _23853_ (.A(_13938_),
    .B(_13283_),
    .Y(_13993_));
 sky130_fd_sc_hd__inv_2 _23854_ (.A(_13272_),
    .Y(_13995_));
 sky130_fd_sc_hd__nand2_1 _23855_ (.A(_13993_),
    .B(_13995_),
    .Y(_13996_));
 sky130_fd_sc_hd__nand3_1 _23856_ (.A(_13938_),
    .B(_13272_),
    .C(_13283_),
    .Y(_13997_));
 sky130_fd_sc_hd__nand2_1 _23857_ (.A(_13996_),
    .B(_13997_),
    .Y(_13998_));
 sky130_fd_sc_hd__nand2_1 _23858_ (.A(_13998_),
    .B(_12894_),
    .Y(_13999_));
 sky130_fd_sc_hd__nand3_1 _23859_ (.A(_13996_),
    .B(_11754_),
    .C(_13997_),
    .Y(_14000_));
 sky130_fd_sc_hd__nand3_1 _23860_ (.A(_13999_),
    .B(_14000_),
    .C(_13945_),
    .Y(_14001_));
 sky130_fd_sc_hd__nor2_1 _23861_ (.A(_14001_),
    .B(_13927_),
    .Y(_14002_));
 sky130_fd_sc_hd__nand2_2 _23862_ (.A(_13907_),
    .B(_14002_),
    .Y(_14003_));
 sky130_fd_sc_hd__nor2_1 _23863_ (.A(_14001_),
    .B(_13932_),
    .Y(_14004_));
 sky130_fd_sc_hd__nand2_1 _23864_ (.A(_13999_),
    .B(_14000_),
    .Y(_14006_));
 sky130_fd_sc_hd__o21ai_1 _23865_ (.A1(_13943_),
    .A2(_14006_),
    .B1(_14000_),
    .Y(_14007_));
 sky130_fd_sc_hd__nor2_1 _23866_ (.A(_14004_),
    .B(_14007_),
    .Y(_14008_));
 sky130_fd_sc_hd__nand2_2 _23867_ (.A(_14003_),
    .B(_14008_),
    .Y(_14009_));
 sky130_fd_sc_hd__clkinvlp_2 _23868_ (.A(_13488_),
    .Y(_14010_));
 sky130_fd_sc_hd__inv_2 _23869_ (.A(_13498_),
    .Y(_14011_));
 sky130_fd_sc_hd__nand2_1 _23870_ (.A(_13452_),
    .B(_14011_),
    .Y(_14012_));
 sky130_fd_sc_hd__nand2_1 _23871_ (.A(_14012_),
    .B(_13497_),
    .Y(_14013_));
 sky130_fd_sc_hd__or2_1 _23872_ (.A(_14010_),
    .B(_14013_),
    .X(_14014_));
 sky130_fd_sc_hd__nand2_1 _23873_ (.A(_14013_),
    .B(_14010_),
    .Y(_14015_));
 sky130_fd_sc_hd__nand2_1 _23874_ (.A(_14014_),
    .B(_14015_),
    .Y(_14017_));
 sky130_fd_sc_hd__nand2_1 _23875_ (.A(_14017_),
    .B(_12914_),
    .Y(_14018_));
 sky130_fd_sc_hd__nand3_1 _23876_ (.A(_14014_),
    .B(_11774_),
    .C(_14015_),
    .Y(_14019_));
 sky130_fd_sc_hd__nand2_1 _23877_ (.A(_14018_),
    .B(_14019_),
    .Y(_14020_));
 sky130_fd_sc_hd__or2_1 _23878_ (.A(_14011_),
    .B(_13452_),
    .X(_14021_));
 sky130_fd_sc_hd__nand2_1 _23879_ (.A(_14021_),
    .B(_14012_),
    .Y(_14022_));
 sky130_fd_sc_hd__inv_2 _23880_ (.A(_14022_),
    .Y(_14023_));
 sky130_fd_sc_hd__nand2_1 _23881_ (.A(_14023_),
    .B(_11199_),
    .Y(_14024_));
 sky130_fd_sc_hd__nand2_1 _23882_ (.A(_14022_),
    .B(_13461_),
    .Y(_14025_));
 sky130_fd_sc_hd__nand2_1 _23883_ (.A(_14024_),
    .B(_14025_),
    .Y(_14026_));
 sky130_fd_sc_hd__inv_2 _23884_ (.A(_14026_),
    .Y(_14028_));
 sky130_fd_sc_hd__nand2b_1 _23885_ (.A_N(_14020_),
    .B(_14028_),
    .Y(_14029_));
 sky130_fd_sc_hd__inv_2 _23886_ (.A(_14029_),
    .Y(_14030_));
 sky130_fd_sc_hd__nand2_1 _23887_ (.A(_14009_),
    .B(_14030_),
    .Y(_14031_));
 sky130_fd_sc_hd__inv_2 _23888_ (.A(_14024_),
    .Y(_14032_));
 sky130_fd_sc_hd__a21boi_1 _23889_ (.A1(_14018_),
    .A2(_14032_),
    .B1_N(_14019_),
    .Y(_14033_));
 sky130_fd_sc_hd__nand2_1 _23890_ (.A(_14031_),
    .B(_14033_),
    .Y(_14034_));
 sky130_fd_sc_hd__inv_2 _23891_ (.A(_13546_),
    .Y(_14035_));
 sky130_fd_sc_hd__nand2_1 _23892_ (.A(_13505_),
    .B(_14035_),
    .Y(_14036_));
 sky130_fd_sc_hd__nand3_1 _23893_ (.A(_13501_),
    .B(_13504_),
    .C(_13546_),
    .Y(_14037_));
 sky130_fd_sc_hd__nand2_1 _23894_ (.A(_14036_),
    .B(_14037_),
    .Y(_14039_));
 sky130_fd_sc_hd__inv_2 _23895_ (.A(_14039_),
    .Y(_14040_));
 sky130_fd_sc_hd__nand2_1 _23896_ (.A(_14040_),
    .B(_11797_),
    .Y(_14041_));
 sky130_fd_sc_hd__nand2_1 _23897_ (.A(_14039_),
    .B(_12939_),
    .Y(_14042_));
 sky130_fd_sc_hd__nand2_1 _23898_ (.A(_14041_),
    .B(_14042_),
    .Y(_14043_));
 sky130_fd_sc_hd__inv_2 _23899_ (.A(_14043_),
    .Y(_14044_));
 sky130_fd_sc_hd__nand2_1 _23900_ (.A(_14034_),
    .B(_14044_),
    .Y(_14045_));
 sky130_fd_sc_hd__buf_6 _23901_ (.A(_13842_),
    .X(_14046_));
 sky130_fd_sc_hd__nand3_1 _23902_ (.A(_14031_),
    .B(_14043_),
    .C(_14033_),
    .Y(_14047_));
 sky130_fd_sc_hd__nand3_1 _23903_ (.A(_14045_),
    .B(_14046_),
    .C(_14047_),
    .Y(_14048_));
 sky130_fd_sc_hd__nand2_1 _23904_ (.A(\div1i.quot[5] ),
    .B(_14040_),
    .Y(_14050_));
 sky130_fd_sc_hd__nand2_1 _23905_ (.A(_14048_),
    .B(_14050_),
    .Y(_14051_));
 sky130_fd_sc_hd__nand2_1 _23906_ (.A(_14051_),
    .B(_11808_),
    .Y(_14052_));
 sky130_fd_sc_hd__nand3_1 _23907_ (.A(_14048_),
    .B(_11811_),
    .C(_14050_),
    .Y(_14053_));
 sky130_fd_sc_hd__nand2_1 _23908_ (.A(_14052_),
    .B(_14053_),
    .Y(_14054_));
 sky130_fd_sc_hd__nand2_1 _23909_ (.A(_14009_),
    .B(_14028_),
    .Y(_14055_));
 sky130_fd_sc_hd__nand2_1 _23910_ (.A(_14055_),
    .B(_14024_),
    .Y(_14056_));
 sky130_fd_sc_hd__xor2_1 _23911_ (.A(_14020_),
    .B(_14056_),
    .X(_14057_));
 sky130_fd_sc_hd__nand2_1 _23912_ (.A(_14057_),
    .B(_14046_),
    .Y(_14058_));
 sky130_fd_sc_hd__nand2_1 _23913_ (.A(\div1i.quot[5] ),
    .B(_14017_),
    .Y(_14059_));
 sky130_fd_sc_hd__nand2_1 _23914_ (.A(_14058_),
    .B(_14059_),
    .Y(_14061_));
 sky130_fd_sc_hd__nand2_1 _23915_ (.A(_14061_),
    .B(_13537_),
    .Y(_14062_));
 sky130_fd_sc_hd__nand3_2 _23916_ (.A(_14058_),
    .B(_07400_),
    .C(_14059_),
    .Y(_14063_));
 sky130_fd_sc_hd__nand2_1 _23917_ (.A(_14062_),
    .B(_14063_),
    .Y(_14064_));
 sky130_fd_sc_hd__nor2_1 _23918_ (.A(_14054_),
    .B(_14064_),
    .Y(_14065_));
 sky130_fd_sc_hd__nand3_1 _23919_ (.A(_14003_),
    .B(_14008_),
    .C(_14026_),
    .Y(_14066_));
 sky130_fd_sc_hd__nand3_1 _23920_ (.A(_14055_),
    .B(_13842_),
    .C(_14066_),
    .Y(_14067_));
 sky130_fd_sc_hd__nand2_1 _23921_ (.A(net226),
    .B(_14023_),
    .Y(_14068_));
 sky130_fd_sc_hd__nand2_1 _23922_ (.A(_14067_),
    .B(_14068_),
    .Y(_14069_));
 sky130_fd_sc_hd__or2_1 _23923_ (.A(_13502_),
    .B(_14069_),
    .X(_14070_));
 sky130_fd_sc_hd__nand2_1 _23924_ (.A(_14069_),
    .B(_13502_),
    .Y(_14072_));
 sky130_fd_sc_hd__nand2_2 _23925_ (.A(_14070_),
    .B(_14072_),
    .Y(_14073_));
 sky130_fd_sc_hd__nand2_1 _23926_ (.A(_13946_),
    .B(_13943_),
    .Y(_14074_));
 sky130_fd_sc_hd__xor2_1 _23927_ (.A(_14006_),
    .B(_14074_),
    .X(_14075_));
 sky130_fd_sc_hd__nand2_1 _23928_ (.A(_14075_),
    .B(_14046_),
    .Y(_14076_));
 sky130_fd_sc_hd__nand2_1 _23929_ (.A(\div1i.quot[5] ),
    .B(_13998_),
    .Y(_14077_));
 sky130_fd_sc_hd__nand2_1 _23930_ (.A(_14076_),
    .B(_14077_),
    .Y(_14078_));
 sky130_fd_sc_hd__nand2_1 _23931_ (.A(_14078_),
    .B(_11838_),
    .Y(_14079_));
 sky130_fd_sc_hd__nand3_2 _23932_ (.A(_14076_),
    .B(_11840_),
    .C(_14077_),
    .Y(_14080_));
 sky130_fd_sc_hd__nand3b_1 _23933_ (.A_N(_14073_),
    .B(_14079_),
    .C(_14080_),
    .Y(_14081_));
 sky130_fd_sc_hd__inv_4 _23934_ (.A(_14081_),
    .Y(_14083_));
 sky130_fd_sc_hd__nand3_4 _23935_ (.A(_13992_),
    .B(_14065_),
    .C(_14083_),
    .Y(_14084_));
 sky130_fd_sc_hd__inv_2 _23936_ (.A(_14072_),
    .Y(_14085_));
 sky130_fd_sc_hd__o21bai_2 _23937_ (.A1(_14073_),
    .A2(_14080_),
    .B1_N(_14085_),
    .Y(_14086_));
 sky130_fd_sc_hd__o21ai_1 _23938_ (.A1(_14054_),
    .A2(_14063_),
    .B1(_14052_),
    .Y(_14087_));
 sky130_fd_sc_hd__a21oi_2 _23939_ (.A1(_14065_),
    .A2(_14086_),
    .B1(_14087_),
    .Y(_14088_));
 sky130_fd_sc_hd__nand2_2 _23940_ (.A(_14084_),
    .B(_14088_),
    .Y(_14089_));
 sky130_fd_sc_hd__nand2_1 _23941_ (.A(_14036_),
    .B(_13543_),
    .Y(_14090_));
 sky130_fd_sc_hd__inv_2 _23942_ (.A(_13536_),
    .Y(_14091_));
 sky130_fd_sc_hd__nand2_1 _23943_ (.A(_14090_),
    .B(_14091_),
    .Y(_14092_));
 sky130_fd_sc_hd__nand3_1 _23944_ (.A(_14036_),
    .B(_13536_),
    .C(_13543_),
    .Y(_14094_));
 sky130_fd_sc_hd__nand2_1 _23945_ (.A(_14092_),
    .B(_14094_),
    .Y(_14095_));
 sky130_fd_sc_hd__nand2_1 _23946_ (.A(_14095_),
    .B(_12992_),
    .Y(_14096_));
 sky130_fd_sc_hd__nand3_1 _23947_ (.A(_14092_),
    .B(_11858_),
    .C(_14094_),
    .Y(_14097_));
 sky130_fd_sc_hd__nand3_1 _23948_ (.A(_14044_),
    .B(_14096_),
    .C(_14097_),
    .Y(_14098_));
 sky130_fd_sc_hd__inv_2 _23949_ (.A(_14098_),
    .Y(_14099_));
 sky130_fd_sc_hd__nand3_2 _23950_ (.A(_14009_),
    .B(_14030_),
    .C(_14099_),
    .Y(_14100_));
 sky130_fd_sc_hd__inv_2 _23951_ (.A(_14096_),
    .Y(_14101_));
 sky130_fd_sc_hd__o21ai_1 _23952_ (.A1(_14041_),
    .A2(_14101_),
    .B1(_14097_),
    .Y(_14102_));
 sky130_fd_sc_hd__nor2_1 _23953_ (.A(_14033_),
    .B(_14098_),
    .Y(_14103_));
 sky130_fd_sc_hd__nor2_1 _23954_ (.A(_14102_),
    .B(_14103_),
    .Y(_14105_));
 sky130_fd_sc_hd__nand2_1 _23955_ (.A(_14100_),
    .B(_14105_),
    .Y(_14106_));
 sky130_fd_sc_hd__inv_2 _23956_ (.A(_13551_),
    .Y(_14107_));
 sky130_fd_sc_hd__nand2_1 _23957_ (.A(_13596_),
    .B(_13597_),
    .Y(_14108_));
 sky130_fd_sc_hd__nand2_1 _23958_ (.A(_14107_),
    .B(_14108_),
    .Y(_14109_));
 sky130_fd_sc_hd__inv_2 _23959_ (.A(_14108_),
    .Y(_14110_));
 sky130_fd_sc_hd__nand2_1 _23960_ (.A(_13551_),
    .B(_14110_),
    .Y(_14111_));
 sky130_fd_sc_hd__nand2_1 _23961_ (.A(_14109_),
    .B(_14111_),
    .Y(_14112_));
 sky130_fd_sc_hd__buf_6 _23962_ (.A(_10749_),
    .X(_14113_));
 sky130_fd_sc_hd__nand2_1 _23963_ (.A(_14112_),
    .B(_14113_),
    .Y(_14114_));
 sky130_fd_sc_hd__nand3_2 _23964_ (.A(_14109_),
    .B(_08554_),
    .C(_14111_),
    .Y(_14116_));
 sky130_fd_sc_hd__nand2_1 _23965_ (.A(_14114_),
    .B(_14116_),
    .Y(_14117_));
 sky130_fd_sc_hd__inv_2 _23966_ (.A(_14117_),
    .Y(_14118_));
 sky130_fd_sc_hd__nand2_1 _23967_ (.A(_14106_),
    .B(_14118_),
    .Y(_14119_));
 sky130_fd_sc_hd__nand2_1 _23968_ (.A(_14119_),
    .B(_14116_),
    .Y(_14120_));
 sky130_fd_sc_hd__nand2_1 _23969_ (.A(_14111_),
    .B(_13597_),
    .Y(_14121_));
 sky130_fd_sc_hd__xor2_2 _23970_ (.A(_13587_),
    .B(_14121_),
    .X(_14122_));
 sky130_fd_sc_hd__inv_2 _23971_ (.A(_14122_),
    .Y(_14123_));
 sky130_fd_sc_hd__nand2_1 _23972_ (.A(_14123_),
    .B(_12495_),
    .Y(_14124_));
 sky130_fd_sc_hd__nand2_1 _23973_ (.A(_14122_),
    .B(_13042_),
    .Y(_14125_));
 sky130_fd_sc_hd__nand2_1 _23974_ (.A(_14124_),
    .B(_14125_),
    .Y(_14127_));
 sky130_fd_sc_hd__inv_2 _23975_ (.A(_14127_),
    .Y(_14128_));
 sky130_fd_sc_hd__nand2_1 _23976_ (.A(_14120_),
    .B(_14128_),
    .Y(_14129_));
 sky130_fd_sc_hd__nand3_1 _23977_ (.A(_14119_),
    .B(_14127_),
    .C(_14116_),
    .Y(_14130_));
 sky130_fd_sc_hd__nand2_1 _23978_ (.A(_14129_),
    .B(_14130_),
    .Y(_14131_));
 sky130_fd_sc_hd__nand2_1 _23979_ (.A(_14131_),
    .B(_14046_),
    .Y(_14132_));
 sky130_fd_sc_hd__nand2_1 _23980_ (.A(_14122_),
    .B(\div1i.quot[5] ),
    .Y(_14133_));
 sky130_fd_sc_hd__nand2_1 _23981_ (.A(_14132_),
    .B(_14133_),
    .Y(_14134_));
 sky130_fd_sc_hd__nand2_1 _23982_ (.A(_14134_),
    .B(_12506_),
    .Y(_14135_));
 sky130_fd_sc_hd__nand3_1 _23983_ (.A(_14132_),
    .B(_11376_),
    .C(_14133_),
    .Y(_14136_));
 sky130_fd_sc_hd__nand2_1 _23984_ (.A(_14135_),
    .B(_14136_),
    .Y(_14138_));
 sky130_fd_sc_hd__inv_2 _23985_ (.A(_14138_),
    .Y(_14139_));
 sky130_fd_sc_hd__nand3_1 _23986_ (.A(_14124_),
    .B(_14125_),
    .C(_14118_),
    .Y(_14140_));
 sky130_fd_sc_hd__inv_2 _23987_ (.A(_14140_),
    .Y(_14141_));
 sky130_fd_sc_hd__nand2_1 _23988_ (.A(_14141_),
    .B(_14106_),
    .Y(_14142_));
 sky130_fd_sc_hd__inv_2 _23989_ (.A(_14125_),
    .Y(_14143_));
 sky130_fd_sc_hd__o21a_1 _23990_ (.A1(_14116_),
    .A2(_14143_),
    .B1(_14124_),
    .X(_14144_));
 sky130_fd_sc_hd__nand2_1 _23991_ (.A(_14142_),
    .B(_14144_),
    .Y(_14145_));
 sky130_fd_sc_hd__o21bai_1 _23992_ (.A1(_13598_),
    .A2(_14107_),
    .B1_N(_13650_),
    .Y(_14146_));
 sky130_fd_sc_hd__or2_1 _23993_ (.A(_13619_),
    .B(_14146_),
    .X(_14147_));
 sky130_fd_sc_hd__nand2_1 _23994_ (.A(_14146_),
    .B(_13619_),
    .Y(_14149_));
 sky130_fd_sc_hd__nand2_1 _23995_ (.A(_14147_),
    .B(_14149_),
    .Y(_14150_));
 sky130_fd_sc_hd__inv_2 _23996_ (.A(_14150_),
    .Y(_14151_));
 sky130_fd_sc_hd__nand2_1 _23997_ (.A(_14151_),
    .B(_11935_),
    .Y(_14152_));
 sky130_fd_sc_hd__nand2_1 _23998_ (.A(_14150_),
    .B(_13633_),
    .Y(_14153_));
 sky130_fd_sc_hd__nand2_1 _23999_ (.A(_14152_),
    .B(_14153_),
    .Y(_14154_));
 sky130_fd_sc_hd__inv_2 _24000_ (.A(_14154_),
    .Y(_14155_));
 sky130_fd_sc_hd__nand2_1 _24001_ (.A(_14145_),
    .B(_14155_),
    .Y(_14156_));
 sky130_fd_sc_hd__nand3_1 _24002_ (.A(_14142_),
    .B(_14144_),
    .C(_14154_),
    .Y(_14157_));
 sky130_fd_sc_hd__nand3_1 _24003_ (.A(_14156_),
    .B(_14157_),
    .C(_14046_),
    .Y(_14158_));
 sky130_fd_sc_hd__nand2_1 _24004_ (.A(_14151_),
    .B(\div1i.quot[5] ),
    .Y(_14160_));
 sky130_fd_sc_hd__nand2_1 _24005_ (.A(_14158_),
    .B(_14160_),
    .Y(_14161_));
 sky130_fd_sc_hd__nand2_1 _24006_ (.A(_14161_),
    .B(_11946_),
    .Y(_14162_));
 sky130_fd_sc_hd__nand3_1 _24007_ (.A(_14158_),
    .B(_11948_),
    .C(_14160_),
    .Y(_14163_));
 sky130_fd_sc_hd__nand2_2 _24008_ (.A(_14162_),
    .B(_14163_),
    .Y(_14164_));
 sky130_fd_sc_hd__inv_2 _24009_ (.A(_14164_),
    .Y(_14165_));
 sky130_fd_sc_hd__nand2_1 _24010_ (.A(_14139_),
    .B(_14165_),
    .Y(_14166_));
 sky130_fd_sc_hd__nand3_1 _24011_ (.A(_14100_),
    .B(_14105_),
    .C(_14117_),
    .Y(_14167_));
 sky130_fd_sc_hd__nand3_1 _24012_ (.A(_14119_),
    .B(_14167_),
    .C(_14046_),
    .Y(_14168_));
 sky130_fd_sc_hd__or2_1 _24013_ (.A(_14112_),
    .B(_14046_),
    .X(_14169_));
 sky130_fd_sc_hd__nand2_1 _24014_ (.A(_14168_),
    .B(_14169_),
    .Y(_14171_));
 sky130_fd_sc_hd__or2_1 _24015_ (.A(_13022_),
    .B(_14171_),
    .X(_14172_));
 sky130_fd_sc_hd__nand2_1 _24016_ (.A(_14171_),
    .B(_13022_),
    .Y(_14173_));
 sky130_fd_sc_hd__nand2_2 _24017_ (.A(_14172_),
    .B(_14173_),
    .Y(_14174_));
 sky130_fd_sc_hd__nand2_1 _24018_ (.A(_14096_),
    .B(_14097_),
    .Y(_14175_));
 sky130_fd_sc_hd__nand2_1 _24019_ (.A(_14045_),
    .B(_14041_),
    .Y(_14176_));
 sky130_fd_sc_hd__xor2_1 _24020_ (.A(_14175_),
    .B(_14176_),
    .X(_14177_));
 sky130_fd_sc_hd__nand2_1 _24021_ (.A(_14177_),
    .B(_14046_),
    .Y(_14178_));
 sky130_fd_sc_hd__nand2_1 _24022_ (.A(\div1i.quot[5] ),
    .B(_14095_),
    .Y(_14179_));
 sky130_fd_sc_hd__nand3_2 _24023_ (.A(_14178_),
    .B(_11899_),
    .C(_14179_),
    .Y(_14180_));
 sky130_fd_sc_hd__nand2_1 _24024_ (.A(_14178_),
    .B(_14179_),
    .Y(_14182_));
 sky130_fd_sc_hd__nand2_1 _24025_ (.A(_14182_),
    .B(_11896_),
    .Y(_14183_));
 sky130_fd_sc_hd__nand3b_1 _24026_ (.A_N(_14174_),
    .B(_14180_),
    .C(_14183_),
    .Y(_14184_));
 sky130_fd_sc_hd__nor2_1 _24027_ (.A(_14166_),
    .B(_14184_),
    .Y(_14185_));
 sky130_fd_sc_hd__nand2_4 _24028_ (.A(_14089_),
    .B(_14185_),
    .Y(_14186_));
 sky130_fd_sc_hd__o21ai_1 _24029_ (.A1(_14174_),
    .A2(_14180_),
    .B1(_14173_),
    .Y(_14187_));
 sky130_fd_sc_hd__nor2_1 _24030_ (.A(_14164_),
    .B(_14138_),
    .Y(_14188_));
 sky130_fd_sc_hd__inv_2 _24031_ (.A(_14163_),
    .Y(_14189_));
 sky130_fd_sc_hd__o21ai_1 _24032_ (.A1(_14136_),
    .A2(_14189_),
    .B1(_14162_),
    .Y(_14190_));
 sky130_fd_sc_hd__a21oi_2 _24033_ (.A1(_14187_),
    .A2(_14188_),
    .B1(_14190_),
    .Y(_14191_));
 sky130_fd_sc_hd__nand2_2 _24034_ (.A(_14191_),
    .B(_14186_),
    .Y(_14193_));
 sky130_fd_sc_hd__nand2_1 _24035_ (.A(_14149_),
    .B(_13617_),
    .Y(_14194_));
 sky130_fd_sc_hd__xor2_1 _24036_ (.A(_13645_),
    .B(_14194_),
    .X(_14195_));
 sky130_fd_sc_hd__nand3_1 _24037_ (.A(_14156_),
    .B(_14046_),
    .C(_14152_),
    .Y(_14196_));
 sky130_fd_sc_hd__xnor2_2 _24038_ (.A(_14195_),
    .B(_14196_),
    .Y(_14197_));
 sky130_fd_sc_hd__nand2_4 _24039_ (.A(_14193_),
    .B(_14197_),
    .Y(_14198_));
 sky130_fd_sc_hd__clkinvlp_2 _24040_ (.A(_14197_),
    .Y(_14199_));
 sky130_fd_sc_hd__nand3_4 _24041_ (.A(_14186_),
    .B(_14191_),
    .C(_14199_),
    .Y(_14200_));
 sky130_fd_sc_hd__nand2_8 _24042_ (.A(_14198_),
    .B(_14200_),
    .Y(_14201_));
 sky130_fd_sc_hd__buf_8 _24043_ (.A(_14201_),
    .X(_14202_));
 sky130_fd_sc_hd__buf_6 _24044_ (.A(net232),
    .X(\div1i.quot[4] ));
 sky130_fd_sc_hd__nand2_1 _24045_ (.A(_13794_),
    .B(_13881_),
    .Y(_14204_));
 sky130_fd_sc_hd__inv_2 _24046_ (.A(_13886_),
    .Y(_14205_));
 sky130_fd_sc_hd__nand2_1 _24047_ (.A(_14204_),
    .B(_14205_),
    .Y(_14206_));
 sky130_fd_sc_hd__inv_2 _24048_ (.A(_13861_),
    .Y(_14207_));
 sky130_fd_sc_hd__nand2_1 _24049_ (.A(_14206_),
    .B(_14207_),
    .Y(_14208_));
 sky130_fd_sc_hd__nand2_1 _24050_ (.A(_14208_),
    .B(_13860_),
    .Y(_14209_));
 sky130_fd_sc_hd__inv_2 _24051_ (.A(_13849_),
    .Y(_14210_));
 sky130_fd_sc_hd__nand2_1 _24052_ (.A(_14209_),
    .B(_14210_),
    .Y(_14211_));
 sky130_fd_sc_hd__nand3_1 _24053_ (.A(_14208_),
    .B(_13849_),
    .C(_13860_),
    .Y(_14212_));
 sky130_fd_sc_hd__nand2_1 _24054_ (.A(_14211_),
    .B(_14212_),
    .Y(_14214_));
 sky130_fd_sc_hd__nand2_2 _24055_ (.A(_14214_),
    .B(_11983_),
    .Y(_14215_));
 sky130_fd_sc_hd__nand3_1 _24056_ (.A(_14204_),
    .B(_13861_),
    .C(_14205_),
    .Y(_14216_));
 sky130_fd_sc_hd__nand3_2 _24057_ (.A(_14208_),
    .B(_11986_),
    .C(_14216_),
    .Y(_14217_));
 sky130_fd_sc_hd__inv_2 _24058_ (.A(_14217_),
    .Y(_14218_));
 sky130_fd_sc_hd__nand3_2 _24059_ (.A(_14211_),
    .B(_11990_),
    .C(_14212_),
    .Y(_14219_));
 sky130_fd_sc_hd__nand3_1 _24060_ (.A(_14215_),
    .B(_14218_),
    .C(_14219_),
    .Y(_14220_));
 sky130_fd_sc_hd__nand2_1 _24061_ (.A(_14220_),
    .B(_14219_),
    .Y(_14221_));
 sky130_fd_sc_hd__inv_2 _24062_ (.A(_13880_),
    .Y(_14222_));
 sky130_fd_sc_hd__nand2_1 _24063_ (.A(_13794_),
    .B(_14222_),
    .Y(_14223_));
 sky130_fd_sc_hd__nand2_1 _24064_ (.A(_14223_),
    .B(_13878_),
    .Y(_14225_));
 sky130_fd_sc_hd__inv_2 _24065_ (.A(_13870_),
    .Y(_14226_));
 sky130_fd_sc_hd__nand2_1 _24066_ (.A(_14225_),
    .B(_14226_),
    .Y(_14227_));
 sky130_fd_sc_hd__nand3_1 _24067_ (.A(_14223_),
    .B(_13870_),
    .C(_13878_),
    .Y(_14228_));
 sky130_fd_sc_hd__nand2_1 _24068_ (.A(_14227_),
    .B(_14228_),
    .Y(_14229_));
 sky130_fd_sc_hd__nand2_1 _24069_ (.A(_14229_),
    .B(_12002_),
    .Y(_14230_));
 sky130_fd_sc_hd__or2_1 _24070_ (.A(_14222_),
    .B(_13794_),
    .X(_14231_));
 sky130_fd_sc_hd__nand2_1 _24071_ (.A(_14231_),
    .B(_14223_),
    .Y(_14232_));
 sky130_fd_sc_hd__inv_2 _24072_ (.A(_14232_),
    .Y(_14233_));
 sky130_fd_sc_hd__nand2_1 _24073_ (.A(_14233_),
    .B(_12008_),
    .Y(_14234_));
 sky130_fd_sc_hd__inv_2 _24074_ (.A(_14234_),
    .Y(_14236_));
 sky130_fd_sc_hd__inv_2 _24075_ (.A(_14229_),
    .Y(_14237_));
 sky130_fd_sc_hd__nand2_1 _24076_ (.A(_14237_),
    .B(_12012_),
    .Y(_14238_));
 sky130_fd_sc_hd__inv_2 _24077_ (.A(_14238_),
    .Y(_14239_));
 sky130_fd_sc_hd__a21oi_2 _24078_ (.A1(_14230_),
    .A2(_14236_),
    .B1(_14239_),
    .Y(_14240_));
 sky130_fd_sc_hd__nand2_1 _24079_ (.A(_14208_),
    .B(_14216_),
    .Y(_14241_));
 sky130_fd_sc_hd__nand2_1 _24080_ (.A(_14241_),
    .B(_12017_),
    .Y(_14242_));
 sky130_fd_sc_hd__nand2_1 _24081_ (.A(_14242_),
    .B(_14217_),
    .Y(_14243_));
 sky130_fd_sc_hd__inv_2 _24082_ (.A(_14243_),
    .Y(_14244_));
 sky130_fd_sc_hd__nand3_2 _24083_ (.A(_14215_),
    .B(_14244_),
    .C(_14219_),
    .Y(_14245_));
 sky130_fd_sc_hd__nor2_1 _24084_ (.A(_14240_),
    .B(_14245_),
    .Y(_14247_));
 sky130_fd_sc_hd__nor2_1 _24085_ (.A(_14221_),
    .B(_14247_),
    .Y(_14248_));
 sky130_fd_sc_hd__inv_2 _24086_ (.A(_14245_),
    .Y(_14249_));
 sky130_fd_sc_hd__nand2_1 _24087_ (.A(_13689_),
    .B(_13692_),
    .Y(_14250_));
 sky130_fd_sc_hd__nand2_1 _24088_ (.A(_14250_),
    .B(_13693_),
    .Y(_14251_));
 sky130_fd_sc_hd__nand2_1 _24089_ (.A(_14251_),
    .B(_13695_),
    .Y(_14252_));
 sky130_fd_sc_hd__nand2_1 _24090_ (.A(_14252_),
    .B(_12030_),
    .Y(_14253_));
 sky130_fd_sc_hd__o21ai_1 _24091_ (.A1(_12032_),
    .A2(\div1i.quot[5] ),
    .B1(_12033_),
    .Y(_14254_));
 sky130_fd_sc_hd__nand3_1 _24092_ (.A(_14251_),
    .B(_12035_),
    .C(_13695_),
    .Y(_14255_));
 sky130_fd_sc_hd__inv_2 _24093_ (.A(_14255_),
    .Y(_14256_));
 sky130_fd_sc_hd__a21o_1 _24094_ (.A1(_14253_),
    .A2(_14254_),
    .B1(_14256_),
    .X(_14258_));
 sky130_fd_sc_hd__nand2_1 _24095_ (.A(_13696_),
    .B(_13680_),
    .Y(_14259_));
 sky130_fd_sc_hd__nand2_1 _24096_ (.A(_13695_),
    .B(_13689_),
    .Y(_14260_));
 sky130_fd_sc_hd__xor2_1 _24097_ (.A(_14259_),
    .B(_14260_),
    .X(_14261_));
 sky130_fd_sc_hd__nand2_1 _24098_ (.A(_14261_),
    .B(_12043_),
    .Y(_14262_));
 sky130_fd_sc_hd__nand2_1 _24099_ (.A(_14258_),
    .B(_14262_),
    .Y(_14263_));
 sky130_fd_sc_hd__inv_2 _24100_ (.A(_14261_),
    .Y(_14264_));
 sky130_fd_sc_hd__nand2_1 _24101_ (.A(_14264_),
    .B(_12047_),
    .Y(_14265_));
 sky130_fd_sc_hd__nand2_1 _24102_ (.A(_14263_),
    .B(_14265_),
    .Y(_14266_));
 sky130_fd_sc_hd__nand2_1 _24103_ (.A(_13691_),
    .B(_13695_),
    .Y(_14267_));
 sky130_fd_sc_hd__nand2_1 _24104_ (.A(_14267_),
    .B(_13696_),
    .Y(_14269_));
 sky130_fd_sc_hd__nand2_1 _24105_ (.A(_14269_),
    .B(_13782_),
    .Y(_14270_));
 sky130_fd_sc_hd__nand3_1 _24106_ (.A(_14267_),
    .B(_13696_),
    .C(_13783_),
    .Y(_14271_));
 sky130_fd_sc_hd__nand2_1 _24107_ (.A(_14270_),
    .B(_14271_),
    .Y(_14272_));
 sky130_fd_sc_hd__nand2_1 _24108_ (.A(_14272_),
    .B(_12056_),
    .Y(_14273_));
 sky130_fd_sc_hd__nand3_1 _24109_ (.A(_14270_),
    .B(_12058_),
    .C(_14271_),
    .Y(_14274_));
 sky130_fd_sc_hd__nand2_1 _24110_ (.A(_14273_),
    .B(_14274_),
    .Y(_14275_));
 sky130_fd_sc_hd__inv_2 _24111_ (.A(_14275_),
    .Y(_14276_));
 sky130_fd_sc_hd__nand2_1 _24112_ (.A(_14266_),
    .B(_14276_),
    .Y(_14277_));
 sky130_fd_sc_hd__nand2_2 _24113_ (.A(_14277_),
    .B(_14274_),
    .Y(_14278_));
 sky130_fd_sc_hd__nand2_1 _24114_ (.A(_14271_),
    .B(_13780_),
    .Y(_14280_));
 sky130_fd_sc_hd__xor2_2 _24115_ (.A(_13772_),
    .B(_14280_),
    .X(_14281_));
 sky130_fd_sc_hd__nand2_1 _24116_ (.A(_14281_),
    .B(_13182_),
    .Y(_14282_));
 sky130_fd_sc_hd__nand2_1 _24117_ (.A(_14278_),
    .B(_14282_),
    .Y(_14283_));
 sky130_fd_sc_hd__or2_1 _24118_ (.A(_13182_),
    .B(_14281_),
    .X(_14284_));
 sky130_fd_sc_hd__nand2_1 _24119_ (.A(_14283_),
    .B(_14284_),
    .Y(_14285_));
 sky130_fd_sc_hd__nor2_1 _24120_ (.A(_13772_),
    .B(_13782_),
    .Y(_14286_));
 sky130_fd_sc_hd__nand3_1 _24121_ (.A(_14267_),
    .B(_14286_),
    .C(_13696_),
    .Y(_14287_));
 sky130_fd_sc_hd__inv_2 _24122_ (.A(_13789_),
    .Y(_14288_));
 sky130_fd_sc_hd__nand2_1 _24123_ (.A(_14287_),
    .B(_14288_),
    .Y(_14289_));
 sky130_fd_sc_hd__nand2_1 _24124_ (.A(_14289_),
    .B(_13760_),
    .Y(_00037_));
 sky130_fd_sc_hd__nand2_1 _24125_ (.A(_00037_),
    .B(_13757_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _24126_ (.A(_00038_),
    .B(_13750_),
    .Y(_00039_));
 sky130_fd_sc_hd__nand3_1 _24127_ (.A(_00037_),
    .B(_13749_),
    .C(_13757_),
    .Y(_00040_));
 sky130_fd_sc_hd__nand2_1 _24128_ (.A(_00039_),
    .B(_00040_),
    .Y(_00041_));
 sky130_fd_sc_hd__nand2_1 _24129_ (.A(_00041_),
    .B(_13197_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand3_1 _24130_ (.A(_14287_),
    .B(_13759_),
    .C(_14288_),
    .Y(_00043_));
 sky130_fd_sc_hd__nand2_1 _24131_ (.A(_00037_),
    .B(_00043_),
    .Y(_00044_));
 sky130_fd_sc_hd__nand2_1 _24132_ (.A(_00044_),
    .B(_12085_),
    .Y(_00045_));
 sky130_fd_sc_hd__nand3_2 _24133_ (.A(_00037_),
    .B(_12087_),
    .C(_00043_),
    .Y(_00046_));
 sky130_fd_sc_hd__nand2_1 _24134_ (.A(_00045_),
    .B(_00046_),
    .Y(_00048_));
 sky130_fd_sc_hd__inv_2 _24135_ (.A(_00048_),
    .Y(_00049_));
 sky130_fd_sc_hd__nand3_1 _24136_ (.A(_00039_),
    .B(_10939_),
    .C(_00040_),
    .Y(_00050_));
 sky130_fd_sc_hd__nand3_1 _24137_ (.A(_00042_),
    .B(_00049_),
    .C(_00050_),
    .Y(_00051_));
 sky130_fd_sc_hd__inv_2 _24138_ (.A(_00051_),
    .Y(_00052_));
 sky130_fd_sc_hd__nand2_1 _24139_ (.A(_14285_),
    .B(_00052_),
    .Y(_00053_));
 sky130_fd_sc_hd__inv_2 _24140_ (.A(_00046_),
    .Y(_00054_));
 sky130_fd_sc_hd__a21boi_1 _24141_ (.A1(_00042_),
    .A2(_00054_),
    .B1_N(_00050_),
    .Y(_00055_));
 sky130_fd_sc_hd__nand2_1 _24142_ (.A(_00053_),
    .B(_00055_),
    .Y(_00056_));
 sky130_fd_sc_hd__nand2_1 _24143_ (.A(_14238_),
    .B(_14230_),
    .Y(_00057_));
 sky130_fd_sc_hd__inv_2 _24144_ (.A(_00057_),
    .Y(_00059_));
 sky130_fd_sc_hd__nand2_1 _24145_ (.A(_14232_),
    .B(_12101_),
    .Y(_00060_));
 sky130_fd_sc_hd__nand2_1 _24146_ (.A(_14234_),
    .B(_00060_),
    .Y(_00061_));
 sky130_fd_sc_hd__inv_2 _24147_ (.A(_00061_),
    .Y(_00062_));
 sky130_fd_sc_hd__nand2_1 _24148_ (.A(_00059_),
    .B(_00062_),
    .Y(_00063_));
 sky130_fd_sc_hd__inv_2 _24149_ (.A(_00063_),
    .Y(_00064_));
 sky130_fd_sc_hd__nand3_1 _24150_ (.A(_14249_),
    .B(_00056_),
    .C(_00064_),
    .Y(_00065_));
 sky130_fd_sc_hd__nand2_2 _24151_ (.A(_14248_),
    .B(_00065_),
    .Y(_00066_));
 sky130_fd_sc_hd__inv_2 _24152_ (.A(_13975_),
    .Y(_00067_));
 sky130_fd_sc_hd__inv_2 _24153_ (.A(_13984_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_1 _24154_ (.A(_13889_),
    .B(_00068_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_1 _24155_ (.A(_00070_),
    .B(_13982_),
    .Y(_00071_));
 sky130_fd_sc_hd__or2_1 _24156_ (.A(_00067_),
    .B(_00071_),
    .X(_00072_));
 sky130_fd_sc_hd__nand2_1 _24157_ (.A(_00071_),
    .B(_00067_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_1 _24158_ (.A(_00072_),
    .B(_00073_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_1 _24159_ (.A(_00074_),
    .B(_12118_),
    .Y(_00075_));
 sky130_fd_sc_hd__nand3_1 _24160_ (.A(_00072_),
    .B(_12120_),
    .C(_00073_),
    .Y(_00076_));
 sky130_fd_sc_hd__nand2_1 _24161_ (.A(_00075_),
    .B(_00076_),
    .Y(_00077_));
 sky130_fd_sc_hd__inv_2 _24162_ (.A(_00077_),
    .Y(_00078_));
 sky130_fd_sc_hd__or2_1 _24163_ (.A(_00068_),
    .B(_13889_),
    .X(_00079_));
 sky130_fd_sc_hd__nand2_1 _24164_ (.A(_00079_),
    .B(_00070_),
    .Y(_00081_));
 sky130_fd_sc_hd__inv_2 _24165_ (.A(_00081_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand2_1 _24166_ (.A(_00082_),
    .B(_11671_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_1 _24167_ (.A(_00081_),
    .B(_12817_),
    .Y(_00084_));
 sky130_fd_sc_hd__nand2_1 _24168_ (.A(_00083_),
    .B(_00084_),
    .Y(_00085_));
 sky130_fd_sc_hd__inv_2 _24169_ (.A(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_1 _24170_ (.A(_00078_),
    .B(_00086_),
    .Y(_00087_));
 sky130_fd_sc_hd__inv_2 _24171_ (.A(_00087_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_1 _24172_ (.A(_00066_),
    .B(_00088_),
    .Y(_00089_));
 sky130_fd_sc_hd__inv_2 _24173_ (.A(_00083_),
    .Y(_00090_));
 sky130_fd_sc_hd__a21boi_2 _24174_ (.A1(_00075_),
    .A2(_00090_),
    .B1_N(_00076_),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_1 _24175_ (.A(_00089_),
    .B(_00092_),
    .Y(_00093_));
 sky130_fd_sc_hd__nand2_1 _24176_ (.A(_13889_),
    .B(_13985_),
    .Y(_00094_));
 sky130_fd_sc_hd__inv_2 _24177_ (.A(_13989_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_1 _24178_ (.A(_00094_),
    .B(_00095_),
    .Y(_00096_));
 sky130_fd_sc_hd__inv_2 _24179_ (.A(_13966_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_1 _24180_ (.A(_00096_),
    .B(_00097_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand3_1 _24181_ (.A(_00094_),
    .B(_13966_),
    .C(_00095_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand2_1 _24182_ (.A(_00098_),
    .B(_00099_),
    .Y(_00100_));
 sky130_fd_sc_hd__inv_2 _24183_ (.A(_00100_),
    .Y(_00101_));
 sky130_fd_sc_hd__nand2_1 _24184_ (.A(_00101_),
    .B(_12147_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_1 _24185_ (.A(_00100_),
    .B(_12149_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_1 _24186_ (.A(_00103_),
    .B(_00104_),
    .Y(_00105_));
 sky130_fd_sc_hd__inv_2 _24187_ (.A(_00105_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_1 _24188_ (.A(_00093_),
    .B(_00106_),
    .Y(_00107_));
 sky130_fd_sc_hd__inv_6 _24189_ (.A(_14201_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand3_1 _24190_ (.A(_00089_),
    .B(_00105_),
    .C(_00092_),
    .Y(_00109_));
 sky130_fd_sc_hd__nand3_1 _24191_ (.A(_00107_),
    .B(_00108_),
    .C(_00109_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_1 _24192_ (.A(net232),
    .B(_00101_),
    .Y(_00111_));
 sky130_fd_sc_hd__nand2_1 _24193_ (.A(_00110_),
    .B(_00111_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_1 _24194_ (.A(_00112_),
    .B(_11701_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand3_1 _24195_ (.A(_00110_),
    .B(_11703_),
    .C(_00111_),
    .Y(_00115_));
 sky130_fd_sc_hd__nand2_1 _24196_ (.A(_00114_),
    .B(_00115_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_1 _24197_ (.A(_00066_),
    .B(_00086_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_1 _24198_ (.A(_00117_),
    .B(_00083_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_1 _24199_ (.A(_00118_),
    .B(_00078_),
    .Y(_00119_));
 sky130_fd_sc_hd__nand3_1 _24200_ (.A(_00117_),
    .B(_00077_),
    .C(_00083_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _24201_ (.A(_00119_),
    .B(_00120_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_1 _24202_ (.A(_00121_),
    .B(_00108_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_1 _24203_ (.A(net232),
    .B(_00074_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_1 _24204_ (.A(_00122_),
    .B(_00123_),
    .Y(_00125_));
 sky130_fd_sc_hd__nand2_1 _24205_ (.A(_00125_),
    .B(_11715_),
    .Y(_00126_));
 sky130_fd_sc_hd__nand3_2 _24206_ (.A(_00122_),
    .B(_11717_),
    .C(_00123_),
    .Y(_00127_));
 sky130_fd_sc_hd__nand2_1 _24207_ (.A(_00126_),
    .B(_00127_),
    .Y(_00128_));
 sky130_fd_sc_hd__nor2_1 _24208_ (.A(_00116_),
    .B(_00128_),
    .Y(_00129_));
 sky130_fd_sc_hd__nand2_1 _24209_ (.A(_00064_),
    .B(_00056_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _24210_ (.A(_00130_),
    .B(_14240_),
    .Y(_00131_));
 sky130_fd_sc_hd__nand2_1 _24211_ (.A(_00131_),
    .B(_14244_),
    .Y(_00132_));
 sky130_fd_sc_hd__nand2_1 _24212_ (.A(_00132_),
    .B(_14217_),
    .Y(_00133_));
 sky130_fd_sc_hd__nand3_1 _24213_ (.A(_00133_),
    .B(_14219_),
    .C(_14215_),
    .Y(_00134_));
 sky130_fd_sc_hd__nand2_1 _24214_ (.A(_14215_),
    .B(_14219_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand3_1 _24215_ (.A(_00132_),
    .B(_14217_),
    .C(_00136_),
    .Y(_00137_));
 sky130_fd_sc_hd__nand2_1 _24216_ (.A(_00134_),
    .B(_00137_),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2_1 _24217_ (.A(_00138_),
    .B(_00108_),
    .Y(_00139_));
 sky130_fd_sc_hd__nand2_1 _24218_ (.A(net232),
    .B(_14214_),
    .Y(_00140_));
 sky130_fd_sc_hd__nand3_1 _24219_ (.A(_00139_),
    .B(_12187_),
    .C(_00140_),
    .Y(_00141_));
 sky130_fd_sc_hd__or2_1 _24220_ (.A(_00086_),
    .B(_00066_),
    .X(_00142_));
 sky130_fd_sc_hd__nand3_1 _24221_ (.A(_00142_),
    .B(_00108_),
    .C(_00117_),
    .Y(_00143_));
 sky130_fd_sc_hd__nand2_1 _24222_ (.A(net232),
    .B(_00082_),
    .Y(_00144_));
 sky130_fd_sc_hd__nand3_1 _24223_ (.A(_00143_),
    .B(_13304_),
    .C(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__inv_2 _24224_ (.A(_00145_),
    .Y(_00147_));
 sky130_fd_sc_hd__a21o_1 _24225_ (.A1(_00143_),
    .A2(_00144_),
    .B1(_13304_),
    .X(_00148_));
 sky130_fd_sc_hd__o21ai_1 _24226_ (.A1(_00141_),
    .A2(_00147_),
    .B1(_00148_),
    .Y(_00149_));
 sky130_fd_sc_hd__inv_2 _24227_ (.A(_00115_),
    .Y(_00150_));
 sky130_fd_sc_hd__o21ai_1 _24228_ (.A1(_00127_),
    .A2(_00150_),
    .B1(_00114_),
    .Y(_00151_));
 sky130_fd_sc_hd__a21oi_1 _24229_ (.A1(_00129_),
    .A2(_00149_),
    .B1(_00151_),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _24230_ (.A(_14252_),
    .Y(_00153_));
 sky130_fd_sc_hd__nand2_1 _24231_ (.A(_14201_),
    .B(_00153_),
    .Y(_00154_));
 sky130_fd_sc_hd__nand2_1 _24232_ (.A(_14253_),
    .B(_14255_),
    .Y(_00155_));
 sky130_fd_sc_hd__xor2_1 _24233_ (.A(_14254_),
    .B(_00155_),
    .X(_00156_));
 sky130_fd_sc_hd__nand3b_1 _24234_ (.A_N(_00156_),
    .B(_14198_),
    .C(_14200_),
    .Y(_00158_));
 sky130_fd_sc_hd__nand2_1 _24235_ (.A(_00154_),
    .B(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__nand2_1 _24236_ (.A(_00159_),
    .B(_13679_),
    .Y(_00160_));
 sky130_fd_sc_hd__buf_6 _24237_ (.A(_12032_),
    .X(_00161_));
 sky130_fd_sc_hd__nor2_1 _24238_ (.A(_00161_),
    .B(_14046_),
    .Y(_00162_));
 sky130_fd_sc_hd__or2_1 _24239_ (.A(_11412_),
    .B(_00162_),
    .X(_00163_));
 sky130_fd_sc_hd__nand2_1 _24240_ (.A(_00163_),
    .B(_13693_),
    .Y(_00164_));
 sky130_fd_sc_hd__inv_2 _24241_ (.A(_00164_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _24242_ (.A(_14201_),
    .B(_00165_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand3_1 _24243_ (.A(_14198_),
    .B(_14200_),
    .C(_00162_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _24244_ (.A(_00166_),
    .B(_00167_),
    .Y(_00169_));
 sky130_fd_sc_hd__nand2_2 _24245_ (.A(_00169_),
    .B(_11421_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_1 _24246_ (.A(_00160_),
    .B(_00170_),
    .Y(_00171_));
 sky130_fd_sc_hd__inv_2 _24247_ (.A(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__nand3_1 _24248_ (.A(_00166_),
    .B(_11426_),
    .C(_00167_),
    .Y(_00173_));
 sky130_fd_sc_hd__buf_6 _24249_ (.A(_12033_),
    .X(_00174_));
 sky130_fd_sc_hd__nand3_2 _24250_ (.A(_14201_),
    .B(_00174_),
    .C(_12221_),
    .Y(_00175_));
 sky130_fd_sc_hd__inv_2 _24251_ (.A(_00175_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand3_2 _24252_ (.A(_00170_),
    .B(_00173_),
    .C(_00176_),
    .Y(_00177_));
 sky130_fd_sc_hd__or2_1 _24253_ (.A(_13679_),
    .B(_00159_),
    .X(_00178_));
 sky130_fd_sc_hd__a21boi_2 _24254_ (.A1(_00172_),
    .A2(_00177_),
    .B1_N(_00178_),
    .Y(_00180_));
 sky130_fd_sc_hd__clkinvlp_2 _24255_ (.A(_00044_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _24256_ (.A(_14202_),
    .B(_00181_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _24257_ (.A(_14285_),
    .B(_00049_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand3_1 _24258_ (.A(_14283_),
    .B(_00048_),
    .C(_14284_),
    .Y(_00184_));
 sky130_fd_sc_hd__nand2_1 _24259_ (.A(_00183_),
    .B(_00184_),
    .Y(_00185_));
 sky130_fd_sc_hd__inv_2 _24260_ (.A(_00185_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand3_1 _24261_ (.A(_14198_),
    .B(_14200_),
    .C(_00186_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _24262_ (.A(_00182_),
    .B(_00187_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _24263_ (.A(_00188_),
    .B(_11482_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand3_2 _24264_ (.A(_00182_),
    .B(_11484_),
    .C(_00187_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_2 _24265_ (.A(_00191_),
    .B(_00189_),
    .Y(_00192_));
 sky130_fd_sc_hd__inv_2 _24266_ (.A(_00192_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _24267_ (.A(_14202_),
    .B(_14281_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _24268_ (.A(_14284_),
    .B(_14282_),
    .Y(_00195_));
 sky130_fd_sc_hd__xor2_1 _24269_ (.A(_14278_),
    .B(_00195_),
    .X(_00196_));
 sky130_fd_sc_hd__nand3_1 _24270_ (.A(_14198_),
    .B(_14200_),
    .C(_00196_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand2_1 _24271_ (.A(_00194_),
    .B(_00197_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _24272_ (.A(_00198_),
    .B(_11496_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand3_2 _24273_ (.A(_00194_),
    .B(_11494_),
    .C(_00197_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_2 _24274_ (.A(_00200_),
    .B(_00199_),
    .Y(_00202_));
 sky130_fd_sc_hd__inv_2 _24275_ (.A(_00202_),
    .Y(_00203_));
 sky130_fd_sc_hd__nand2_1 _24276_ (.A(_00193_),
    .B(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__inv_2 _24277_ (.A(_14272_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _24278_ (.A(_14201_),
    .B(_00205_),
    .Y(_00206_));
 sky130_fd_sc_hd__or2_1 _24279_ (.A(_14276_),
    .B(_14266_),
    .X(_00207_));
 sky130_fd_sc_hd__nand2_1 _24280_ (.A(_00207_),
    .B(_14277_),
    .Y(_00208_));
 sky130_fd_sc_hd__inv_4 _24281_ (.A(_00208_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand3_1 _24282_ (.A(_14198_),
    .B(_14200_),
    .C(_00209_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _24283_ (.A(_00206_),
    .B(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _24284_ (.A(_00211_),
    .B(_11105_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand3_1 _24285_ (.A(_00206_),
    .B(_12261_),
    .C(_00210_),
    .Y(_00214_));
 sky130_fd_sc_hd__nand2_1 _24286_ (.A(_00213_),
    .B(_00214_),
    .Y(_00215_));
 sky130_fd_sc_hd__inv_2 _24287_ (.A(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _24288_ (.A(_14201_),
    .B(_14264_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_1 _24289_ (.A(_14265_),
    .B(_14262_),
    .Y(_00218_));
 sky130_fd_sc_hd__xnor2_1 _24290_ (.A(_14258_),
    .B(_00218_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand3_1 _24291_ (.A(_14198_),
    .B(_14200_),
    .C(_00219_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _24292_ (.A(_00217_),
    .B(_00220_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _24293_ (.A(_00221_),
    .B(_12270_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand3_1 _24294_ (.A(_00217_),
    .B(_11117_),
    .C(_00220_),
    .Y(_00224_));
 sky130_fd_sc_hd__nand2_2 _24295_ (.A(_00222_),
    .B(_00224_),
    .Y(_00225_));
 sky130_fd_sc_hd__inv_4 _24296_ (.A(_00225_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _24297_ (.A(_00216_),
    .B(_00226_),
    .Y(_00227_));
 sky130_fd_sc_hd__nor2_1 _24298_ (.A(_00204_),
    .B(_00227_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _24299_ (.A(_00180_),
    .B(_00228_),
    .Y(_00229_));
 sky130_fd_sc_hd__clkinvlp_2 _24300_ (.A(_00214_),
    .Y(_00230_));
 sky130_fd_sc_hd__o21ai_2 _24301_ (.A1(_00222_),
    .A2(_00230_),
    .B1(_00213_),
    .Y(_00231_));
 sky130_fd_sc_hd__nor2_1 _24302_ (.A(_00192_),
    .B(_00202_),
    .Y(_00232_));
 sky130_fd_sc_hd__inv_2 _24303_ (.A(_00191_),
    .Y(_00233_));
 sky130_fd_sc_hd__o21ai_1 _24304_ (.A1(_00200_),
    .A2(_00233_),
    .B1(_00189_),
    .Y(_00235_));
 sky130_fd_sc_hd__a21oi_1 _24305_ (.A1(_00231_),
    .A2(_00232_),
    .B1(_00235_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_2 _24306_ (.A(_00236_),
    .B(_00229_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _24307_ (.A(_00056_),
    .B(_00062_),
    .Y(_00238_));
 sky130_fd_sc_hd__or2_1 _24308_ (.A(_00062_),
    .B(_00056_),
    .X(_00239_));
 sky130_fd_sc_hd__nand3_1 _24309_ (.A(_00108_),
    .B(_00238_),
    .C(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _24310_ (.A(_14202_),
    .B(_14233_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _24311_ (.A(_00240_),
    .B(_00241_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _24312_ (.A(_00242_),
    .B(_11614_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand3_1 _24313_ (.A(_00240_),
    .B(_11616_),
    .C(_00241_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _24314_ (.A(_00243_),
    .B(_00244_),
    .Y(_00246_));
 sky130_fd_sc_hd__inv_2 _24315_ (.A(_00246_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _24316_ (.A(_00042_),
    .B(_00050_),
    .Y(_00248_));
 sky130_fd_sc_hd__nand2_1 _24317_ (.A(_00183_),
    .B(_00046_),
    .Y(_00249_));
 sky130_fd_sc_hd__xor2_1 _24318_ (.A(_00248_),
    .B(_00249_),
    .X(_00250_));
 sky130_fd_sc_hd__nand2_1 _24319_ (.A(_00250_),
    .B(_00108_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _24320_ (.A(_14202_),
    .B(_00041_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _24321_ (.A(_00251_),
    .B(_00252_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _24322_ (.A(_00253_),
    .B(_12771_),
    .Y(_00254_));
 sky130_fd_sc_hd__nand3_2 _24323_ (.A(_00251_),
    .B(_08951_),
    .C(_00252_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _24324_ (.A(_00254_),
    .B(_00255_),
    .Y(_00257_));
 sky130_fd_sc_hd__inv_2 _24325_ (.A(_00257_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _24326_ (.A(_00247_),
    .B(_00258_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _24327_ (.A(_00238_),
    .B(_14234_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _24328_ (.A(_00260_),
    .B(_00059_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand3_1 _24329_ (.A(_00238_),
    .B(_00057_),
    .C(_14234_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _24330_ (.A(_00261_),
    .B(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _24331_ (.A(_00263_),
    .B(_00108_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _24332_ (.A(_14202_),
    .B(_14229_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _24333_ (.A(_00264_),
    .B(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__nand2_1 _24334_ (.A(_00266_),
    .B(_11600_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand3_2 _24335_ (.A(_00264_),
    .B(_11603_),
    .C(_00265_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _24336_ (.A(_00268_),
    .B(_00269_),
    .Y(_00270_));
 sky130_fd_sc_hd__or2_1 _24337_ (.A(_14241_),
    .B(_00108_),
    .X(_00271_));
 sky130_fd_sc_hd__nand3_1 _24338_ (.A(_00130_),
    .B(_14243_),
    .C(_14240_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand3_1 _24339_ (.A(_00132_),
    .B(_00108_),
    .C(_00272_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _24340_ (.A(_00271_),
    .B(_00273_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _24341_ (.A(_00274_),
    .B(_11586_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand3_2 _24342_ (.A(_00271_),
    .B(_00273_),
    .C(_11588_),
    .Y(_00276_));
 sky130_fd_sc_hd__nand2_2 _24343_ (.A(_00275_),
    .B(_00276_),
    .Y(_00277_));
 sky130_fd_sc_hd__nor2_1 _24344_ (.A(_00270_),
    .B(_00277_),
    .Y(_00279_));
 sky130_fd_sc_hd__nor2b_1 _24345_ (.A(_00259_),
    .B_N(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _24346_ (.A(_00237_),
    .B(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__inv_2 _24347_ (.A(_00244_),
    .Y(_00282_));
 sky130_fd_sc_hd__o21ai_2 _24348_ (.A1(_00255_),
    .A2(_00282_),
    .B1(_00243_),
    .Y(_00283_));
 sky130_fd_sc_hd__inv_2 _24349_ (.A(_00276_),
    .Y(_00284_));
 sky130_fd_sc_hd__o21ai_1 _24350_ (.A1(_00269_),
    .A2(_00284_),
    .B1(_00275_),
    .Y(_00285_));
 sky130_fd_sc_hd__a21oi_1 _24351_ (.A1(_00279_),
    .A2(_00283_),
    .B1(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_2 _24352_ (.A(_00281_),
    .B(_00286_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_1 _24353_ (.A(_00139_),
    .B(_00140_),
    .Y(_00288_));
 sky130_fd_sc_hd__nand2_1 _24354_ (.A(_00288_),
    .B(_11185_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _24355_ (.A(_00290_),
    .B(_00141_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _24356_ (.A(_00148_),
    .B(_00145_),
    .Y(_00292_));
 sky130_fd_sc_hd__nor2_1 _24357_ (.A(_00291_),
    .B(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand3_2 _24358_ (.A(_00287_),
    .B(_00129_),
    .C(_00293_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_2 _24359_ (.A(_00152_),
    .B(_00294_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _24360_ (.A(_14079_),
    .B(_14080_),
    .Y(_00296_));
 sky130_fd_sc_hd__inv_2 _24361_ (.A(_00296_),
    .Y(_00297_));
 sky130_fd_sc_hd__or2_1 _24362_ (.A(_00297_),
    .B(_13992_),
    .X(_00298_));
 sky130_fd_sc_hd__nand2_1 _24363_ (.A(_13992_),
    .B(_00297_),
    .Y(_00299_));
 sky130_fd_sc_hd__nand2_1 _24364_ (.A(_00298_),
    .B(_00299_),
    .Y(_00301_));
 sky130_fd_sc_hd__inv_2 _24365_ (.A(_00301_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _24366_ (.A(_00302_),
    .B(_11199_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _24367_ (.A(_00301_),
    .B(_13461_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _24368_ (.A(_00303_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__inv_2 _24369_ (.A(_00305_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _24370_ (.A(_00098_),
    .B(_13965_),
    .Y(_00307_));
 sky130_fd_sc_hd__inv_2 _24371_ (.A(_13954_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _24372_ (.A(_00307_),
    .B(_00308_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand3_1 _24373_ (.A(_00098_),
    .B(_13954_),
    .C(_13965_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _24374_ (.A(_00309_),
    .B(_00310_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _24375_ (.A(_00312_),
    .B(_12894_),
    .Y(_00313_));
 sky130_fd_sc_hd__nand3_1 _24376_ (.A(_00309_),
    .B(_11754_),
    .C(_00310_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand3_1 _24377_ (.A(_00106_),
    .B(_00313_),
    .C(_00314_),
    .Y(_00315_));
 sky130_fd_sc_hd__inv_2 _24378_ (.A(_00315_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand3_1 _24379_ (.A(_00066_),
    .B(_00088_),
    .C(_00316_),
    .Y(_00317_));
 sky130_fd_sc_hd__inv_2 _24380_ (.A(_00313_),
    .Y(_00318_));
 sky130_fd_sc_hd__o21ai_1 _24381_ (.A1(_00103_),
    .A2(_00318_),
    .B1(_00314_),
    .Y(_00319_));
 sky130_fd_sc_hd__nor2_1 _24382_ (.A(_00092_),
    .B(_00315_),
    .Y(_00320_));
 sky130_fd_sc_hd__nor2_1 _24383_ (.A(_00319_),
    .B(_00320_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_2 _24384_ (.A(_00317_),
    .B(_00321_),
    .Y(_00323_));
 sky130_fd_sc_hd__or2_1 _24385_ (.A(_00306_),
    .B(_00323_),
    .X(_00324_));
 sky130_fd_sc_hd__buf_6 _24386_ (.A(_00108_),
    .X(_00325_));
 sky130_fd_sc_hd__nand2_1 _24387_ (.A(_00323_),
    .B(_00306_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand3_1 _24388_ (.A(_00324_),
    .B(_00325_),
    .C(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _24389_ (.A(\div1i.quot[4] ),
    .B(_00302_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _24390_ (.A(_00327_),
    .B(_00328_),
    .Y(_00329_));
 sky130_fd_sc_hd__xor2_2 _24391_ (.A(_06754_),
    .B(_00329_),
    .X(_00330_));
 sky130_fd_sc_hd__nand2_1 _24392_ (.A(_00313_),
    .B(_00314_),
    .Y(_00331_));
 sky130_fd_sc_hd__nand2_1 _24393_ (.A(_00107_),
    .B(_00103_),
    .Y(_00332_));
 sky130_fd_sc_hd__xor2_1 _24394_ (.A(_00331_),
    .B(_00332_),
    .X(_00334_));
 sky130_fd_sc_hd__nand2_1 _24395_ (.A(_00334_),
    .B(_00325_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _24396_ (.A(\div1i.quot[4] ),
    .B(_00312_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _24397_ (.A(_00335_),
    .B(_00336_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _24398_ (.A(_00337_),
    .B(_11838_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand3_1 _24399_ (.A(_00335_),
    .B(_11840_),
    .C(_00336_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _24400_ (.A(_00338_),
    .B(_00339_),
    .Y(_00340_));
 sky130_fd_sc_hd__nor2_1 _24401_ (.A(_00330_),
    .B(_00340_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _24402_ (.A(_00295_),
    .B(_00341_),
    .Y(_00342_));
 sky130_fd_sc_hd__nand2_1 _24403_ (.A(_00329_),
    .B(_13502_),
    .Y(_00343_));
 sky130_fd_sc_hd__o21a_1 _24404_ (.A1(_00339_),
    .A2(_00330_),
    .B1(_00343_),
    .X(_00345_));
 sky130_fd_sc_hd__nand2_1 _24405_ (.A(_00342_),
    .B(_00345_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _24406_ (.A(_13992_),
    .B(_14083_),
    .Y(_00347_));
 sky130_fd_sc_hd__inv_2 _24407_ (.A(_14086_),
    .Y(_00348_));
 sky130_fd_sc_hd__a21o_1 _24408_ (.A1(_00347_),
    .A2(_00348_),
    .B1(_14064_),
    .X(_00349_));
 sky130_fd_sc_hd__nand3_1 _24409_ (.A(_00347_),
    .B(_14064_),
    .C(_00348_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _24410_ (.A(_00349_),
    .B(_00350_),
    .Y(_00351_));
 sky130_fd_sc_hd__inv_2 _24411_ (.A(_00351_),
    .Y(_00352_));
 sky130_fd_sc_hd__nand2_1 _24412_ (.A(_00352_),
    .B(_11797_),
    .Y(_00353_));
 sky130_fd_sc_hd__nand2_1 _24413_ (.A(_00351_),
    .B(_12939_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand2_1 _24414_ (.A(_00353_),
    .B(_00354_),
    .Y(_00356_));
 sky130_fd_sc_hd__inv_4 _24415_ (.A(_00356_),
    .Y(_00357_));
 sky130_fd_sc_hd__nand2_1 _24416_ (.A(_00299_),
    .B(_14080_),
    .Y(_00358_));
 sky130_fd_sc_hd__xor2_2 _24417_ (.A(_14073_),
    .B(_00358_),
    .X(_00359_));
 sky130_fd_sc_hd__inv_2 _24418_ (.A(_00359_),
    .Y(_00360_));
 sky130_fd_sc_hd__nand2_1 _24419_ (.A(_00360_),
    .B(_11774_),
    .Y(_00361_));
 sky130_fd_sc_hd__nand2_1 _24420_ (.A(_00359_),
    .B(_12914_),
    .Y(_00362_));
 sky130_fd_sc_hd__nand2_1 _24421_ (.A(_00361_),
    .B(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__or2_1 _24422_ (.A(_00305_),
    .B(_00363_),
    .X(_00364_));
 sky130_fd_sc_hd__inv_4 _24423_ (.A(_00364_),
    .Y(_00365_));
 sky130_fd_sc_hd__nand2_1 _24424_ (.A(_00323_),
    .B(_00365_),
    .Y(_00367_));
 sky130_fd_sc_hd__inv_2 _24425_ (.A(_00303_),
    .Y(_00368_));
 sky130_fd_sc_hd__a21boi_1 _24426_ (.A1(_00368_),
    .A2(_00362_),
    .B1_N(_00361_),
    .Y(_00369_));
 sky130_fd_sc_hd__nand2_1 _24427_ (.A(_00367_),
    .B(_00369_),
    .Y(_00370_));
 sky130_fd_sc_hd__or2_1 _24428_ (.A(_00357_),
    .B(_00370_),
    .X(_00371_));
 sky130_fd_sc_hd__nand2_1 _24429_ (.A(_00370_),
    .B(_00357_),
    .Y(_00372_));
 sky130_fd_sc_hd__nand3_1 _24430_ (.A(_00371_),
    .B(_00325_),
    .C(_00372_),
    .Y(_00373_));
 sky130_fd_sc_hd__nand2_1 _24431_ (.A(\div1i.quot[4] ),
    .B(_00352_),
    .Y(_00374_));
 sky130_fd_sc_hd__nand2_1 _24432_ (.A(_00373_),
    .B(_00374_),
    .Y(_00375_));
 sky130_fd_sc_hd__xor2_2 _24433_ (.A(_11811_),
    .B(_00375_),
    .X(_00376_));
 sky130_fd_sc_hd__nand2_1 _24434_ (.A(_00326_),
    .B(_00303_),
    .Y(_00378_));
 sky130_fd_sc_hd__xor2_1 _24435_ (.A(_00363_),
    .B(_00378_),
    .X(_00379_));
 sky130_fd_sc_hd__nand2_1 _24436_ (.A(_00379_),
    .B(_00325_),
    .Y(_00380_));
 sky130_fd_sc_hd__nand2_1 _24437_ (.A(\div1i.quot[4] ),
    .B(_00359_),
    .Y(_00381_));
 sky130_fd_sc_hd__nand2_1 _24438_ (.A(_00380_),
    .B(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__or2_1 _24439_ (.A(_13537_),
    .B(_00382_),
    .X(_00383_));
 sky130_fd_sc_hd__nand2_1 _24440_ (.A(_00382_),
    .B(_13537_),
    .Y(_00384_));
 sky130_fd_sc_hd__nand2_1 _24441_ (.A(_00383_),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__nor2_1 _24442_ (.A(_00376_),
    .B(_00385_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _24443_ (.A(_00346_),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _24444_ (.A(_00375_),
    .B(_11808_),
    .Y(_00389_));
 sky130_fd_sc_hd__o21a_1 _24445_ (.A1(_00383_),
    .A2(_00376_),
    .B1(_00389_),
    .X(_00390_));
 sky130_fd_sc_hd__nand2_2 _24446_ (.A(_00387_),
    .B(_00390_),
    .Y(_00391_));
 sky130_fd_sc_hd__a21o_1 _24447_ (.A1(_14180_),
    .A2(_14183_),
    .B1(_14089_),
    .X(_00392_));
 sky130_fd_sc_hd__nand3_1 _24448_ (.A(_14089_),
    .B(_14180_),
    .C(_14183_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _24449_ (.A(_00392_),
    .B(_00393_),
    .Y(_00394_));
 sky130_fd_sc_hd__or2_1 _24450_ (.A(_14113_),
    .B(_00394_),
    .X(_00395_));
 sky130_fd_sc_hd__nand2_1 _24451_ (.A(_00394_),
    .B(_14113_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _24452_ (.A(_00395_),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__inv_4 _24453_ (.A(_00397_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _24454_ (.A(_00349_),
    .B(_14063_),
    .Y(_00400_));
 sky130_fd_sc_hd__inv_2 _24455_ (.A(_14054_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _24456_ (.A(_00400_),
    .B(_00401_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand3_1 _24457_ (.A(_00349_),
    .B(_14054_),
    .C(_14063_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _24458_ (.A(_00402_),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__nand2_1 _24459_ (.A(_00404_),
    .B(_12992_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand3_1 _24460_ (.A(_00402_),
    .B(_11858_),
    .C(_00403_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand3_1 _24461_ (.A(_00357_),
    .B(_00405_),
    .C(_00406_),
    .Y(_00407_));
 sky130_fd_sc_hd__inv_2 _24462_ (.A(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__nand3_1 _24463_ (.A(_00323_),
    .B(_00365_),
    .C(_00408_),
    .Y(_00409_));
 sky130_fd_sc_hd__inv_2 _24464_ (.A(_00353_),
    .Y(_00411_));
 sky130_fd_sc_hd__inv_2 _24465_ (.A(_00406_),
    .Y(_00412_));
 sky130_fd_sc_hd__a21o_1 _24466_ (.A1(_00405_),
    .A2(_00411_),
    .B1(_00412_),
    .X(_00413_));
 sky130_fd_sc_hd__nor2_1 _24467_ (.A(_00369_),
    .B(_00407_),
    .Y(_00414_));
 sky130_fd_sc_hd__nor2_1 _24468_ (.A(_00413_),
    .B(_00414_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_2 _24469_ (.A(_00409_),
    .B(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__or2_1 _24470_ (.A(_00398_),
    .B(_00416_),
    .X(_00417_));
 sky130_fd_sc_hd__nand2_1 _24471_ (.A(_00416_),
    .B(_00398_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _24472_ (.A(_00417_),
    .B(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _24473_ (.A(_00419_),
    .B(_00325_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _24474_ (.A(\div1i.quot[4] ),
    .B(_00394_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _24475_ (.A(_00420_),
    .B(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _24476_ (.A(_00423_),
    .B(_08020_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand3_1 _24477_ (.A(_00420_),
    .B(_13022_),
    .C(_00422_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_2 _24478_ (.A(_00424_),
    .B(_00425_),
    .Y(_00426_));
 sky130_fd_sc_hd__inv_2 _24479_ (.A(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__nand2_1 _24480_ (.A(_00405_),
    .B(_00406_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _24481_ (.A(_00372_),
    .B(_00353_),
    .Y(_00429_));
 sky130_fd_sc_hd__xor2_1 _24482_ (.A(_00428_),
    .B(_00429_),
    .X(_00430_));
 sky130_fd_sc_hd__nand2_1 _24483_ (.A(_00430_),
    .B(_00325_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _24484_ (.A(_00404_),
    .B(\div1i.quot[4] ),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _24485_ (.A(_00431_),
    .B(_00433_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _24486_ (.A(_00434_),
    .B(_11896_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand3_2 _24487_ (.A(_00431_),
    .B(_11899_),
    .C(_00433_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand3_1 _24488_ (.A(_00427_),
    .B(_00435_),
    .C(_00436_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _24489_ (.A(_00418_),
    .B(_00395_),
    .Y(_00438_));
 sky130_fd_sc_hd__nand2_1 _24490_ (.A(_00393_),
    .B(_14180_),
    .Y(_00439_));
 sky130_fd_sc_hd__xor2_2 _24491_ (.A(_14174_),
    .B(_00439_),
    .X(_00440_));
 sky130_fd_sc_hd__inv_2 _24492_ (.A(_00440_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand2_1 _24493_ (.A(_00441_),
    .B(_12495_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _24494_ (.A(_00440_),
    .B(_13042_),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _24495_ (.A(_00442_),
    .B(_00444_),
    .Y(_00445_));
 sky130_fd_sc_hd__inv_2 _24496_ (.A(_00445_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _24497_ (.A(_00438_),
    .B(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__nand3_1 _24498_ (.A(_00418_),
    .B(_00445_),
    .C(_00395_),
    .Y(_00448_));
 sky130_fd_sc_hd__nand2_1 _24499_ (.A(_00447_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _24500_ (.A(_00449_),
    .B(_00325_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _24501_ (.A(_00440_),
    .B(\div1i.quot[4] ),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _24502_ (.A(_00450_),
    .B(_00451_),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _24503_ (.A(_00452_),
    .B(_12506_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand3_1 _24504_ (.A(_00450_),
    .B(_11376_),
    .C(_00451_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _24505_ (.A(_00453_),
    .B(_00455_),
    .Y(_00456_));
 sky130_fd_sc_hd__inv_2 _24506_ (.A(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__nand2_1 _24507_ (.A(_00446_),
    .B(_00398_),
    .Y(_00458_));
 sky130_fd_sc_hd__inv_2 _24508_ (.A(_00458_),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _24509_ (.A(_00416_),
    .B(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__o21a_1 _24510_ (.A1(_00395_),
    .A2(_00445_),
    .B1(_00442_),
    .X(_00461_));
 sky130_fd_sc_hd__nand2_1 _24511_ (.A(_00460_),
    .B(_00461_),
    .Y(_00462_));
 sky130_fd_sc_hd__a21oi_1 _24512_ (.A1(_14084_),
    .A2(_14088_),
    .B1(_14184_),
    .Y(_00463_));
 sky130_fd_sc_hd__or2_1 _24513_ (.A(_14187_),
    .B(_00463_),
    .X(_00464_));
 sky130_fd_sc_hd__or2_1 _24514_ (.A(_14139_),
    .B(_00464_),
    .X(_00466_));
 sky130_fd_sc_hd__nand2_1 _24515_ (.A(_00464_),
    .B(_14139_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _24516_ (.A(_00466_),
    .B(_00467_),
    .Y(_00468_));
 sky130_fd_sc_hd__inv_2 _24517_ (.A(_00468_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _24518_ (.A(_00469_),
    .B(_11935_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _24519_ (.A(_00468_),
    .B(_13633_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _24520_ (.A(_00470_),
    .B(_00471_),
    .Y(_00472_));
 sky130_fd_sc_hd__inv_2 _24521_ (.A(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand2_1 _24522_ (.A(_00462_),
    .B(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand3_1 _24523_ (.A(_00460_),
    .B(_00461_),
    .C(_00472_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand3_1 _24524_ (.A(_00474_),
    .B(_00325_),
    .C(_00475_),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _24525_ (.A(_00469_),
    .B(\div1i.quot[4] ),
    .Y(_00478_));
 sky130_fd_sc_hd__nand2_1 _24526_ (.A(_00477_),
    .B(_00478_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _24527_ (.A(_00479_),
    .B(_11946_),
    .Y(_00480_));
 sky130_fd_sc_hd__nand3_1 _24528_ (.A(_00477_),
    .B(_11948_),
    .C(_00478_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_2 _24529_ (.A(_00480_),
    .B(_00481_),
    .Y(_00482_));
 sky130_fd_sc_hd__inv_2 _24530_ (.A(_00482_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _24531_ (.A(_00457_),
    .B(_00483_),
    .Y(_00484_));
 sky130_fd_sc_hd__nor2_1 _24532_ (.A(_00437_),
    .B(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_4 _24533_ (.A(_00391_),
    .B(_00485_),
    .Y(_00486_));
 sky130_fd_sc_hd__o21ai_1 _24534_ (.A1(_00436_),
    .A2(_00426_),
    .B1(_00425_),
    .Y(_00488_));
 sky130_fd_sc_hd__nor2_1 _24535_ (.A(_00482_),
    .B(_00456_),
    .Y(_00489_));
 sky130_fd_sc_hd__o21ai_1 _24536_ (.A1(_00455_),
    .A2(_00482_),
    .B1(_00480_),
    .Y(_00490_));
 sky130_fd_sc_hd__a21oi_2 _24537_ (.A1(_00488_),
    .A2(_00489_),
    .B1(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__nand2_4 _24538_ (.A(_00486_),
    .B(_00491_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _24539_ (.A(_00467_),
    .B(_14136_),
    .Y(_00493_));
 sky130_fd_sc_hd__xor2_2 _24540_ (.A(_14164_),
    .B(_00493_),
    .X(_00494_));
 sky130_fd_sc_hd__nand3_1 _24541_ (.A(_00474_),
    .B(_00325_),
    .C(_00470_),
    .Y(_00495_));
 sky130_fd_sc_hd__xnor2_2 _24542_ (.A(_00494_),
    .B(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_8 _24543_ (.A(_00492_),
    .B(_00496_),
    .Y(_00497_));
 sky130_fd_sc_hd__clkinvlp_2 _24544_ (.A(_00496_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand3_4 _24545_ (.A(_00486_),
    .B(_00491_),
    .C(_00499_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_8 _24546_ (.A(_00497_),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__buf_8 _24547_ (.A(_00501_),
    .X(_00502_));
 sky130_fd_sc_hd__buf_6 _24548_ (.A(net228),
    .X(\div1i.quot[3] ));
 sky130_fd_sc_hd__nand2_1 _24549_ (.A(_00170_),
    .B(_00173_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _24550_ (.A(_00503_),
    .B(_00175_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _24551_ (.A(_00504_),
    .B(_00177_),
    .Y(_00505_));
 sky130_fd_sc_hd__inv_2 _24552_ (.A(_00505_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _24553_ (.A(net228),
    .B(_00506_),
    .Y(_00507_));
 sky130_fd_sc_hd__o21ai_2 _24554_ (.A1(_00161_),
    .A2(\div1i.quot[4] ),
    .B1(_00174_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_1 _24555_ (.A(_00505_),
    .B(_12030_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand3_1 _24556_ (.A(_00504_),
    .B(_12035_),
    .C(_00177_),
    .Y(_00511_));
 sky130_fd_sc_hd__nand2_1 _24557_ (.A(_00510_),
    .B(_00511_),
    .Y(_00512_));
 sky130_fd_sc_hd__xor2_1 _24558_ (.A(_00509_),
    .B(_00512_),
    .X(_00513_));
 sky130_fd_sc_hd__nand3b_1 _24559_ (.A_N(_00513_),
    .B(_00497_),
    .C(_00500_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _24560_ (.A(_00507_),
    .B(_00514_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _24561_ (.A(_00515_),
    .B(_13679_),
    .Y(_00516_));
 sky130_fd_sc_hd__nor2_1 _24562_ (.A(_00161_),
    .B(_00325_),
    .Y(_00517_));
 sky130_fd_sc_hd__or2_1 _24563_ (.A(_11412_),
    .B(_00517_),
    .X(_00518_));
 sky130_fd_sc_hd__nand2_1 _24564_ (.A(_00518_),
    .B(_00175_),
    .Y(_00520_));
 sky130_fd_sc_hd__inv_2 _24565_ (.A(_00520_),
    .Y(_00521_));
 sky130_fd_sc_hd__nand2_1 _24566_ (.A(_00502_),
    .B(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand3_1 _24567_ (.A(_00497_),
    .B(_00500_),
    .C(_00517_),
    .Y(_00523_));
 sky130_fd_sc_hd__nand2_1 _24568_ (.A(_00522_),
    .B(_00523_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_2 _24569_ (.A(_00524_),
    .B(_11421_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _24570_ (.A(_00516_),
    .B(_00525_),
    .Y(_00526_));
 sky130_fd_sc_hd__inv_2 _24571_ (.A(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand3_1 _24572_ (.A(_00522_),
    .B(_11426_),
    .C(_00523_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand3_2 _24573_ (.A(_00502_),
    .B(_00174_),
    .C(_12221_),
    .Y(_00529_));
 sky130_fd_sc_hd__inv_2 _24574_ (.A(_00529_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand3_2 _24575_ (.A(_00525_),
    .B(_00528_),
    .C(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__or2_4 _24576_ (.A(_13679_),
    .B(_00515_),
    .X(_00533_));
 sky130_fd_sc_hd__inv_2 _24577_ (.A(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__a21oi_2 _24578_ (.A1(_00527_),
    .A2(_00532_),
    .B1(_00534_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _24579_ (.A(_00172_),
    .B(_00177_),
    .Y(_00536_));
 sky130_fd_sc_hd__nand2_1 _24580_ (.A(_00536_),
    .B(_00178_),
    .Y(_00537_));
 sky130_fd_sc_hd__inv_2 _24581_ (.A(_00231_),
    .Y(_00538_));
 sky130_fd_sc_hd__o21ai_1 _24582_ (.A1(_00227_),
    .A2(_00537_),
    .B1(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__or2_1 _24583_ (.A(_00203_),
    .B(_00539_),
    .X(_00540_));
 sky130_fd_sc_hd__nand2_1 _24584_ (.A(_00539_),
    .B(_00203_),
    .Y(_00542_));
 sky130_fd_sc_hd__nand2_1 _24585_ (.A(_00540_),
    .B(_00542_),
    .Y(_00543_));
 sky130_fd_sc_hd__inv_2 _24586_ (.A(_00543_),
    .Y(_00544_));
 sky130_fd_sc_hd__nand2_1 _24587_ (.A(_00501_),
    .B(_00544_),
    .Y(_00545_));
 sky130_fd_sc_hd__nand2_1 _24588_ (.A(_00544_),
    .B(_12087_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _24589_ (.A(_00543_),
    .B(_12085_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _24590_ (.A(_00546_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__inv_2 _24591_ (.A(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _24592_ (.A(_00180_),
    .B(_00226_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _24593_ (.A(_00537_),
    .B(_00225_),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_1 _24594_ (.A(_00550_),
    .B(_00551_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_1 _24595_ (.A(_00553_),
    .B(_12056_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand3_1 _24596_ (.A(_00550_),
    .B(_12058_),
    .C(_00551_),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _24597_ (.A(_00554_),
    .B(_00555_),
    .Y(_00556_));
 sky130_fd_sc_hd__inv_2 _24598_ (.A(_00556_),
    .Y(_00557_));
 sky130_fd_sc_hd__inv_2 _24599_ (.A(_00511_),
    .Y(_00558_));
 sky130_fd_sc_hd__a21o_1 _24600_ (.A1(_00510_),
    .A2(_00509_),
    .B1(_00558_),
    .X(_00559_));
 sky130_fd_sc_hd__nand2_1 _24601_ (.A(_00178_),
    .B(_00160_),
    .Y(_00560_));
 sky130_fd_sc_hd__nand2_1 _24602_ (.A(_00177_),
    .B(_00170_),
    .Y(_00561_));
 sky130_fd_sc_hd__xor2_1 _24603_ (.A(_00560_),
    .B(_00561_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _24604_ (.A(_00562_),
    .B(_12043_),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_1 _24605_ (.A(_00559_),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__inv_2 _24606_ (.A(_00562_),
    .Y(_00566_));
 sky130_fd_sc_hd__nand2_1 _24607_ (.A(_00566_),
    .B(_12047_),
    .Y(_00567_));
 sky130_fd_sc_hd__nand2_1 _24608_ (.A(_00565_),
    .B(_00567_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _24609_ (.A(_00557_),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_1 _24610_ (.A(_00569_),
    .B(_00555_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _24611_ (.A(_00550_),
    .B(_00222_),
    .Y(_00571_));
 sky130_fd_sc_hd__xor2_1 _24612_ (.A(_00215_),
    .B(_00571_),
    .X(_00572_));
 sky130_fd_sc_hd__nand2_1 _24613_ (.A(_00572_),
    .B(_13182_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _24614_ (.A(_00570_),
    .B(_00573_),
    .Y(_00575_));
 sky130_fd_sc_hd__inv_2 _24615_ (.A(_00572_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _24616_ (.A(_00576_),
    .B(_08176_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _24617_ (.A(_00575_),
    .B(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hd__or2_1 _24618_ (.A(_00549_),
    .B(_00578_),
    .X(_00579_));
 sky130_fd_sc_hd__nand2_1 _24619_ (.A(_00578_),
    .B(_00549_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_1 _24620_ (.A(_00579_),
    .B(_00580_),
    .Y(_00581_));
 sky130_fd_sc_hd__inv_2 _24621_ (.A(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand3_1 _24622_ (.A(_00497_),
    .B(_00500_),
    .C(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _24623_ (.A(_00545_),
    .B(_00583_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _24624_ (.A(_00584_),
    .B(_11482_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand3_1 _24625_ (.A(_00545_),
    .B(_11484_),
    .C(_00583_),
    .Y(_00587_));
 sky130_fd_sc_hd__nand2_1 _24626_ (.A(_00586_),
    .B(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__inv_2 _24627_ (.A(_00588_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _24628_ (.A(_00501_),
    .B(_00576_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _24629_ (.A(_00577_),
    .B(_00573_),
    .Y(_00591_));
 sky130_fd_sc_hd__xnor2_1 _24630_ (.A(_00570_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand3_1 _24631_ (.A(_00497_),
    .B(_00500_),
    .C(_00592_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _24632_ (.A(_00590_),
    .B(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _24633_ (.A(_00594_),
    .B(_11494_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand3_1 _24634_ (.A(_00590_),
    .B(_11496_),
    .C(_00593_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_2 _24635_ (.A(_00595_),
    .B(_00597_),
    .Y(_00598_));
 sky130_fd_sc_hd__inv_2 _24636_ (.A(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _24637_ (.A(_00589_),
    .B(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__inv_2 _24638_ (.A(_00553_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_1 _24639_ (.A(_00501_),
    .B(_00601_),
    .Y(_00602_));
 sky130_fd_sc_hd__or2_1 _24640_ (.A(_00568_),
    .B(_00557_),
    .X(_00603_));
 sky130_fd_sc_hd__nand2_1 _24641_ (.A(_00603_),
    .B(_00569_),
    .Y(_00604_));
 sky130_fd_sc_hd__inv_4 _24642_ (.A(_00604_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand3_1 _24643_ (.A(_00497_),
    .B(_00500_),
    .C(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__nand2_1 _24644_ (.A(_00602_),
    .B(_00606_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _24645_ (.A(_00608_),
    .B(_11105_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand3_1 _24646_ (.A(_00602_),
    .B(_12261_),
    .C(_00606_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_2 _24647_ (.A(_00609_),
    .B(_00610_),
    .Y(_00611_));
 sky130_fd_sc_hd__inv_2 _24648_ (.A(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _24649_ (.A(_00501_),
    .B(_00566_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _24650_ (.A(_00567_),
    .B(_00564_),
    .Y(_00614_));
 sky130_fd_sc_hd__xnor2_1 _24651_ (.A(_00559_),
    .B(_00614_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand3_1 _24652_ (.A(_00497_),
    .B(_00500_),
    .C(_00615_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _24653_ (.A(_00613_),
    .B(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _24654_ (.A(_00617_),
    .B(_12270_),
    .Y(_00619_));
 sky130_fd_sc_hd__nand3_1 _24655_ (.A(_00613_),
    .B(_11117_),
    .C(_00616_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _24656_ (.A(_00619_),
    .B(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hd__inv_2 _24657_ (.A(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _24658_ (.A(_00612_),
    .B(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__nor2_1 _24659_ (.A(_00600_),
    .B(_00623_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _24660_ (.A(_00535_),
    .B(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__inv_2 _24661_ (.A(_00610_),
    .Y(_00626_));
 sky130_fd_sc_hd__o21ai_2 _24662_ (.A1(_00619_),
    .A2(_00626_),
    .B1(_00609_),
    .Y(_00627_));
 sky130_fd_sc_hd__nor2_1 _24663_ (.A(_00588_),
    .B(_00598_),
    .Y(_00628_));
 sky130_fd_sc_hd__inv_2 _24664_ (.A(_00587_),
    .Y(_00630_));
 sky130_fd_sc_hd__o21ai_1 _24665_ (.A1(_00595_),
    .A2(_00630_),
    .B1(_00586_),
    .Y(_00631_));
 sky130_fd_sc_hd__a21oi_1 _24666_ (.A1(_00627_),
    .A2(_00628_),
    .B1(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_2 _24667_ (.A(_00625_),
    .B(_00632_),
    .Y(_00633_));
 sky130_fd_sc_hd__inv_2 _24668_ (.A(_00259_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _24669_ (.A(_00237_),
    .B(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hd__inv_2 _24670_ (.A(_00283_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _24671_ (.A(_00635_),
    .B(_00636_),
    .Y(_00637_));
 sky130_fd_sc_hd__inv_2 _24672_ (.A(_00270_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _24673_ (.A(_00637_),
    .B(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__nand3_1 _24674_ (.A(_00635_),
    .B(_00270_),
    .C(_00636_),
    .Y(_00641_));
 sky130_fd_sc_hd__nand2_1 _24675_ (.A(_00639_),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__inv_2 _24676_ (.A(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hd__nand2_1 _24677_ (.A(_00643_),
    .B(_11986_),
    .Y(_00644_));
 sky130_fd_sc_hd__nand2_1 _24678_ (.A(_00642_),
    .B(_12017_),
    .Y(_00645_));
 sky130_fd_sc_hd__nand2_1 _24679_ (.A(_00644_),
    .B(_00645_),
    .Y(_00646_));
 sky130_fd_sc_hd__inv_2 _24680_ (.A(_00646_),
    .Y(_00647_));
 sky130_fd_sc_hd__nand2_1 _24681_ (.A(_00542_),
    .B(_00200_),
    .Y(_00648_));
 sky130_fd_sc_hd__or2_1 _24682_ (.A(_00193_),
    .B(_00648_),
    .X(_00649_));
 sky130_fd_sc_hd__nand2_1 _24683_ (.A(_00648_),
    .B(_00193_),
    .Y(_00650_));
 sky130_fd_sc_hd__nand3_1 _24684_ (.A(_00649_),
    .B(_10939_),
    .C(_00650_),
    .Y(_00652_));
 sky130_fd_sc_hd__nand2_1 _24685_ (.A(_00652_),
    .B(_00546_),
    .Y(_00653_));
 sky130_fd_sc_hd__inv_2 _24686_ (.A(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__nand2_1 _24687_ (.A(_00580_),
    .B(_00654_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand2_2 _24688_ (.A(_00237_),
    .B(_00258_),
    .Y(_00656_));
 sky130_fd_sc_hd__nand2_1 _24689_ (.A(_00656_),
    .B(_00255_),
    .Y(_00657_));
 sky130_fd_sc_hd__xor2_1 _24690_ (.A(_00246_),
    .B(_00657_),
    .X(_00658_));
 sky130_fd_sc_hd__nand2_1 _24691_ (.A(_00658_),
    .B(_12002_),
    .Y(_00659_));
 sky130_fd_sc_hd__or2_1 _24692_ (.A(_00247_),
    .B(_00657_),
    .X(_00660_));
 sky130_fd_sc_hd__nand2_1 _24693_ (.A(_00657_),
    .B(_00247_),
    .Y(_00661_));
 sky130_fd_sc_hd__nand3_1 _24694_ (.A(_00660_),
    .B(_12012_),
    .C(_00661_),
    .Y(_00663_));
 sky130_fd_sc_hd__or2_1 _24695_ (.A(_00258_),
    .B(_00237_),
    .X(_00664_));
 sky130_fd_sc_hd__nand2_1 _24696_ (.A(_00664_),
    .B(_00656_),
    .Y(_00665_));
 sky130_fd_sc_hd__nand2_1 _24697_ (.A(_00665_),
    .B(_12101_),
    .Y(_00666_));
 sky130_fd_sc_hd__nand3_2 _24698_ (.A(_00664_),
    .B(_12008_),
    .C(_00656_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _24699_ (.A(_00666_),
    .B(_00667_),
    .Y(_00668_));
 sky130_fd_sc_hd__inv_2 _24700_ (.A(_00668_),
    .Y(_00669_));
 sky130_fd_sc_hd__nand3_1 _24701_ (.A(_00659_),
    .B(_00663_),
    .C(_00669_),
    .Y(_00670_));
 sky130_fd_sc_hd__inv_2 _24702_ (.A(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__nand2_1 _24703_ (.A(_00649_),
    .B(_00650_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand2_1 _24704_ (.A(_00672_),
    .B(_13197_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand3_2 _24705_ (.A(_00655_),
    .B(_00671_),
    .C(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__clkinvlp_2 _24706_ (.A(_00667_),
    .Y(_00676_));
 sky130_fd_sc_hd__a21boi_1 _24707_ (.A1(_00659_),
    .A2(_00676_),
    .B1_N(_00663_),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _24708_ (.A(_00675_),
    .B(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__or2_1 _24709_ (.A(_00647_),
    .B(_00678_),
    .X(_00679_));
 sky130_fd_sc_hd__inv_6 _24710_ (.A(_00501_),
    .Y(_00680_));
 sky130_fd_sc_hd__nand2_1 _24711_ (.A(_00678_),
    .B(_00647_),
    .Y(_00681_));
 sky130_fd_sc_hd__nand3_1 _24712_ (.A(_00679_),
    .B(_00680_),
    .C(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__nand2_1 _24713_ (.A(net228),
    .B(_00643_),
    .Y(_00683_));
 sky130_fd_sc_hd__nand2_1 _24714_ (.A(_00682_),
    .B(_00683_),
    .Y(_00685_));
 sky130_fd_sc_hd__nand2_1 _24715_ (.A(_00685_),
    .B(_11586_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand3_1 _24716_ (.A(_00682_),
    .B(_11588_),
    .C(_00683_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand2_1 _24717_ (.A(_00686_),
    .B(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__nand3_1 _24718_ (.A(_00655_),
    .B(_00674_),
    .C(_00669_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _24719_ (.A(_00689_),
    .B(_00667_),
    .Y(_00690_));
 sky130_fd_sc_hd__nand3_1 _24720_ (.A(_00690_),
    .B(_00663_),
    .C(_00659_),
    .Y(_00691_));
 sky130_fd_sc_hd__nand2_1 _24721_ (.A(_00659_),
    .B(_00663_),
    .Y(_00692_));
 sky130_fd_sc_hd__nand3_1 _24722_ (.A(_00689_),
    .B(_00692_),
    .C(_00667_),
    .Y(_00693_));
 sky130_fd_sc_hd__a21o_1 _24723_ (.A1(_00691_),
    .A2(_00693_),
    .B1(_00502_),
    .X(_00694_));
 sky130_fd_sc_hd__nand2_1 _24724_ (.A(_00502_),
    .B(_00658_),
    .Y(_00696_));
 sky130_fd_sc_hd__nand2_1 _24725_ (.A(_00694_),
    .B(_00696_),
    .Y(_00697_));
 sky130_fd_sc_hd__nand2_1 _24726_ (.A(_00697_),
    .B(_11600_),
    .Y(_00698_));
 sky130_fd_sc_hd__nand3_2 _24727_ (.A(_00694_),
    .B(_11603_),
    .C(_00696_),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _24728_ (.A(_00698_),
    .B(_00699_),
    .Y(_00700_));
 sky130_fd_sc_hd__nor2_2 _24729_ (.A(_00688_),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hd__a21o_1 _24730_ (.A1(_00655_),
    .A2(_00674_),
    .B1(_00669_),
    .X(_00702_));
 sky130_fd_sc_hd__nand3_1 _24731_ (.A(_00680_),
    .B(_00689_),
    .C(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__a21o_1 _24732_ (.A1(_00497_),
    .A2(_00500_),
    .B1(_00665_),
    .X(_00704_));
 sky130_fd_sc_hd__nand2_1 _24733_ (.A(_00703_),
    .B(_00704_),
    .Y(_00705_));
 sky130_fd_sc_hd__nand2_1 _24734_ (.A(_00705_),
    .B(_11614_),
    .Y(_00707_));
 sky130_fd_sc_hd__nand3_1 _24735_ (.A(_00703_),
    .B(_11616_),
    .C(_00704_),
    .Y(_00708_));
 sky130_fd_sc_hd__nand2_1 _24736_ (.A(_00707_),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _24737_ (.A(_00674_),
    .B(_00652_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand2_1 _24738_ (.A(_00580_),
    .B(_00546_),
    .Y(_00711_));
 sky130_fd_sc_hd__xor2_1 _24739_ (.A(_00710_),
    .B(_00711_),
    .X(_00712_));
 sky130_fd_sc_hd__nand2_1 _24740_ (.A(_00680_),
    .B(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__nand2_1 _24741_ (.A(_00502_),
    .B(_00672_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2_1 _24742_ (.A(_00713_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__or2_1 _24743_ (.A(_12771_),
    .B(_00715_),
    .X(_00716_));
 sky130_fd_sc_hd__nand2_1 _24744_ (.A(_00715_),
    .B(_12771_),
    .Y(_00718_));
 sky130_fd_sc_hd__nand2_1 _24745_ (.A(_00716_),
    .B(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__nor2_1 _24746_ (.A(_00709_),
    .B(_00719_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand2_1 _24747_ (.A(_00701_),
    .B(_00720_),
    .Y(_00721_));
 sky130_fd_sc_hd__inv_2 _24748_ (.A(_00721_),
    .Y(_00722_));
 sky130_fd_sc_hd__nand2_1 _24749_ (.A(_00633_),
    .B(_00722_),
    .Y(_00723_));
 sky130_fd_sc_hd__o21ai_1 _24750_ (.A1(_00716_),
    .A2(_00709_),
    .B1(_00707_),
    .Y(_00724_));
 sky130_fd_sc_hd__o21ai_1 _24751_ (.A1(_00699_),
    .A2(_00688_),
    .B1(_00686_),
    .Y(_00725_));
 sky130_fd_sc_hd__a21oi_1 _24752_ (.A1(_00724_),
    .A2(_00701_),
    .B1(_00725_),
    .Y(_00726_));
 sky130_fd_sc_hd__nand2_2 _24753_ (.A(_00723_),
    .B(_00726_),
    .Y(_00727_));
 sky130_fd_sc_hd__inv_2 _24754_ (.A(_00675_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand2_1 _24755_ (.A(_00639_),
    .B(_00269_),
    .Y(_00730_));
 sky130_fd_sc_hd__inv_2 _24756_ (.A(_00277_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _24757_ (.A(_00730_),
    .B(_00731_),
    .Y(_00732_));
 sky130_fd_sc_hd__nand3_1 _24758_ (.A(_00639_),
    .B(_00277_),
    .C(_00269_),
    .Y(_00733_));
 sky130_fd_sc_hd__nand2_1 _24759_ (.A(_00732_),
    .B(_00733_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _24760_ (.A(_00734_),
    .B(_11983_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand3_1 _24761_ (.A(_00732_),
    .B(_11990_),
    .C(_00733_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand3_1 _24762_ (.A(_00647_),
    .B(_00735_),
    .C(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__inv_2 _24763_ (.A(_00737_),
    .Y(_00738_));
 sky130_fd_sc_hd__nand2_1 _24764_ (.A(_00729_),
    .B(_00738_),
    .Y(_00740_));
 sky130_fd_sc_hd__nor2_1 _24765_ (.A(_00677_),
    .B(_00737_),
    .Y(_00741_));
 sky130_fd_sc_hd__nand2_1 _24766_ (.A(_00735_),
    .B(_00736_),
    .Y(_00742_));
 sky130_fd_sc_hd__o21ai_1 _24767_ (.A1(_00644_),
    .A2(_00742_),
    .B1(_00736_),
    .Y(_00743_));
 sky130_fd_sc_hd__nor2_1 _24768_ (.A(_00741_),
    .B(_00743_),
    .Y(_00744_));
 sky130_fd_sc_hd__nand2_1 _24769_ (.A(_00740_),
    .B(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__inv_2 _24770_ (.A(_00292_),
    .Y(_00746_));
 sky130_fd_sc_hd__inv_2 _24771_ (.A(_00291_),
    .Y(_00747_));
 sky130_fd_sc_hd__nand2_1 _24772_ (.A(_00287_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__nand2_1 _24773_ (.A(_00748_),
    .B(_00141_),
    .Y(_00749_));
 sky130_fd_sc_hd__or2_1 _24774_ (.A(_00746_),
    .B(_00749_),
    .X(_00751_));
 sky130_fd_sc_hd__nand2_1 _24775_ (.A(_00749_),
    .B(_00746_),
    .Y(_00752_));
 sky130_fd_sc_hd__nand2_1 _24776_ (.A(_00751_),
    .B(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _24777_ (.A(_00753_),
    .B(_12118_),
    .Y(_00754_));
 sky130_fd_sc_hd__nand3_1 _24778_ (.A(_00751_),
    .B(_12120_),
    .C(_00752_),
    .Y(_00755_));
 sky130_fd_sc_hd__nand2_1 _24779_ (.A(_00754_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__inv_2 _24780_ (.A(_00756_),
    .Y(_00757_));
 sky130_fd_sc_hd__or2_1 _24781_ (.A(_00747_),
    .B(_00287_),
    .X(_00758_));
 sky130_fd_sc_hd__nand2_1 _24782_ (.A(_00758_),
    .B(_00748_),
    .Y(_00759_));
 sky130_fd_sc_hd__inv_4 _24783_ (.A(_00759_),
    .Y(_00760_));
 sky130_fd_sc_hd__nand2_1 _24784_ (.A(_00760_),
    .B(_11671_),
    .Y(_00762_));
 sky130_fd_sc_hd__nand2_1 _24785_ (.A(_00759_),
    .B(_12817_),
    .Y(_00763_));
 sky130_fd_sc_hd__nand2_1 _24786_ (.A(_00762_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__inv_4 _24787_ (.A(_00764_),
    .Y(_00765_));
 sky130_fd_sc_hd__nand2_1 _24788_ (.A(_00757_),
    .B(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hd__inv_2 _24789_ (.A(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__nand2_1 _24790_ (.A(_00745_),
    .B(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__inv_2 _24791_ (.A(_00762_),
    .Y(_00769_));
 sky130_fd_sc_hd__a21boi_2 _24792_ (.A1(_00754_),
    .A2(_00769_),
    .B1_N(_00755_),
    .Y(_00770_));
 sky130_fd_sc_hd__nand2_1 _24793_ (.A(_00768_),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__nand2_1 _24794_ (.A(_00287_),
    .B(_00293_),
    .Y(_00773_));
 sky130_fd_sc_hd__inv_2 _24795_ (.A(_00149_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _24796_ (.A(_00773_),
    .B(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__inv_2 _24797_ (.A(_00128_),
    .Y(_00776_));
 sky130_fd_sc_hd__nand2_1 _24798_ (.A(_00775_),
    .B(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__nand3_1 _24799_ (.A(_00773_),
    .B(_00774_),
    .C(_00128_),
    .Y(_00778_));
 sky130_fd_sc_hd__nand2_1 _24800_ (.A(_00777_),
    .B(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hd__nand2_1 _24801_ (.A(_00779_),
    .B(_12149_),
    .Y(_00780_));
 sky130_fd_sc_hd__nand3_1 _24802_ (.A(_00777_),
    .B(_00778_),
    .C(_12147_),
    .Y(_00781_));
 sky130_fd_sc_hd__nand2_1 _24803_ (.A(_00780_),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _24804_ (.A(_00782_),
    .Y(_00784_));
 sky130_fd_sc_hd__nand2_1 _24805_ (.A(_00771_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hd__nand3_1 _24806_ (.A(_00768_),
    .B(_00782_),
    .C(_00770_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand3_1 _24807_ (.A(_00785_),
    .B(_00680_),
    .C(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__or2_1 _24808_ (.A(_00779_),
    .B(_00680_),
    .X(_00788_));
 sky130_fd_sc_hd__nand2_1 _24809_ (.A(_00787_),
    .B(_00788_),
    .Y(_00789_));
 sky130_fd_sc_hd__nand2_1 _24810_ (.A(_00789_),
    .B(_11701_),
    .Y(_00790_));
 sky130_fd_sc_hd__nand3_1 _24811_ (.A(_00787_),
    .B(_11703_),
    .C(_00788_),
    .Y(_00791_));
 sky130_fd_sc_hd__nand2_2 _24812_ (.A(_00790_),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__nand2_1 _24813_ (.A(_00745_),
    .B(_00765_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_1 _24814_ (.A(_00793_),
    .B(_00762_),
    .Y(_00795_));
 sky130_fd_sc_hd__nand2_1 _24815_ (.A(_00795_),
    .B(_00757_),
    .Y(_00796_));
 sky130_fd_sc_hd__nand3_1 _24816_ (.A(_00793_),
    .B(_00756_),
    .C(_00762_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand2_1 _24817_ (.A(_00796_),
    .B(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__nand2_1 _24818_ (.A(_00798_),
    .B(_00680_),
    .Y(_00799_));
 sky130_fd_sc_hd__nand2_1 _24819_ (.A(\div1i.quot[3] ),
    .B(_00753_),
    .Y(_00800_));
 sky130_fd_sc_hd__nand2_1 _24820_ (.A(_00799_),
    .B(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__nand2_1 _24821_ (.A(_00801_),
    .B(_11715_),
    .Y(_00802_));
 sky130_fd_sc_hd__nand3_2 _24822_ (.A(_00799_),
    .B(_11717_),
    .C(_00800_),
    .Y(_00803_));
 sky130_fd_sc_hd__nand2_1 _24823_ (.A(_00802_),
    .B(_00803_),
    .Y(_00804_));
 sky130_fd_sc_hd__nor2_1 _24824_ (.A(_00792_),
    .B(_00804_),
    .Y(_00806_));
 sky130_fd_sc_hd__or2_1 _24825_ (.A(_00765_),
    .B(_00745_),
    .X(_00807_));
 sky130_fd_sc_hd__nand3_1 _24826_ (.A(_00807_),
    .B(_00680_),
    .C(_00793_),
    .Y(_00808_));
 sky130_fd_sc_hd__nand2_1 _24827_ (.A(net228),
    .B(_00760_),
    .Y(_00809_));
 sky130_fd_sc_hd__nand2_1 _24828_ (.A(_00808_),
    .B(_00809_),
    .Y(_00810_));
 sky130_fd_sc_hd__nand2_1 _24829_ (.A(_00810_),
    .B(_06149_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand3_1 _24830_ (.A(_00808_),
    .B(_13304_),
    .C(_00809_),
    .Y(_00812_));
 sky130_fd_sc_hd__nand2_1 _24831_ (.A(_00811_),
    .B(_00812_),
    .Y(_00813_));
 sky130_fd_sc_hd__nand2_1 _24832_ (.A(_00681_),
    .B(_00644_),
    .Y(_00814_));
 sky130_fd_sc_hd__xor2_1 _24833_ (.A(_00742_),
    .B(_00814_),
    .X(_00815_));
 sky130_fd_sc_hd__nand2_1 _24834_ (.A(_00815_),
    .B(_00680_),
    .Y(_00817_));
 sky130_fd_sc_hd__nand2_1 _24835_ (.A(\div1i.quot[3] ),
    .B(_00734_),
    .Y(_00818_));
 sky130_fd_sc_hd__nand2_1 _24836_ (.A(_00817_),
    .B(_00818_),
    .Y(_00819_));
 sky130_fd_sc_hd__nand2_1 _24837_ (.A(_00819_),
    .B(_11185_),
    .Y(_00820_));
 sky130_fd_sc_hd__nand3_1 _24838_ (.A(_00817_),
    .B(_12187_),
    .C(_00818_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand2_1 _24839_ (.A(_00820_),
    .B(_00821_),
    .Y(_00822_));
 sky130_fd_sc_hd__nor2_1 _24840_ (.A(_00813_),
    .B(_00822_),
    .Y(_00823_));
 sky130_fd_sc_hd__nand2_1 _24841_ (.A(_00806_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__inv_2 _24842_ (.A(_00824_),
    .Y(_00825_));
 sky130_fd_sc_hd__nand2_1 _24843_ (.A(_00727_),
    .B(_00825_),
    .Y(_00826_));
 sky130_fd_sc_hd__o21ai_1 _24844_ (.A1(_00821_),
    .A2(_00813_),
    .B1(_00811_),
    .Y(_00828_));
 sky130_fd_sc_hd__o21ai_1 _24845_ (.A1(_00803_),
    .A2(_00792_),
    .B1(_00790_),
    .Y(_00829_));
 sky130_fd_sc_hd__a21oi_1 _24846_ (.A1(_00806_),
    .A2(_00828_),
    .B1(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__nand2_2 _24847_ (.A(_00826_),
    .B(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__nand2_1 _24848_ (.A(_00777_),
    .B(_00127_),
    .Y(_00832_));
 sky130_fd_sc_hd__inv_2 _24849_ (.A(_00116_),
    .Y(_00833_));
 sky130_fd_sc_hd__nand2_1 _24850_ (.A(_00832_),
    .B(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__nand3_1 _24851_ (.A(_00777_),
    .B(_00116_),
    .C(_00127_),
    .Y(_00835_));
 sky130_fd_sc_hd__nand2_1 _24852_ (.A(_00834_),
    .B(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__nand2_1 _24853_ (.A(_00836_),
    .B(_12894_),
    .Y(_00837_));
 sky130_fd_sc_hd__nand3_1 _24854_ (.A(_00834_),
    .B(_11754_),
    .C(_00835_),
    .Y(_00839_));
 sky130_fd_sc_hd__nand3_1 _24855_ (.A(_00837_),
    .B(_00839_),
    .C(_00784_),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2_1 _24856_ (.A(_00840_),
    .B(_00766_),
    .Y(_00841_));
 sky130_fd_sc_hd__nand2_1 _24857_ (.A(_00745_),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2_1 _24858_ (.A(_00840_),
    .B(_00770_),
    .Y(_00843_));
 sky130_fd_sc_hd__nand2_1 _24859_ (.A(_00837_),
    .B(_00839_),
    .Y(_00844_));
 sky130_fd_sc_hd__o21ai_1 _24860_ (.A1(_00781_),
    .A2(_00844_),
    .B1(_00839_),
    .Y(_00845_));
 sky130_fd_sc_hd__nor2_1 _24861_ (.A(_00843_),
    .B(_00845_),
    .Y(_00846_));
 sky130_fd_sc_hd__nand2_1 _24862_ (.A(_00842_),
    .B(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__clkinvlp_2 _24863_ (.A(_00330_),
    .Y(_00848_));
 sky130_fd_sc_hd__inv_2 _24864_ (.A(_00340_),
    .Y(_00850_));
 sky130_fd_sc_hd__nand2_1 _24865_ (.A(_00295_),
    .B(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__nand2_1 _24866_ (.A(_00851_),
    .B(_00339_),
    .Y(_00852_));
 sky130_fd_sc_hd__or2_1 _24867_ (.A(_00848_),
    .B(_00852_),
    .X(_00853_));
 sky130_fd_sc_hd__nand2_1 _24868_ (.A(_00852_),
    .B(_00848_),
    .Y(_00854_));
 sky130_fd_sc_hd__nand2_1 _24869_ (.A(_00853_),
    .B(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__nand2_1 _24870_ (.A(_00855_),
    .B(_12914_),
    .Y(_00856_));
 sky130_fd_sc_hd__nand3_1 _24871_ (.A(_00853_),
    .B(_11774_),
    .C(_00854_),
    .Y(_00857_));
 sky130_fd_sc_hd__nand2_1 _24872_ (.A(_00856_),
    .B(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__or2_1 _24873_ (.A(_00850_),
    .B(_00295_),
    .X(_00859_));
 sky130_fd_sc_hd__nand2_1 _24874_ (.A(_00859_),
    .B(_00851_),
    .Y(_00861_));
 sky130_fd_sc_hd__inv_2 _24875_ (.A(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _24876_ (.A(_00862_),
    .B(_11199_),
    .Y(_00863_));
 sky130_fd_sc_hd__nand2_1 _24877_ (.A(_00861_),
    .B(_13461_),
    .Y(_00864_));
 sky130_fd_sc_hd__nand2_1 _24878_ (.A(_00863_),
    .B(_00864_),
    .Y(_00865_));
 sky130_fd_sc_hd__inv_2 _24879_ (.A(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__nand2b_1 _24880_ (.A_N(_00858_),
    .B(_00866_),
    .Y(_00867_));
 sky130_fd_sc_hd__inv_2 _24881_ (.A(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__nand2_1 _24882_ (.A(_00847_),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _24883_ (.A(_00863_),
    .Y(_00870_));
 sky130_fd_sc_hd__a21boi_2 _24884_ (.A1(_00856_),
    .A2(_00870_),
    .B1_N(_00857_),
    .Y(_00872_));
 sky130_fd_sc_hd__nand2_1 _24885_ (.A(_00869_),
    .B(_00872_),
    .Y(_00873_));
 sky130_fd_sc_hd__inv_2 _24886_ (.A(_00385_),
    .Y(_00874_));
 sky130_fd_sc_hd__nand2_1 _24887_ (.A(_00346_),
    .B(_00874_),
    .Y(_00875_));
 sky130_fd_sc_hd__nand3_1 _24888_ (.A(_00342_),
    .B(_00345_),
    .C(_00385_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand2_1 _24889_ (.A(_00875_),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__inv_2 _24890_ (.A(_00877_),
    .Y(_00878_));
 sky130_fd_sc_hd__nand2_1 _24891_ (.A(_00878_),
    .B(_11797_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _24892_ (.A(_00877_),
    .B(_12939_),
    .Y(_00880_));
 sky130_fd_sc_hd__nand2_1 _24893_ (.A(_00879_),
    .B(_00880_),
    .Y(_00881_));
 sky130_fd_sc_hd__inv_2 _24894_ (.A(_00881_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand2_1 _24895_ (.A(_00873_),
    .B(_00883_),
    .Y(_00884_));
 sky130_fd_sc_hd__buf_6 _24896_ (.A(_00680_),
    .X(_00885_));
 sky130_fd_sc_hd__nand3_1 _24897_ (.A(_00869_),
    .B(_00881_),
    .C(_00872_),
    .Y(_00886_));
 sky130_fd_sc_hd__nand3_1 _24898_ (.A(_00884_),
    .B(_00885_),
    .C(_00886_),
    .Y(_00887_));
 sky130_fd_sc_hd__nand2_1 _24899_ (.A(\div1i.quot[3] ),
    .B(_00878_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_1 _24900_ (.A(_00887_),
    .B(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__nand2_1 _24901_ (.A(_00889_),
    .B(_11808_),
    .Y(_00890_));
 sky130_fd_sc_hd__nand3_1 _24902_ (.A(_00887_),
    .B(_11811_),
    .C(_00888_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_1 _24903_ (.A(_00890_),
    .B(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__nand2_1 _24904_ (.A(_00847_),
    .B(_00866_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_1 _24905_ (.A(_00894_),
    .B(_00863_),
    .Y(_00895_));
 sky130_fd_sc_hd__xor2_1 _24906_ (.A(_00858_),
    .B(_00895_),
    .X(_00896_));
 sky130_fd_sc_hd__nand2_1 _24907_ (.A(_00896_),
    .B(_00885_),
    .Y(_00897_));
 sky130_fd_sc_hd__nand2_1 _24908_ (.A(\div1i.quot[3] ),
    .B(_00855_),
    .Y(_00898_));
 sky130_fd_sc_hd__nand2_1 _24909_ (.A(_00897_),
    .B(_00898_),
    .Y(_00899_));
 sky130_fd_sc_hd__nand2_1 _24910_ (.A(_00899_),
    .B(_13537_),
    .Y(_00900_));
 sky130_fd_sc_hd__nand3_2 _24911_ (.A(_00897_),
    .B(_07400_),
    .C(_00898_),
    .Y(_00901_));
 sky130_fd_sc_hd__nand2_1 _24912_ (.A(_00900_),
    .B(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__nor2_1 _24913_ (.A(_00892_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__nand3_1 _24914_ (.A(_00842_),
    .B(_00846_),
    .C(_00865_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand3_1 _24915_ (.A(_00894_),
    .B(_00680_),
    .C(_00905_),
    .Y(_00906_));
 sky130_fd_sc_hd__nand2_1 _24916_ (.A(net228),
    .B(_00862_),
    .Y(_00907_));
 sky130_fd_sc_hd__nand2_1 _24917_ (.A(_00906_),
    .B(_00907_),
    .Y(_00908_));
 sky130_fd_sc_hd__or2_1 _24918_ (.A(_13502_),
    .B(_00908_),
    .X(_00909_));
 sky130_fd_sc_hd__nand2_1 _24919_ (.A(_00908_),
    .B(_13502_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand2_1 _24920_ (.A(_00909_),
    .B(_00910_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _24921_ (.A(_00785_),
    .B(_00781_),
    .Y(_00912_));
 sky130_fd_sc_hd__xor2_1 _24922_ (.A(_00844_),
    .B(_00912_),
    .X(_00913_));
 sky130_fd_sc_hd__nand2_1 _24923_ (.A(_00913_),
    .B(_00885_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand2_1 _24924_ (.A(\div1i.quot[3] ),
    .B(_00836_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand2_1 _24925_ (.A(_00914_),
    .B(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__nand2_1 _24926_ (.A(_00917_),
    .B(_11838_),
    .Y(_00918_));
 sky130_fd_sc_hd__nand3_2 _24927_ (.A(_00914_),
    .B(_11840_),
    .C(_00916_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand3b_1 _24928_ (.A_N(_00911_),
    .B(_00918_),
    .C(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__inv_4 _24929_ (.A(_00920_),
    .Y(_00921_));
 sky130_fd_sc_hd__nand3_1 _24930_ (.A(_00831_),
    .B(_00903_),
    .C(_00921_),
    .Y(_00922_));
 sky130_fd_sc_hd__inv_2 _24931_ (.A(_00910_),
    .Y(_00923_));
 sky130_fd_sc_hd__o21bai_1 _24932_ (.A1(_00911_),
    .A2(_00919_),
    .B1_N(_00923_),
    .Y(_00924_));
 sky130_fd_sc_hd__o21ai_1 _24933_ (.A1(_00892_),
    .A2(_00901_),
    .B1(_00890_),
    .Y(_00925_));
 sky130_fd_sc_hd__a21oi_1 _24934_ (.A1(_00903_),
    .A2(_00924_),
    .B1(_00925_),
    .Y(_00927_));
 sky130_fd_sc_hd__nand2_2 _24935_ (.A(_00922_),
    .B(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__nand2_1 _24936_ (.A(_00875_),
    .B(_00383_),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _24937_ (.A(_00376_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand2_1 _24938_ (.A(_00929_),
    .B(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand3_1 _24939_ (.A(_00875_),
    .B(_00376_),
    .C(_00383_),
    .Y(_00932_));
 sky130_fd_sc_hd__nand2_1 _24940_ (.A(_00931_),
    .B(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_1 _24941_ (.A(_00933_),
    .B(_12992_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand3_1 _24942_ (.A(_00931_),
    .B(_11858_),
    .C(_00932_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand3_1 _24943_ (.A(_00883_),
    .B(_00934_),
    .C(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__inv_2 _24944_ (.A(_00936_),
    .Y(_00938_));
 sky130_fd_sc_hd__nand3_1 _24945_ (.A(_00847_),
    .B(_00868_),
    .C(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__inv_2 _24946_ (.A(_00934_),
    .Y(_00940_));
 sky130_fd_sc_hd__o21ai_1 _24947_ (.A1(_00879_),
    .A2(_00940_),
    .B1(_00935_),
    .Y(_00941_));
 sky130_fd_sc_hd__nor2_1 _24948_ (.A(_00872_),
    .B(_00936_),
    .Y(_00942_));
 sky130_fd_sc_hd__nor2_1 _24949_ (.A(_00941_),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__nand2_1 _24950_ (.A(_00939_),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__inv_2 _24951_ (.A(_00391_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand2_1 _24952_ (.A(_00435_),
    .B(_00436_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _24953_ (.A(_00945_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__inv_2 _24954_ (.A(_00946_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_1 _24955_ (.A(_00391_),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand2_1 _24956_ (.A(_00947_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand2_1 _24957_ (.A(_00951_),
    .B(_14113_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand3_2 _24958_ (.A(_00947_),
    .B(_08554_),
    .C(_00950_),
    .Y(_00953_));
 sky130_fd_sc_hd__nand2_1 _24959_ (.A(_00952_),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__inv_2 _24960_ (.A(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand2_1 _24961_ (.A(_00944_),
    .B(_00955_),
    .Y(_00956_));
 sky130_fd_sc_hd__nand3_1 _24962_ (.A(_00939_),
    .B(_00943_),
    .C(_00954_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand3_1 _24963_ (.A(_00956_),
    .B(_00957_),
    .C(_00885_),
    .Y(_00958_));
 sky130_fd_sc_hd__or2_1 _24964_ (.A(_00951_),
    .B(_00885_),
    .X(_00960_));
 sky130_fd_sc_hd__nand2_1 _24965_ (.A(_00958_),
    .B(_00960_),
    .Y(_00961_));
 sky130_fd_sc_hd__or2_1 _24966_ (.A(_13022_),
    .B(_00961_),
    .X(_00962_));
 sky130_fd_sc_hd__nand2_1 _24967_ (.A(_00961_),
    .B(_13022_),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_1 _24968_ (.A(_00962_),
    .B(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hd__inv_2 _24969_ (.A(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _24970_ (.A(_00934_),
    .B(_00935_),
    .Y(_00966_));
 sky130_fd_sc_hd__nand2_1 _24971_ (.A(_00884_),
    .B(_00879_),
    .Y(_00967_));
 sky130_fd_sc_hd__xor2_1 _24972_ (.A(_00966_),
    .B(_00967_),
    .X(_00968_));
 sky130_fd_sc_hd__nand2_1 _24973_ (.A(_00968_),
    .B(_00885_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_1 _24974_ (.A(\div1i.quot[3] ),
    .B(_00933_),
    .Y(_00971_));
 sky130_fd_sc_hd__nand2_1 _24975_ (.A(_00969_),
    .B(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_1 _24976_ (.A(_00972_),
    .B(_11896_),
    .Y(_00973_));
 sky130_fd_sc_hd__nand3_2 _24977_ (.A(_00969_),
    .B(_11899_),
    .C(_00971_),
    .Y(_00974_));
 sky130_fd_sc_hd__nand3_1 _24978_ (.A(_00965_),
    .B(_00973_),
    .C(_00974_),
    .Y(_00975_));
 sky130_fd_sc_hd__nand2_1 _24979_ (.A(_00956_),
    .B(_00953_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_1 _24980_ (.A(_00950_),
    .B(_00436_),
    .Y(_00977_));
 sky130_fd_sc_hd__xor2_2 _24981_ (.A(_00426_),
    .B(_00977_),
    .X(_00978_));
 sky130_fd_sc_hd__inv_2 _24982_ (.A(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__nand2_1 _24983_ (.A(_00979_),
    .B(_12495_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _24984_ (.A(_00978_),
    .B(_13042_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _24985_ (.A(_00980_),
    .B(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__inv_2 _24986_ (.A(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _24987_ (.A(_00976_),
    .B(_00984_),
    .Y(_00985_));
 sky130_fd_sc_hd__nand3_1 _24988_ (.A(_00956_),
    .B(_00983_),
    .C(_00953_),
    .Y(_00986_));
 sky130_fd_sc_hd__nand2_1 _24989_ (.A(_00985_),
    .B(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__nand2_1 _24990_ (.A(_00987_),
    .B(_00885_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _24991_ (.A(_00978_),
    .B(\div1i.quot[3] ),
    .Y(_00989_));
 sky130_fd_sc_hd__nand2_1 _24992_ (.A(_00988_),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__nand2_1 _24993_ (.A(_00990_),
    .B(_12506_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand3_1 _24994_ (.A(_00988_),
    .B(_11376_),
    .C(_00989_),
    .Y(_00993_));
 sky130_fd_sc_hd__nand2_1 _24995_ (.A(_00991_),
    .B(_00993_),
    .Y(_00994_));
 sky130_fd_sc_hd__inv_2 _24996_ (.A(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__nand3_1 _24997_ (.A(_00980_),
    .B(_00982_),
    .C(_00955_),
    .Y(_00996_));
 sky130_fd_sc_hd__inv_2 _24998_ (.A(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_1 _24999_ (.A(_00997_),
    .B(_00944_),
    .Y(_00998_));
 sky130_fd_sc_hd__inv_2 _25000_ (.A(_00982_),
    .Y(_00999_));
 sky130_fd_sc_hd__o21a_1 _25001_ (.A1(_00953_),
    .A2(_00999_),
    .B1(_00980_),
    .X(_01000_));
 sky130_fd_sc_hd__nand2_1 _25002_ (.A(_00998_),
    .B(_01000_),
    .Y(_01001_));
 sky130_fd_sc_hd__o21bai_1 _25003_ (.A1(_00437_),
    .A2(_00945_),
    .B1_N(_00488_),
    .Y(_01002_));
 sky130_fd_sc_hd__or2_1 _25004_ (.A(_00457_),
    .B(_01002_),
    .X(_01004_));
 sky130_fd_sc_hd__nand2_1 _25005_ (.A(_01002_),
    .B(_00457_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand2_1 _25006_ (.A(_01004_),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__inv_2 _25007_ (.A(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__nand2_1 _25008_ (.A(_01007_),
    .B(_11935_),
    .Y(_01008_));
 sky130_fd_sc_hd__nand2_1 _25009_ (.A(_01006_),
    .B(_13633_),
    .Y(_01009_));
 sky130_fd_sc_hd__nand2_1 _25010_ (.A(_01008_),
    .B(_01009_),
    .Y(_01010_));
 sky130_fd_sc_hd__inv_2 _25011_ (.A(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__nand2_1 _25012_ (.A(_01001_),
    .B(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hd__nand3_1 _25013_ (.A(_00998_),
    .B(_01000_),
    .C(_01010_),
    .Y(_01013_));
 sky130_fd_sc_hd__nand3_1 _25014_ (.A(_01012_),
    .B(_01013_),
    .C(_00885_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _25015_ (.A(_01007_),
    .B(\div1i.quot[3] ),
    .Y(_01016_));
 sky130_fd_sc_hd__nand2_1 _25016_ (.A(_01015_),
    .B(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__nand2_1 _25017_ (.A(_01017_),
    .B(_11946_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand3_1 _25018_ (.A(_01015_),
    .B(_11948_),
    .C(_01016_),
    .Y(_01019_));
 sky130_fd_sc_hd__nand2_1 _25019_ (.A(_01018_),
    .B(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__inv_2 _25020_ (.A(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _25021_ (.A(_00995_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__nor2_1 _25022_ (.A(_00975_),
    .B(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__nand2_4 _25023_ (.A(_00928_),
    .B(_01023_),
    .Y(_01024_));
 sky130_fd_sc_hd__o21ai_1 _25024_ (.A1(_00964_),
    .A2(_00974_),
    .B1(_00963_),
    .Y(_01026_));
 sky130_fd_sc_hd__nor2_1 _25025_ (.A(_01020_),
    .B(_00994_),
    .Y(_01027_));
 sky130_fd_sc_hd__inv_2 _25026_ (.A(_01019_),
    .Y(_01028_));
 sky130_fd_sc_hd__o21ai_1 _25027_ (.A1(_00993_),
    .A2(_01028_),
    .B1(_01018_),
    .Y(_01029_));
 sky130_fd_sc_hd__a21oi_2 _25028_ (.A1(_01026_),
    .A2(_01027_),
    .B1(_01029_),
    .Y(_01030_));
 sky130_fd_sc_hd__nand2_2 _25029_ (.A(_01024_),
    .B(_01030_),
    .Y(_01031_));
 sky130_fd_sc_hd__nand2_1 _25030_ (.A(_01005_),
    .B(_00455_),
    .Y(_01032_));
 sky130_fd_sc_hd__xor2_1 _25031_ (.A(_00482_),
    .B(_01032_),
    .X(_01033_));
 sky130_fd_sc_hd__nand3_1 _25032_ (.A(_01012_),
    .B(_00885_),
    .C(_01008_),
    .Y(_01034_));
 sky130_fd_sc_hd__xnor2_2 _25033_ (.A(_01033_),
    .B(_01034_),
    .Y(_01035_));
 sky130_fd_sc_hd__nand2_4 _25034_ (.A(_01031_),
    .B(_01035_),
    .Y(_01037_));
 sky130_fd_sc_hd__clkinvlp_2 _25035_ (.A(_01035_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand3_4 _25036_ (.A(_01024_),
    .B(_01030_),
    .C(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__nand2_8 _25037_ (.A(_01037_),
    .B(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__buf_8 _25038_ (.A(_01040_),
    .X(_01041_));
 sky130_fd_sc_hd__buf_4 _25039_ (.A(_01041_),
    .X(\div1i.quot[2] ));
 sky130_fd_sc_hd__nand2_1 _25040_ (.A(_00633_),
    .B(_00720_),
    .Y(_01042_));
 sky130_fd_sc_hd__inv_2 _25041_ (.A(_00724_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand2_1 _25042_ (.A(_01042_),
    .B(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__inv_2 _25043_ (.A(_00700_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand2_1 _25044_ (.A(_01044_),
    .B(_01045_),
    .Y(_01047_));
 sky130_fd_sc_hd__nand2_1 _25045_ (.A(_01047_),
    .B(_00699_),
    .Y(_01048_));
 sky130_fd_sc_hd__inv_2 _25046_ (.A(_00688_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand2_1 _25047_ (.A(_01048_),
    .B(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand3_1 _25048_ (.A(_01047_),
    .B(_00688_),
    .C(_00699_),
    .Y(_01051_));
 sky130_fd_sc_hd__nand2_1 _25049_ (.A(_01050_),
    .B(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__nand2_1 _25050_ (.A(_01052_),
    .B(_11983_),
    .Y(_01053_));
 sky130_fd_sc_hd__nand3_1 _25051_ (.A(_01042_),
    .B(_00700_),
    .C(_01043_),
    .Y(_01054_));
 sky130_fd_sc_hd__nand3_2 _25052_ (.A(_01047_),
    .B(_11986_),
    .C(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__inv_2 _25053_ (.A(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__nand3_2 _25054_ (.A(_01050_),
    .B(_11990_),
    .C(_01051_),
    .Y(_01058_));
 sky130_fd_sc_hd__nand3_1 _25055_ (.A(_01053_),
    .B(_01056_),
    .C(_01058_),
    .Y(_01059_));
 sky130_fd_sc_hd__nand2_1 _25056_ (.A(_01059_),
    .B(_01058_),
    .Y(_01060_));
 sky130_fd_sc_hd__inv_2 _25057_ (.A(_00719_),
    .Y(_01061_));
 sky130_fd_sc_hd__nand2_1 _25058_ (.A(_00633_),
    .B(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__nand2_1 _25059_ (.A(_01062_),
    .B(_00716_),
    .Y(_01063_));
 sky130_fd_sc_hd__inv_2 _25060_ (.A(_00709_),
    .Y(_01064_));
 sky130_fd_sc_hd__nand2_1 _25061_ (.A(_01063_),
    .B(_01064_),
    .Y(_01065_));
 sky130_fd_sc_hd__nand3_1 _25062_ (.A(_01062_),
    .B(_00709_),
    .C(_00716_),
    .Y(_01066_));
 sky130_fd_sc_hd__nand2_1 _25063_ (.A(_01065_),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _25064_ (.A(_01067_),
    .B(_12002_),
    .Y(_01069_));
 sky130_fd_sc_hd__or2_1 _25065_ (.A(_01061_),
    .B(_00633_),
    .X(_01070_));
 sky130_fd_sc_hd__nand2_1 _25066_ (.A(_01070_),
    .B(_01062_),
    .Y(_01071_));
 sky130_fd_sc_hd__inv_2 _25067_ (.A(_01071_),
    .Y(_01072_));
 sky130_fd_sc_hd__nand2_1 _25068_ (.A(_01072_),
    .B(_12008_),
    .Y(_01073_));
 sky130_fd_sc_hd__inv_2 _25069_ (.A(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__inv_2 _25070_ (.A(_01067_),
    .Y(_01075_));
 sky130_fd_sc_hd__nand2_1 _25071_ (.A(_01075_),
    .B(_12012_),
    .Y(_01076_));
 sky130_fd_sc_hd__inv_2 _25072_ (.A(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__a21oi_2 _25073_ (.A1(_01069_),
    .A2(_01074_),
    .B1(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand2_1 _25074_ (.A(_01047_),
    .B(_01054_),
    .Y(_01080_));
 sky130_fd_sc_hd__nand2_1 _25075_ (.A(_01080_),
    .B(_12017_),
    .Y(_01081_));
 sky130_fd_sc_hd__nand2_1 _25076_ (.A(_01081_),
    .B(_01055_),
    .Y(_01082_));
 sky130_fd_sc_hd__inv_2 _25077_ (.A(_01082_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand3_1 _25078_ (.A(_01053_),
    .B(_01083_),
    .C(_01058_),
    .Y(_01084_));
 sky130_fd_sc_hd__nor2_1 _25079_ (.A(_01078_),
    .B(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__nor2_1 _25080_ (.A(_01060_),
    .B(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__inv_2 _25081_ (.A(_01084_),
    .Y(_01087_));
 sky130_fd_sc_hd__nand2_1 _25082_ (.A(_00525_),
    .B(_00528_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2_1 _25083_ (.A(_01088_),
    .B(_00529_),
    .Y(_01089_));
 sky130_fd_sc_hd__nand2_1 _25084_ (.A(_01089_),
    .B(_00532_),
    .Y(_01091_));
 sky130_fd_sc_hd__nand2_1 _25085_ (.A(_01091_),
    .B(_12030_),
    .Y(_01092_));
 sky130_fd_sc_hd__o21ai_2 _25086_ (.A1(_00161_),
    .A2(\div1i.quot[3] ),
    .B1(_00174_),
    .Y(_01093_));
 sky130_fd_sc_hd__nand3_1 _25087_ (.A(_01089_),
    .B(_12035_),
    .C(_00532_),
    .Y(_01094_));
 sky130_fd_sc_hd__inv_2 _25088_ (.A(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hd__a21o_1 _25089_ (.A1(_01092_),
    .A2(_01093_),
    .B1(_01095_),
    .X(_01096_));
 sky130_fd_sc_hd__nand2_1 _25090_ (.A(_00533_),
    .B(_00516_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_1 _25091_ (.A(_00532_),
    .B(_00525_),
    .Y(_01098_));
 sky130_fd_sc_hd__xor2_2 _25092_ (.A(_01097_),
    .B(_01098_),
    .X(_01099_));
 sky130_fd_sc_hd__nand2_1 _25093_ (.A(_01099_),
    .B(_12043_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_1 _25094_ (.A(_01096_),
    .B(_01100_),
    .Y(_01102_));
 sky130_fd_sc_hd__inv_2 _25095_ (.A(_01099_),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _25096_ (.A(_01103_),
    .B(_12047_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _25097_ (.A(_01102_),
    .B(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand2_1 _25098_ (.A(_00527_),
    .B(_00532_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand2_1 _25099_ (.A(_01106_),
    .B(_00533_),
    .Y(_01107_));
 sky130_fd_sc_hd__nand2_1 _25100_ (.A(_01107_),
    .B(_00621_),
    .Y(_01108_));
 sky130_fd_sc_hd__nand3_1 _25101_ (.A(_01106_),
    .B(_00533_),
    .C(_00622_),
    .Y(_01109_));
 sky130_fd_sc_hd__nand2_1 _25102_ (.A(_01108_),
    .B(_01109_),
    .Y(_01110_));
 sky130_fd_sc_hd__nand2_1 _25103_ (.A(_01110_),
    .B(_12056_),
    .Y(_01111_));
 sky130_fd_sc_hd__nand3_1 _25104_ (.A(_01108_),
    .B(_12058_),
    .C(_01109_),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _25105_ (.A(_01111_),
    .B(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__inv_2 _25106_ (.A(_01114_),
    .Y(_01115_));
 sky130_fd_sc_hd__nand2_1 _25107_ (.A(_01105_),
    .B(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _25108_ (.A(_01116_),
    .B(_01113_),
    .Y(_01117_));
 sky130_fd_sc_hd__nand2_1 _25109_ (.A(_01109_),
    .B(_00619_),
    .Y(_01118_));
 sky130_fd_sc_hd__xor2_2 _25110_ (.A(_00611_),
    .B(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__nand2_1 _25111_ (.A(_01119_),
    .B(_13182_),
    .Y(_01120_));
 sky130_fd_sc_hd__nand2_1 _25112_ (.A(_01117_),
    .B(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__or2_1 _25113_ (.A(_13182_),
    .B(_01119_),
    .X(_01122_));
 sky130_fd_sc_hd__nand2_1 _25114_ (.A(_01121_),
    .B(_01122_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _25115_ (.A(_00611_),
    .B(_00621_),
    .Y(_01125_));
 sky130_fd_sc_hd__nand3_1 _25116_ (.A(_01106_),
    .B(_01125_),
    .C(_00533_),
    .Y(_01126_));
 sky130_fd_sc_hd__inv_2 _25117_ (.A(_00627_),
    .Y(_01127_));
 sky130_fd_sc_hd__nand2_1 _25118_ (.A(_01126_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__nand2_1 _25119_ (.A(_01128_),
    .B(_00599_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_1 _25120_ (.A(_01129_),
    .B(_00595_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _25121_ (.A(_01130_),
    .B(_00589_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand3_1 _25122_ (.A(_01129_),
    .B(_00588_),
    .C(_00595_),
    .Y(_01132_));
 sky130_fd_sc_hd__nand2_1 _25123_ (.A(_01131_),
    .B(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__nand2_1 _25124_ (.A(_01133_),
    .B(_13197_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand3_1 _25125_ (.A(_01126_),
    .B(_00598_),
    .C(_01127_),
    .Y(_01136_));
 sky130_fd_sc_hd__nand2_1 _25126_ (.A(_01129_),
    .B(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__nand2_1 _25127_ (.A(_01137_),
    .B(_12085_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand3_2 _25128_ (.A(_01129_),
    .B(_12087_),
    .C(_01136_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand2_1 _25129_ (.A(_01138_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__inv_2 _25130_ (.A(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand3_1 _25131_ (.A(_01131_),
    .B(_10939_),
    .C(_01132_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand3_1 _25132_ (.A(_01135_),
    .B(_01141_),
    .C(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__inv_2 _25133_ (.A(_01143_),
    .Y(_01144_));
 sky130_fd_sc_hd__nand2_1 _25134_ (.A(_01124_),
    .B(_01144_),
    .Y(_01146_));
 sky130_fd_sc_hd__inv_2 _25135_ (.A(_01139_),
    .Y(_01147_));
 sky130_fd_sc_hd__a21boi_1 _25136_ (.A1(_01135_),
    .A2(_01147_),
    .B1_N(_01142_),
    .Y(_01148_));
 sky130_fd_sc_hd__nand2_1 _25137_ (.A(_01146_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__nand2_1 _25138_ (.A(_01076_),
    .B(_01069_),
    .Y(_01150_));
 sky130_fd_sc_hd__inv_2 _25139_ (.A(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hd__nand2_1 _25140_ (.A(_01071_),
    .B(_12101_),
    .Y(_01152_));
 sky130_fd_sc_hd__nand2_1 _25141_ (.A(_01073_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__inv_2 _25142_ (.A(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand2_1 _25143_ (.A(_01151_),
    .B(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__inv_2 _25144_ (.A(_01155_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand3_1 _25145_ (.A(_01087_),
    .B(_01149_),
    .C(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__nand2_2 _25146_ (.A(_01086_),
    .B(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__inv_2 _25147_ (.A(_00813_),
    .Y(_01160_));
 sky130_fd_sc_hd__inv_2 _25148_ (.A(_00822_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2_1 _25149_ (.A(_00727_),
    .B(_01161_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2_1 _25150_ (.A(_01162_),
    .B(_00821_),
    .Y(_01163_));
 sky130_fd_sc_hd__or2_1 _25151_ (.A(_01160_),
    .B(_01163_),
    .X(_01164_));
 sky130_fd_sc_hd__nand2_1 _25152_ (.A(_01163_),
    .B(_01160_),
    .Y(_01165_));
 sky130_fd_sc_hd__nand2_1 _25153_ (.A(_01164_),
    .B(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand2_1 _25154_ (.A(_01166_),
    .B(_12118_),
    .Y(_01168_));
 sky130_fd_sc_hd__nand3_1 _25155_ (.A(_01164_),
    .B(_12120_),
    .C(_01165_),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_1 _25156_ (.A(_01168_),
    .B(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__inv_2 _25157_ (.A(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__or2_1 _25158_ (.A(_01161_),
    .B(_00727_),
    .X(_01172_));
 sky130_fd_sc_hd__nand2_1 _25159_ (.A(_01172_),
    .B(_01162_),
    .Y(_01173_));
 sky130_fd_sc_hd__inv_2 _25160_ (.A(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__nand2_2 _25161_ (.A(_01174_),
    .B(_11671_),
    .Y(_01175_));
 sky130_fd_sc_hd__nand2_1 _25162_ (.A(_01173_),
    .B(_12817_),
    .Y(_01176_));
 sky130_fd_sc_hd__nand2_1 _25163_ (.A(_01175_),
    .B(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__inv_2 _25164_ (.A(_01177_),
    .Y(_01179_));
 sky130_fd_sc_hd__nand2_1 _25165_ (.A(_01171_),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__inv_2 _25166_ (.A(_01180_),
    .Y(_01181_));
 sky130_fd_sc_hd__nand2_1 _25167_ (.A(_01159_),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__inv_2 _25168_ (.A(_01175_),
    .Y(_01183_));
 sky130_fd_sc_hd__a21boi_2 _25169_ (.A1(_01168_),
    .A2(_01183_),
    .B1_N(_01169_),
    .Y(_01184_));
 sky130_fd_sc_hd__nand2_1 _25170_ (.A(_01182_),
    .B(_01184_),
    .Y(_01185_));
 sky130_fd_sc_hd__nand2_1 _25171_ (.A(_00727_),
    .B(_00823_),
    .Y(_01186_));
 sky130_fd_sc_hd__inv_2 _25172_ (.A(_00828_),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _25173_ (.A(_01186_),
    .B(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__inv_2 _25174_ (.A(_00804_),
    .Y(_01190_));
 sky130_fd_sc_hd__nand2_1 _25175_ (.A(_01188_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hd__nand3_1 _25176_ (.A(_01186_),
    .B(_00804_),
    .C(_01187_),
    .Y(_01192_));
 sky130_fd_sc_hd__nand2_1 _25177_ (.A(_01191_),
    .B(_01192_),
    .Y(_01193_));
 sky130_fd_sc_hd__inv_2 _25178_ (.A(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__nand2_1 _25179_ (.A(_01194_),
    .B(_12147_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand2_1 _25180_ (.A(_01193_),
    .B(_12149_),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_1 _25181_ (.A(_01195_),
    .B(_01196_),
    .Y(_01197_));
 sky130_fd_sc_hd__inv_2 _25182_ (.A(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__nand2_1 _25183_ (.A(_01185_),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__inv_6 _25184_ (.A(_01040_),
    .Y(_01201_));
 sky130_fd_sc_hd__nand3_1 _25185_ (.A(_01182_),
    .B(_01197_),
    .C(_01184_),
    .Y(_01202_));
 sky130_fd_sc_hd__nand3_1 _25186_ (.A(_01199_),
    .B(_01201_),
    .C(_01202_),
    .Y(_01203_));
 sky130_fd_sc_hd__nand2_1 _25187_ (.A(_01041_),
    .B(_01194_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _25188_ (.A(_01203_),
    .B(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__nand2_1 _25189_ (.A(_01205_),
    .B(_11701_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand3_1 _25190_ (.A(_01203_),
    .B(_11703_),
    .C(_01204_),
    .Y(_01207_));
 sky130_fd_sc_hd__nand2_1 _25191_ (.A(_01206_),
    .B(_01207_),
    .Y(_01208_));
 sky130_fd_sc_hd__nand2_1 _25192_ (.A(_01159_),
    .B(_01179_),
    .Y(_01209_));
 sky130_fd_sc_hd__nand2_1 _25193_ (.A(_01209_),
    .B(_01175_),
    .Y(_01210_));
 sky130_fd_sc_hd__nand2_1 _25194_ (.A(_01210_),
    .B(_01171_),
    .Y(_01212_));
 sky130_fd_sc_hd__nand3_1 _25195_ (.A(_01209_),
    .B(_01170_),
    .C(_01175_),
    .Y(_01213_));
 sky130_fd_sc_hd__nand2_1 _25196_ (.A(_01212_),
    .B(_01213_),
    .Y(_01214_));
 sky130_fd_sc_hd__nand2_1 _25197_ (.A(_01214_),
    .B(_01201_),
    .Y(_01215_));
 sky130_fd_sc_hd__nand2_1 _25198_ (.A(_01041_),
    .B(_01166_),
    .Y(_01216_));
 sky130_fd_sc_hd__nand2_1 _25199_ (.A(_01215_),
    .B(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_1 _25200_ (.A(_01217_),
    .B(_11715_),
    .Y(_01218_));
 sky130_fd_sc_hd__nand3_2 _25201_ (.A(_01215_),
    .B(_11717_),
    .C(_01216_),
    .Y(_01219_));
 sky130_fd_sc_hd__nand2_1 _25202_ (.A(_01218_),
    .B(_01219_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor2_1 _25203_ (.A(_01208_),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__nand2_1 _25204_ (.A(_01157_),
    .B(_01149_),
    .Y(_01223_));
 sky130_fd_sc_hd__nand2_1 _25205_ (.A(_01223_),
    .B(_01078_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand2_1 _25206_ (.A(_01224_),
    .B(_01083_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_1 _25207_ (.A(_01225_),
    .B(_01055_),
    .Y(_01226_));
 sky130_fd_sc_hd__nand3_1 _25208_ (.A(_01226_),
    .B(_01058_),
    .C(_01053_),
    .Y(_01227_));
 sky130_fd_sc_hd__nand2_1 _25209_ (.A(_01053_),
    .B(_01058_),
    .Y(_01228_));
 sky130_fd_sc_hd__nand3_1 _25210_ (.A(_01225_),
    .B(_01055_),
    .C(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__nand2_1 _25211_ (.A(_01227_),
    .B(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2_1 _25212_ (.A(_01230_),
    .B(_01201_),
    .Y(_01231_));
 sky130_fd_sc_hd__nand2_1 _25213_ (.A(_01041_),
    .B(_01052_),
    .Y(_01232_));
 sky130_fd_sc_hd__nand3_2 _25214_ (.A(_01231_),
    .B(_12187_),
    .C(_01232_),
    .Y(_01234_));
 sky130_fd_sc_hd__or2_1 _25215_ (.A(_01179_),
    .B(_01159_),
    .X(_01235_));
 sky130_fd_sc_hd__nand3_1 _25216_ (.A(_01235_),
    .B(_01201_),
    .C(_01209_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _25217_ (.A(_01041_),
    .B(_01174_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand3_1 _25218_ (.A(_01236_),
    .B(_13304_),
    .C(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__inv_2 _25219_ (.A(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__a21o_1 _25220_ (.A1(_01236_),
    .A2(_01237_),
    .B1(_13304_),
    .X(_01240_));
 sky130_fd_sc_hd__o21ai_2 _25221_ (.A1(_01234_),
    .A2(_01239_),
    .B1(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__inv_2 _25222_ (.A(_01207_),
    .Y(_01242_));
 sky130_fd_sc_hd__o21ai_1 _25223_ (.A1(_01219_),
    .A2(_01242_),
    .B1(_01206_),
    .Y(_01243_));
 sky130_fd_sc_hd__a21oi_1 _25224_ (.A1(_01221_),
    .A2(_01241_),
    .B1(_01243_),
    .Y(_01245_));
 sky130_fd_sc_hd__inv_2 _25225_ (.A(_01091_),
    .Y(_01246_));
 sky130_fd_sc_hd__nand2_1 _25226_ (.A(_01041_),
    .B(_01246_),
    .Y(_01247_));
 sky130_fd_sc_hd__nand2_1 _25227_ (.A(_01092_),
    .B(_01094_),
    .Y(_01248_));
 sky130_fd_sc_hd__xor2_1 _25228_ (.A(_01093_),
    .B(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__nand3b_1 _25229_ (.A_N(_01249_),
    .B(_01037_),
    .C(_01039_),
    .Y(_01250_));
 sky130_fd_sc_hd__nand2_1 _25230_ (.A(_01247_),
    .B(_01250_),
    .Y(_01251_));
 sky130_fd_sc_hd__nand2_1 _25231_ (.A(_01251_),
    .B(_13679_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _25232_ (.A(_00161_),
    .B(_00885_),
    .Y(_01253_));
 sky130_fd_sc_hd__or2_1 _25233_ (.A(_11412_),
    .B(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__nand2_1 _25234_ (.A(_01254_),
    .B(_00529_),
    .Y(_01256_));
 sky130_fd_sc_hd__inv_2 _25235_ (.A(_01256_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2_1 _25236_ (.A(_01040_),
    .B(_01257_),
    .Y(_01258_));
 sky130_fd_sc_hd__nand3_1 _25237_ (.A(_01037_),
    .B(_01039_),
    .C(_01253_),
    .Y(_01259_));
 sky130_fd_sc_hd__nand2_1 _25238_ (.A(_01258_),
    .B(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hd__nand2_2 _25239_ (.A(_01260_),
    .B(_11421_),
    .Y(_01261_));
 sky130_fd_sc_hd__nand2_1 _25240_ (.A(_01252_),
    .B(_01261_),
    .Y(_01262_));
 sky130_fd_sc_hd__inv_2 _25241_ (.A(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__nand3_1 _25242_ (.A(_01258_),
    .B(_11426_),
    .C(_01259_),
    .Y(_01264_));
 sky130_fd_sc_hd__nand3_2 _25243_ (.A(_01041_),
    .B(_00174_),
    .C(_12221_),
    .Y(_01265_));
 sky130_fd_sc_hd__inv_2 _25244_ (.A(_01265_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand3_4 _25245_ (.A(_01261_),
    .B(_01264_),
    .C(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__or2_4 _25246_ (.A(_13679_),
    .B(_01251_),
    .X(_01269_));
 sky130_fd_sc_hd__a21boi_2 _25247_ (.A1(_01263_),
    .A2(_01268_),
    .B1_N(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__clkinvlp_2 _25248_ (.A(_01137_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2_1 _25249_ (.A(_01040_),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hd__nand2_1 _25250_ (.A(_01124_),
    .B(_01141_),
    .Y(_01273_));
 sky130_fd_sc_hd__nand3_1 _25251_ (.A(_01121_),
    .B(_01140_),
    .C(_01122_),
    .Y(_01274_));
 sky130_fd_sc_hd__nand2_1 _25252_ (.A(_01273_),
    .B(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__inv_2 _25253_ (.A(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__nand3_1 _25254_ (.A(_01037_),
    .B(_01039_),
    .C(_01276_),
    .Y(_01278_));
 sky130_fd_sc_hd__nand2_1 _25255_ (.A(_01272_),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hd__nand2_1 _25256_ (.A(_01279_),
    .B(_11482_),
    .Y(_01280_));
 sky130_fd_sc_hd__nand3_1 _25257_ (.A(_01272_),
    .B(_11484_),
    .C(_01278_),
    .Y(_01281_));
 sky130_fd_sc_hd__nand2_1 _25258_ (.A(_01280_),
    .B(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__inv_2 _25259_ (.A(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hd__nand2_1 _25260_ (.A(_01040_),
    .B(_01119_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2_1 _25261_ (.A(_01122_),
    .B(_01120_),
    .Y(_01285_));
 sky130_fd_sc_hd__xor2_1 _25262_ (.A(_01117_),
    .B(_01285_),
    .X(_01286_));
 sky130_fd_sc_hd__nand3_1 _25263_ (.A(_01037_),
    .B(_01039_),
    .C(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__nand2_1 _25264_ (.A(_01284_),
    .B(_01287_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_1 _25265_ (.A(_01289_),
    .B(_11496_),
    .Y(_01290_));
 sky130_fd_sc_hd__nand3_2 _25266_ (.A(_01284_),
    .B(_11494_),
    .C(_01287_),
    .Y(_01291_));
 sky130_fd_sc_hd__nand2_1 _25267_ (.A(_01290_),
    .B(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__inv_2 _25268_ (.A(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__nand2_1 _25269_ (.A(_01283_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__inv_2 _25270_ (.A(_01110_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2_1 _25271_ (.A(_01040_),
    .B(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__or2_1 _25272_ (.A(_01115_),
    .B(_01105_),
    .X(_01297_));
 sky130_fd_sc_hd__nand2_1 _25273_ (.A(_01297_),
    .B(_01116_),
    .Y(_01298_));
 sky130_fd_sc_hd__clkinvlp_2 _25274_ (.A(_01298_),
    .Y(_01300_));
 sky130_fd_sc_hd__nand3_1 _25275_ (.A(_01037_),
    .B(_01039_),
    .C(_01300_),
    .Y(_01301_));
 sky130_fd_sc_hd__nand2_1 _25276_ (.A(_01296_),
    .B(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__nand2_1 _25277_ (.A(_01302_),
    .B(_11105_),
    .Y(_01303_));
 sky130_fd_sc_hd__nand3_1 _25278_ (.A(_01296_),
    .B(_12261_),
    .C(_01301_),
    .Y(_01304_));
 sky130_fd_sc_hd__nand2_1 _25279_ (.A(_01303_),
    .B(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__inv_2 _25280_ (.A(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__nand2_1 _25281_ (.A(_01040_),
    .B(_01103_),
    .Y(_01307_));
 sky130_fd_sc_hd__nand2_1 _25282_ (.A(_01104_),
    .B(_01100_),
    .Y(_01308_));
 sky130_fd_sc_hd__xnor2_1 _25283_ (.A(_01096_),
    .B(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__nand3_1 _25284_ (.A(_01037_),
    .B(_01039_),
    .C(_01309_),
    .Y(_01311_));
 sky130_fd_sc_hd__nand2_1 _25285_ (.A(_01307_),
    .B(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__nand2_1 _25286_ (.A(_01312_),
    .B(_12270_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand3_1 _25287_ (.A(_01307_),
    .B(_11117_),
    .C(_01311_),
    .Y(_01314_));
 sky130_fd_sc_hd__nand2_1 _25288_ (.A(_01313_),
    .B(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__inv_2 _25289_ (.A(_01315_),
    .Y(_01316_));
 sky130_fd_sc_hd__nand2_1 _25290_ (.A(_01306_),
    .B(_01316_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_1 _25291_ (.A(_01294_),
    .B(_01317_),
    .Y(_01318_));
 sky130_fd_sc_hd__nand2_1 _25292_ (.A(_01270_),
    .B(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hd__inv_2 _25293_ (.A(_01304_),
    .Y(_01320_));
 sky130_fd_sc_hd__o21ai_1 _25294_ (.A1(_01313_),
    .A2(_01320_),
    .B1(_01303_),
    .Y(_01322_));
 sky130_fd_sc_hd__nor2_1 _25295_ (.A(_01282_),
    .B(_01292_),
    .Y(_01323_));
 sky130_fd_sc_hd__inv_2 _25296_ (.A(_01281_),
    .Y(_01324_));
 sky130_fd_sc_hd__o21ai_1 _25297_ (.A1(_01291_),
    .A2(_01324_),
    .B1(_01280_),
    .Y(_01325_));
 sky130_fd_sc_hd__a21oi_1 _25298_ (.A1(_01322_),
    .A2(_01323_),
    .B1(_01325_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_2 _25299_ (.A(_01319_),
    .B(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__nand2_1 _25300_ (.A(_01149_),
    .B(_01154_),
    .Y(_01328_));
 sky130_fd_sc_hd__nand2_1 _25301_ (.A(_01328_),
    .B(_01073_),
    .Y(_01329_));
 sky130_fd_sc_hd__nand2_1 _25302_ (.A(_01329_),
    .B(_01151_),
    .Y(_01330_));
 sky130_fd_sc_hd__nand3_1 _25303_ (.A(_01328_),
    .B(_01150_),
    .C(_01073_),
    .Y(_01331_));
 sky130_fd_sc_hd__nand2_1 _25304_ (.A(_01330_),
    .B(_01331_),
    .Y(_01333_));
 sky130_fd_sc_hd__nand2_1 _25305_ (.A(_01333_),
    .B(_01201_),
    .Y(_01334_));
 sky130_fd_sc_hd__nand2_1 _25306_ (.A(_01041_),
    .B(_01067_),
    .Y(_01335_));
 sky130_fd_sc_hd__nand2_1 _25307_ (.A(_01334_),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__nand2_1 _25308_ (.A(_01336_),
    .B(_11600_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand3_2 _25309_ (.A(_01334_),
    .B(_11603_),
    .C(_01335_),
    .Y(_01338_));
 sky130_fd_sc_hd__nand2_1 _25310_ (.A(_01337_),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__or2_1 _25311_ (.A(_01080_),
    .B(_01201_),
    .X(_01340_));
 sky130_fd_sc_hd__nand3_1 _25312_ (.A(_01223_),
    .B(_01082_),
    .C(_01078_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand3_1 _25313_ (.A(_01225_),
    .B(_01201_),
    .C(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__nand2_1 _25314_ (.A(_01340_),
    .B(_01342_),
    .Y(_01344_));
 sky130_fd_sc_hd__nand2_1 _25315_ (.A(_01344_),
    .B(_11586_),
    .Y(_01345_));
 sky130_fd_sc_hd__nand3_1 _25316_ (.A(_01340_),
    .B(_01342_),
    .C(_11588_),
    .Y(_01346_));
 sky130_fd_sc_hd__nand2_2 _25317_ (.A(_01345_),
    .B(_01346_),
    .Y(_01347_));
 sky130_fd_sc_hd__nor2_1 _25318_ (.A(_01339_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hd__or2_1 _25319_ (.A(_01154_),
    .B(_01149_),
    .X(_01349_));
 sky130_fd_sc_hd__nand3_1 _25320_ (.A(_01201_),
    .B(_01328_),
    .C(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hd__nand2_1 _25321_ (.A(_01041_),
    .B(_01072_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2_1 _25322_ (.A(_01350_),
    .B(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__nand2_1 _25323_ (.A(_01352_),
    .B(_11614_),
    .Y(_01353_));
 sky130_fd_sc_hd__nand3_1 _25324_ (.A(_01350_),
    .B(_11616_),
    .C(_01351_),
    .Y(_01355_));
 sky130_fd_sc_hd__nand2_1 _25325_ (.A(_01353_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__nand2_1 _25326_ (.A(_01135_),
    .B(_01142_),
    .Y(_01357_));
 sky130_fd_sc_hd__nand2_1 _25327_ (.A(_01273_),
    .B(_01139_),
    .Y(_01358_));
 sky130_fd_sc_hd__xor2_1 _25328_ (.A(_01357_),
    .B(_01358_),
    .X(_01359_));
 sky130_fd_sc_hd__nand2_1 _25329_ (.A(_01359_),
    .B(_01201_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _25330_ (.A(_01041_),
    .B(_01133_),
    .Y(_01361_));
 sky130_fd_sc_hd__a21o_1 _25331_ (.A1(_01360_),
    .A2(_01361_),
    .B1(_08951_),
    .X(_01362_));
 sky130_fd_sc_hd__nand3_1 _25332_ (.A(_01360_),
    .B(_08951_),
    .C(_01361_),
    .Y(_01363_));
 sky130_fd_sc_hd__nand2_1 _25333_ (.A(_01362_),
    .B(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_1 _25334_ (.A(_01356_),
    .B(_01364_),
    .Y(_01366_));
 sky130_fd_sc_hd__and2_1 _25335_ (.A(_01348_),
    .B(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__nand2_1 _25336_ (.A(_01327_),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__inv_2 _25337_ (.A(_01355_),
    .Y(_01369_));
 sky130_fd_sc_hd__o21ai_1 _25338_ (.A1(_01363_),
    .A2(_01369_),
    .B1(_01353_),
    .Y(_01370_));
 sky130_fd_sc_hd__inv_2 _25339_ (.A(_01346_),
    .Y(_01371_));
 sky130_fd_sc_hd__o21ai_1 _25340_ (.A1(_01338_),
    .A2(_01371_),
    .B1(_01345_),
    .Y(_01372_));
 sky130_fd_sc_hd__a21oi_1 _25341_ (.A1(_01348_),
    .A2(_01370_),
    .B1(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__nand2_2 _25342_ (.A(_01368_),
    .B(_01373_),
    .Y(_01374_));
 sky130_fd_sc_hd__nand2_1 _25343_ (.A(_01231_),
    .B(_01232_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand2_1 _25344_ (.A(_01375_),
    .B(_11185_),
    .Y(_01377_));
 sky130_fd_sc_hd__nand2_1 _25345_ (.A(_01377_),
    .B(_01234_),
    .Y(_01378_));
 sky130_fd_sc_hd__nand2_1 _25346_ (.A(_01240_),
    .B(_01238_),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_1 _25347_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__nand3_1 _25348_ (.A(_01374_),
    .B(_01221_),
    .C(_01380_),
    .Y(_01381_));
 sky130_fd_sc_hd__nand2_2 _25349_ (.A(_01245_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand2_1 _25350_ (.A(_00918_),
    .B(_00919_),
    .Y(_01383_));
 sky130_fd_sc_hd__inv_2 _25351_ (.A(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__or2_1 _25352_ (.A(_01384_),
    .B(_00831_),
    .X(_01385_));
 sky130_fd_sc_hd__nand2_1 _25353_ (.A(_00831_),
    .B(_01384_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand2_1 _25354_ (.A(_01385_),
    .B(_01386_),
    .Y(_01388_));
 sky130_fd_sc_hd__inv_2 _25355_ (.A(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__nand2_1 _25356_ (.A(_01389_),
    .B(_11199_),
    .Y(_01390_));
 sky130_fd_sc_hd__nand2_1 _25357_ (.A(_01388_),
    .B(_13461_),
    .Y(_01391_));
 sky130_fd_sc_hd__nand2_1 _25358_ (.A(_01390_),
    .B(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__inv_2 _25359_ (.A(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__nand2_1 _25360_ (.A(_01191_),
    .B(_00803_),
    .Y(_01394_));
 sky130_fd_sc_hd__inv_2 _25361_ (.A(_00792_),
    .Y(_01395_));
 sky130_fd_sc_hd__nand2_1 _25362_ (.A(_01394_),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hd__nand3_1 _25363_ (.A(_01191_),
    .B(_00792_),
    .C(_00803_),
    .Y(_01397_));
 sky130_fd_sc_hd__nand2_1 _25364_ (.A(_01396_),
    .B(_01397_),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2_1 _25365_ (.A(_01399_),
    .B(_12894_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand3_1 _25366_ (.A(_01396_),
    .B(_11754_),
    .C(_01397_),
    .Y(_01401_));
 sky130_fd_sc_hd__nand3_1 _25367_ (.A(_01198_),
    .B(_01400_),
    .C(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__inv_2 _25368_ (.A(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__nand3_1 _25369_ (.A(_01159_),
    .B(_01181_),
    .C(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__inv_2 _25370_ (.A(_01400_),
    .Y(_01405_));
 sky130_fd_sc_hd__o21ai_1 _25371_ (.A1(_01195_),
    .A2(_01405_),
    .B1(_01401_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _25372_ (.A(_01184_),
    .B(_01402_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _25373_ (.A(_01406_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__nand2_1 _25374_ (.A(_01404_),
    .B(_01408_),
    .Y(_01410_));
 sky130_fd_sc_hd__or2_1 _25375_ (.A(_01393_),
    .B(_01410_),
    .X(_01411_));
 sky130_fd_sc_hd__buf_6 _25376_ (.A(_01201_),
    .X(_01412_));
 sky130_fd_sc_hd__nand2_1 _25377_ (.A(_01410_),
    .B(_01393_),
    .Y(_01413_));
 sky130_fd_sc_hd__nand3_1 _25378_ (.A(_01411_),
    .B(_01412_),
    .C(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__nand2_1 _25379_ (.A(\div1i.quot[2] ),
    .B(_01389_),
    .Y(_01415_));
 sky130_fd_sc_hd__nand2_1 _25380_ (.A(_01414_),
    .B(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__xor2_2 _25381_ (.A(_06754_),
    .B(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__nand2_1 _25382_ (.A(_01400_),
    .B(_01401_),
    .Y(_01418_));
 sky130_fd_sc_hd__nand2_1 _25383_ (.A(_01199_),
    .B(_01195_),
    .Y(_01419_));
 sky130_fd_sc_hd__xor2_1 _25384_ (.A(_01418_),
    .B(_01419_),
    .X(_01421_));
 sky130_fd_sc_hd__nand2_1 _25385_ (.A(_01421_),
    .B(_01412_),
    .Y(_01422_));
 sky130_fd_sc_hd__nand2_1 _25386_ (.A(\div1i.quot[2] ),
    .B(_01399_),
    .Y(_01423_));
 sky130_fd_sc_hd__nand2_1 _25387_ (.A(_01422_),
    .B(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__nand2_1 _25388_ (.A(_01424_),
    .B(_11838_),
    .Y(_01425_));
 sky130_fd_sc_hd__nand3_1 _25389_ (.A(_01422_),
    .B(_11840_),
    .C(_01423_),
    .Y(_01426_));
 sky130_fd_sc_hd__nand2_1 _25390_ (.A(_01425_),
    .B(_01426_),
    .Y(_01427_));
 sky130_fd_sc_hd__nor2_1 _25391_ (.A(_01417_),
    .B(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__nand2_2 _25392_ (.A(_01382_),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand2_1 _25393_ (.A(_01416_),
    .B(_13502_),
    .Y(_01430_));
 sky130_fd_sc_hd__o21a_1 _25394_ (.A1(_01426_),
    .A2(_01417_),
    .B1(_01430_),
    .X(_01432_));
 sky130_fd_sc_hd__nand2_1 _25395_ (.A(_01429_),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_1 _25396_ (.A(_00831_),
    .B(_00921_),
    .Y(_01434_));
 sky130_fd_sc_hd__inv_2 _25397_ (.A(_00924_),
    .Y(_01435_));
 sky130_fd_sc_hd__a21o_1 _25398_ (.A1(_01434_),
    .A2(_01435_),
    .B1(_00902_),
    .X(_01436_));
 sky130_fd_sc_hd__nand3_1 _25399_ (.A(_01434_),
    .B(_00902_),
    .C(_01435_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_1 _25400_ (.A(_01436_),
    .B(_01437_),
    .Y(_01438_));
 sky130_fd_sc_hd__inv_2 _25401_ (.A(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2_1 _25402_ (.A(_01439_),
    .B(_11797_),
    .Y(_01440_));
 sky130_fd_sc_hd__nand2_1 _25403_ (.A(_01438_),
    .B(_12939_),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_1 _25404_ (.A(_01440_),
    .B(_01441_),
    .Y(_01443_));
 sky130_fd_sc_hd__inv_2 _25405_ (.A(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__nand2_1 _25406_ (.A(_01386_),
    .B(_00919_),
    .Y(_01445_));
 sky130_fd_sc_hd__xor2_2 _25407_ (.A(_00911_),
    .B(_01445_),
    .X(_01446_));
 sky130_fd_sc_hd__inv_2 _25408_ (.A(_01446_),
    .Y(_01447_));
 sky130_fd_sc_hd__nand2_1 _25409_ (.A(_01447_),
    .B(_11774_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _25410_ (.A(_01446_),
    .B(_12914_),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_1 _25411_ (.A(_01448_),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__or2_1 _25412_ (.A(_01392_),
    .B(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__inv_4 _25413_ (.A(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__nand2_1 _25414_ (.A(_01410_),
    .B(_01452_),
    .Y(_01454_));
 sky130_fd_sc_hd__inv_2 _25415_ (.A(_01390_),
    .Y(_01455_));
 sky130_fd_sc_hd__a21boi_1 _25416_ (.A1(_01455_),
    .A2(_01449_),
    .B1_N(_01448_),
    .Y(_01456_));
 sky130_fd_sc_hd__nand2_1 _25417_ (.A(_01454_),
    .B(_01456_),
    .Y(_01457_));
 sky130_fd_sc_hd__or2_1 _25418_ (.A(_01444_),
    .B(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__nand2_1 _25419_ (.A(_01457_),
    .B(_01444_),
    .Y(_01459_));
 sky130_fd_sc_hd__nand3_1 _25420_ (.A(_01458_),
    .B(_01412_),
    .C(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _25421_ (.A(\div1i.quot[2] ),
    .B(_01439_),
    .Y(_01461_));
 sky130_fd_sc_hd__nand2_1 _25422_ (.A(_01460_),
    .B(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__xor2_2 _25423_ (.A(_11811_),
    .B(_01462_),
    .X(_01463_));
 sky130_fd_sc_hd__nand2_1 _25424_ (.A(_01413_),
    .B(_01390_),
    .Y(_01465_));
 sky130_fd_sc_hd__xor2_1 _25425_ (.A(_01450_),
    .B(_01465_),
    .X(_01466_));
 sky130_fd_sc_hd__nand2_1 _25426_ (.A(_01466_),
    .B(_01412_),
    .Y(_01467_));
 sky130_fd_sc_hd__nand2_1 _25427_ (.A(\div1i.quot[2] ),
    .B(_01446_),
    .Y(_01468_));
 sky130_fd_sc_hd__nand2_1 _25428_ (.A(_01467_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hd__or2_1 _25429_ (.A(_13537_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__nand2_1 _25430_ (.A(_01469_),
    .B(_13537_),
    .Y(_01471_));
 sky130_fd_sc_hd__nand2_1 _25431_ (.A(_01470_),
    .B(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__nor2_1 _25432_ (.A(_01463_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hd__nand2_1 _25433_ (.A(_01433_),
    .B(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__nand2_1 _25434_ (.A(_01462_),
    .B(_11808_),
    .Y(_01476_));
 sky130_fd_sc_hd__o21a_1 _25435_ (.A1(_01470_),
    .A2(_01463_),
    .B1(_01476_),
    .X(_01477_));
 sky130_fd_sc_hd__nand2_2 _25436_ (.A(_01474_),
    .B(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hd__nand2_1 _25437_ (.A(_00973_),
    .B(_00974_),
    .Y(_01479_));
 sky130_fd_sc_hd__nand2b_1 _25438_ (.A_N(_00928_),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nand2b_1 _25439_ (.A_N(_01479_),
    .B(_00928_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand2_1 _25440_ (.A(_01480_),
    .B(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__or2_1 _25441_ (.A(_14113_),
    .B(_01482_),
    .X(_01483_));
 sky130_fd_sc_hd__nand2_1 _25442_ (.A(_01482_),
    .B(_14113_),
    .Y(_01484_));
 sky130_fd_sc_hd__nand2_1 _25443_ (.A(_01483_),
    .B(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__inv_4 _25444_ (.A(_01485_),
    .Y(_01487_));
 sky130_fd_sc_hd__nand2_1 _25445_ (.A(_01436_),
    .B(_00901_),
    .Y(_01488_));
 sky130_fd_sc_hd__inv_2 _25446_ (.A(_00892_),
    .Y(_01489_));
 sky130_fd_sc_hd__nand2_1 _25447_ (.A(_01488_),
    .B(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hd__nand3_1 _25448_ (.A(_01436_),
    .B(_00892_),
    .C(_00901_),
    .Y(_01491_));
 sky130_fd_sc_hd__nand2_1 _25449_ (.A(_01490_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2_1 _25450_ (.A(_01492_),
    .B(_12992_),
    .Y(_01493_));
 sky130_fd_sc_hd__nand3_2 _25451_ (.A(_01490_),
    .B(_11858_),
    .C(_01491_),
    .Y(_01494_));
 sky130_fd_sc_hd__nand3_1 _25452_ (.A(_01444_),
    .B(_01493_),
    .C(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__inv_2 _25453_ (.A(_01495_),
    .Y(_01496_));
 sky130_fd_sc_hd__nand3_1 _25454_ (.A(_01410_),
    .B(_01452_),
    .C(_01496_),
    .Y(_01498_));
 sky130_fd_sc_hd__inv_2 _25455_ (.A(_01440_),
    .Y(_01499_));
 sky130_fd_sc_hd__inv_2 _25456_ (.A(_01494_),
    .Y(_01500_));
 sky130_fd_sc_hd__a21o_1 _25457_ (.A1(_01493_),
    .A2(_01499_),
    .B1(_01500_),
    .X(_01501_));
 sky130_fd_sc_hd__nor2_1 _25458_ (.A(_01456_),
    .B(_01495_),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _25459_ (.A(_01501_),
    .B(_01502_),
    .Y(_01503_));
 sky130_fd_sc_hd__nand2_1 _25460_ (.A(_01498_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__or2_1 _25461_ (.A(_01487_),
    .B(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__nand2_1 _25462_ (.A(_01504_),
    .B(_01487_),
    .Y(_01506_));
 sky130_fd_sc_hd__nand2_1 _25463_ (.A(_01505_),
    .B(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__nand2_1 _25464_ (.A(_01507_),
    .B(_01412_),
    .Y(_01509_));
 sky130_fd_sc_hd__nand2_1 _25465_ (.A(\div1i.quot[2] ),
    .B(_01482_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand2_1 _25466_ (.A(_01509_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__nand2_1 _25467_ (.A(_01511_),
    .B(_08020_),
    .Y(_01512_));
 sky130_fd_sc_hd__nand3_1 _25468_ (.A(_01509_),
    .B(_13022_),
    .C(_01510_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_1 _25469_ (.A(_01512_),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__inv_2 _25470_ (.A(_01514_),
    .Y(_01515_));
 sky130_fd_sc_hd__nand2_1 _25471_ (.A(_01493_),
    .B(_01494_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand2_1 _25472_ (.A(_01459_),
    .B(_01440_),
    .Y(_01517_));
 sky130_fd_sc_hd__xor2_1 _25473_ (.A(_01516_),
    .B(_01517_),
    .X(_01518_));
 sky130_fd_sc_hd__nand2_1 _25474_ (.A(_01518_),
    .B(_01412_),
    .Y(_01520_));
 sky130_fd_sc_hd__nand2_1 _25475_ (.A(_01492_),
    .B(\div1i.quot[2] ),
    .Y(_01521_));
 sky130_fd_sc_hd__nand2_1 _25476_ (.A(_01520_),
    .B(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__nand2_1 _25477_ (.A(_01522_),
    .B(_11896_),
    .Y(_01523_));
 sky130_fd_sc_hd__nand3_2 _25478_ (.A(_01520_),
    .B(_11899_),
    .C(_01521_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand3_1 _25479_ (.A(_01515_),
    .B(_01523_),
    .C(_01524_),
    .Y(_01525_));
 sky130_fd_sc_hd__nand2_1 _25480_ (.A(_01506_),
    .B(_01483_),
    .Y(_01526_));
 sky130_fd_sc_hd__nand2_1 _25481_ (.A(_01481_),
    .B(_00974_),
    .Y(_01527_));
 sky130_fd_sc_hd__or2_1 _25482_ (.A(_00965_),
    .B(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__nand2_1 _25483_ (.A(_01527_),
    .B(_00965_),
    .Y(_01529_));
 sky130_fd_sc_hd__nand2_1 _25484_ (.A(_01528_),
    .B(_01529_),
    .Y(_01531_));
 sky130_fd_sc_hd__nand2_1 _25485_ (.A(_01531_),
    .B(_13042_),
    .Y(_01532_));
 sky130_fd_sc_hd__nand3_1 _25486_ (.A(_01528_),
    .B(_12495_),
    .C(_01529_),
    .Y(_01533_));
 sky130_fd_sc_hd__nand2_1 _25487_ (.A(_01532_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__inv_2 _25488_ (.A(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__nand2_1 _25489_ (.A(_01526_),
    .B(_01535_),
    .Y(_01536_));
 sky130_fd_sc_hd__nand3_1 _25490_ (.A(_01506_),
    .B(_01534_),
    .C(_01483_),
    .Y(_01537_));
 sky130_fd_sc_hd__nand2_1 _25491_ (.A(_01536_),
    .B(_01537_),
    .Y(_01538_));
 sky130_fd_sc_hd__nand2_1 _25492_ (.A(_01538_),
    .B(_01412_),
    .Y(_01539_));
 sky130_fd_sc_hd__nand2_1 _25493_ (.A(_01531_),
    .B(\div1i.quot[2] ),
    .Y(_01540_));
 sky130_fd_sc_hd__nand2_1 _25494_ (.A(_01539_),
    .B(_01540_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2_1 _25495_ (.A(_01542_),
    .B(_12506_),
    .Y(_01543_));
 sky130_fd_sc_hd__nand3_1 _25496_ (.A(_01539_),
    .B(_11376_),
    .C(_01540_),
    .Y(_01544_));
 sky130_fd_sc_hd__nand2_1 _25497_ (.A(_01543_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__inv_2 _25498_ (.A(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_1 _25499_ (.A(_01535_),
    .B(_01487_),
    .Y(_01547_));
 sky130_fd_sc_hd__inv_2 _25500_ (.A(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__nand2_1 _25501_ (.A(_01504_),
    .B(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__o21a_1 _25502_ (.A1(_01483_),
    .A2(_01534_),
    .B1(_01533_),
    .X(_01550_));
 sky130_fd_sc_hd__nand2_1 _25503_ (.A(_01549_),
    .B(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__a41o_1 _25504_ (.A1(_00928_),
    .A2(_00965_),
    .A3(_00974_),
    .A4(_00973_),
    .B1(_01026_),
    .X(_01553_));
 sky130_fd_sc_hd__or2_1 _25505_ (.A(_00995_),
    .B(_01553_),
    .X(_01554_));
 sky130_fd_sc_hd__nand2_1 _25506_ (.A(_01553_),
    .B(_00995_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _25507_ (.A(_01554_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__inv_2 _25508_ (.A(_01556_),
    .Y(_01557_));
 sky130_fd_sc_hd__nand2_1 _25509_ (.A(_01557_),
    .B(_11935_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_1 _25510_ (.A(_01556_),
    .B(_13633_),
    .Y(_01559_));
 sky130_fd_sc_hd__nand2_1 _25511_ (.A(_01558_),
    .B(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hd__clkinvlp_2 _25512_ (.A(_01560_),
    .Y(_01561_));
 sky130_fd_sc_hd__nand2_1 _25513_ (.A(_01551_),
    .B(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__nand3_1 _25514_ (.A(_01549_),
    .B(_01560_),
    .C(_01550_),
    .Y(_01564_));
 sky130_fd_sc_hd__nand3_1 _25515_ (.A(_01562_),
    .B(_01564_),
    .C(_01412_),
    .Y(_01565_));
 sky130_fd_sc_hd__nand2_1 _25516_ (.A(_01557_),
    .B(\div1i.quot[2] ),
    .Y(_01566_));
 sky130_fd_sc_hd__nand2_1 _25517_ (.A(_01565_),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__nand2_1 _25518_ (.A(_01567_),
    .B(_11946_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand3_1 _25519_ (.A(_01565_),
    .B(_11948_),
    .C(_01566_),
    .Y(_01569_));
 sky130_fd_sc_hd__nand2_2 _25520_ (.A(_01568_),
    .B(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hd__inv_2 _25521_ (.A(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__nand2_1 _25522_ (.A(_01546_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__nor2_2 _25523_ (.A(_01572_),
    .B(_01525_),
    .Y(_01573_));
 sky130_fd_sc_hd__nand2_4 _25524_ (.A(_01478_),
    .B(_01573_),
    .Y(_01575_));
 sky130_fd_sc_hd__o21ai_1 _25525_ (.A1(_01524_),
    .A2(_01514_),
    .B1(_01513_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _25526_ (.A(_01570_),
    .B(_01545_),
    .Y(_01577_));
 sky130_fd_sc_hd__o21ai_1 _25527_ (.A1(_01544_),
    .A2(_01570_),
    .B1(_01568_),
    .Y(_01578_));
 sky130_fd_sc_hd__a21oi_2 _25528_ (.A1(_01576_),
    .A2(_01577_),
    .B1(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__nand2_2 _25529_ (.A(_01575_),
    .B(_01579_),
    .Y(_01580_));
 sky130_fd_sc_hd__nand2_1 _25530_ (.A(_01555_),
    .B(_00993_),
    .Y(_01581_));
 sky130_fd_sc_hd__xor2_1 _25531_ (.A(_01020_),
    .B(_01581_),
    .X(_01582_));
 sky130_fd_sc_hd__nand3_1 _25532_ (.A(_01562_),
    .B(_01412_),
    .C(_01558_),
    .Y(_01583_));
 sky130_fd_sc_hd__xnor2_2 _25533_ (.A(_01582_),
    .B(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__nand2_4 _25534_ (.A(_01580_),
    .B(_01584_),
    .Y(_01586_));
 sky130_fd_sc_hd__clkinvlp_2 _25535_ (.A(_01584_),
    .Y(_01587_));
 sky130_fd_sc_hd__nand3_4 _25536_ (.A(_01575_),
    .B(_01579_),
    .C(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__nand2_8 _25537_ (.A(_01586_),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__buf_8 _25538_ (.A(_01589_),
    .X(_01590_));
 sky130_fd_sc_hd__buf_8 _25539_ (.A(net233),
    .X(\div1i.quot[1] ));
 sky130_fd_sc_hd__nor2_1 _25540_ (.A(_00161_),
    .B(_01412_),
    .Y(_01591_));
 sky130_fd_sc_hd__or2_1 _25541_ (.A(_11412_),
    .B(_01591_),
    .X(_01592_));
 sky130_fd_sc_hd__nand2_1 _25542_ (.A(_01592_),
    .B(_01265_),
    .Y(_01593_));
 sky130_fd_sc_hd__inv_2 _25543_ (.A(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__nand2_1 _25544_ (.A(_01589_),
    .B(_01594_),
    .Y(_01596_));
 sky130_fd_sc_hd__nand3_1 _25545_ (.A(_01586_),
    .B(_01588_),
    .C(_01591_),
    .Y(_01597_));
 sky130_fd_sc_hd__nand2_1 _25546_ (.A(_01596_),
    .B(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_2 _25547_ (.A(_01598_),
    .B(_11421_),
    .Y(_01599_));
 sky130_fd_sc_hd__nand3_1 _25548_ (.A(_01596_),
    .B(_11426_),
    .C(_01597_),
    .Y(_01600_));
 sky130_fd_sc_hd__nand3_2 _25549_ (.A(_01589_),
    .B(_00174_),
    .C(_12221_),
    .Y(_01601_));
 sky130_fd_sc_hd__inv_2 _25550_ (.A(_01601_),
    .Y(_01602_));
 sky130_fd_sc_hd__nand3_2 _25551_ (.A(_01599_),
    .B(_01600_),
    .C(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__inv_2 _25552_ (.A(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_1 _25553_ (.A(_01261_),
    .B(_01264_),
    .Y(_01605_));
 sky130_fd_sc_hd__nand2_1 _25554_ (.A(_01605_),
    .B(_01265_),
    .Y(_01607_));
 sky130_fd_sc_hd__nand2_1 _25555_ (.A(_01607_),
    .B(_01268_),
    .Y(_01608_));
 sky130_fd_sc_hd__inv_2 _25556_ (.A(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_1 _25557_ (.A(_01590_),
    .B(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__o21ai_2 _25558_ (.A1(_00161_),
    .A2(\div1i.quot[2] ),
    .B1(_00174_),
    .Y(_01611_));
 sky130_fd_sc_hd__nand2_1 _25559_ (.A(_01608_),
    .B(_12030_),
    .Y(_01612_));
 sky130_fd_sc_hd__nand3_1 _25560_ (.A(_01607_),
    .B(_12035_),
    .C(_01268_),
    .Y(_01613_));
 sky130_fd_sc_hd__nand2_1 _25561_ (.A(_01612_),
    .B(_01613_),
    .Y(_01614_));
 sky130_fd_sc_hd__xor2_1 _25562_ (.A(_01611_),
    .B(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__nand3b_1 _25563_ (.A_N(_01615_),
    .B(_01586_),
    .C(_01588_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _25564_ (.A(_01610_),
    .B(_01616_),
    .Y(_01618_));
 sky130_fd_sc_hd__nand2_1 _25565_ (.A(_01618_),
    .B(_13679_),
    .Y(_01619_));
 sky130_fd_sc_hd__nand3_2 _25566_ (.A(_01610_),
    .B(_01616_),
    .C(_11799_),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_2 _25567_ (.A(_01619_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__inv_4 _25568_ (.A(_01621_),
    .Y(_01622_));
 sky130_fd_sc_hd__nand2_1 _25569_ (.A(_01604_),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__inv_2 _25570_ (.A(_01599_),
    .Y(_01624_));
 sky130_fd_sc_hd__a21boi_2 _25571_ (.A1(_01624_),
    .A2(_01620_),
    .B1_N(_01619_),
    .Y(_01625_));
 sky130_fd_sc_hd__nand2_2 _25572_ (.A(_01625_),
    .B(_01623_),
    .Y(_01626_));
 sky130_fd_sc_hd__nand2_1 _25573_ (.A(_01263_),
    .B(_01268_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _25574_ (.A(_01305_),
    .B(_01315_),
    .Y(_01629_));
 sky130_fd_sc_hd__a31o_1 _25575_ (.A1(_01627_),
    .A2(_01629_),
    .A3(_01269_),
    .B1(_01322_),
    .X(_01630_));
 sky130_fd_sc_hd__or2_1 _25576_ (.A(_01293_),
    .B(_01630_),
    .X(_01631_));
 sky130_fd_sc_hd__nand2_1 _25577_ (.A(_01630_),
    .B(_01293_),
    .Y(_01632_));
 sky130_fd_sc_hd__nand2_1 _25578_ (.A(_01631_),
    .B(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__inv_2 _25579_ (.A(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__nand2_1 _25580_ (.A(_01590_),
    .B(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__nand2_1 _25581_ (.A(_01633_),
    .B(_12085_),
    .Y(_01636_));
 sky130_fd_sc_hd__nand3_1 _25582_ (.A(_01631_),
    .B(_12087_),
    .C(_01632_),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2_1 _25583_ (.A(_01636_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__inv_2 _25584_ (.A(_01638_),
    .Y(_01640_));
 sky130_fd_sc_hd__nand2_1 _25585_ (.A(_01270_),
    .B(_01316_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_1 _25586_ (.A(_01627_),
    .B(_01269_),
    .Y(_01642_));
 sky130_fd_sc_hd__nand2_1 _25587_ (.A(_01642_),
    .B(_01315_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand2_1 _25588_ (.A(_01641_),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__nand2_1 _25589_ (.A(_01644_),
    .B(_12056_),
    .Y(_01645_));
 sky130_fd_sc_hd__nand3_1 _25590_ (.A(_01641_),
    .B(_12058_),
    .C(_01643_),
    .Y(_01646_));
 sky130_fd_sc_hd__nand2_1 _25591_ (.A(_01645_),
    .B(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__inv_2 _25592_ (.A(_01647_),
    .Y(_01648_));
 sky130_fd_sc_hd__inv_2 _25593_ (.A(_01613_),
    .Y(_01649_));
 sky130_fd_sc_hd__a21o_1 _25594_ (.A1(_01612_),
    .A2(_01611_),
    .B1(_01649_),
    .X(_01651_));
 sky130_fd_sc_hd__nand2_1 _25595_ (.A(_01269_),
    .B(_01252_),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_1 _25596_ (.A(_01268_),
    .B(_01261_),
    .Y(_01653_));
 sky130_fd_sc_hd__xor2_1 _25597_ (.A(_01652_),
    .B(_01653_),
    .X(_01654_));
 sky130_fd_sc_hd__nand2_1 _25598_ (.A(_01654_),
    .B(_12043_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_1 _25599_ (.A(_01651_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__inv_2 _25600_ (.A(_01654_),
    .Y(_01657_));
 sky130_fd_sc_hd__nand2_1 _25601_ (.A(_01657_),
    .B(_12047_),
    .Y(_01658_));
 sky130_fd_sc_hd__nand2_1 _25602_ (.A(_01656_),
    .B(_01658_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_1 _25603_ (.A(_01648_),
    .B(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__nand2_1 _25604_ (.A(_01660_),
    .B(_01646_),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_1 _25605_ (.A(_01641_),
    .B(_01313_),
    .Y(_01663_));
 sky130_fd_sc_hd__xor2_1 _25606_ (.A(_01305_),
    .B(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__nand2_1 _25607_ (.A(_01664_),
    .B(_13182_),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_1 _25608_ (.A(_01662_),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__inv_2 _25609_ (.A(_01664_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _25610_ (.A(_01667_),
    .B(_08176_),
    .Y(_01668_));
 sky130_fd_sc_hd__nand2_1 _25611_ (.A(_01666_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__or2_1 _25612_ (.A(_01640_),
    .B(_01669_),
    .X(_01670_));
 sky130_fd_sc_hd__nand2_1 _25613_ (.A(_01669_),
    .B(_01640_),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2_1 _25614_ (.A(_01670_),
    .B(_01671_),
    .Y(_01673_));
 sky130_fd_sc_hd__inv_2 _25615_ (.A(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__nand3_1 _25616_ (.A(net129),
    .B(net119),
    .C(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__nand2_1 _25617_ (.A(_01635_),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__nand2_1 _25618_ (.A(_01676_),
    .B(_11482_),
    .Y(_01677_));
 sky130_fd_sc_hd__nand3_1 _25619_ (.A(_01635_),
    .B(_11484_),
    .C(_01675_),
    .Y(_01678_));
 sky130_fd_sc_hd__nand2_1 _25620_ (.A(_01677_),
    .B(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__inv_2 _25621_ (.A(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__nand2_1 _25622_ (.A(_01590_),
    .B(_01667_),
    .Y(_01681_));
 sky130_fd_sc_hd__nand2_1 _25623_ (.A(_01668_),
    .B(_01665_),
    .Y(_01682_));
 sky130_fd_sc_hd__xnor2_1 _25624_ (.A(_01662_),
    .B(_01682_),
    .Y(_01684_));
 sky130_fd_sc_hd__nand3_1 _25625_ (.A(net129),
    .B(_01588_),
    .C(_01684_),
    .Y(_01685_));
 sky130_fd_sc_hd__nand2_1 _25626_ (.A(_01681_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__nand2_2 _25627_ (.A(_01686_),
    .B(_11494_),
    .Y(_01687_));
 sky130_fd_sc_hd__nand3_1 _25628_ (.A(_01681_),
    .B(_11496_),
    .C(_01685_),
    .Y(_01688_));
 sky130_fd_sc_hd__nand2_2 _25629_ (.A(_01687_),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__inv_2 _25630_ (.A(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__nand2_1 _25631_ (.A(_01680_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hd__inv_2 _25632_ (.A(_01644_),
    .Y(_01692_));
 sky130_fd_sc_hd__nand2_1 _25633_ (.A(_01590_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__or2_1 _25634_ (.A(_01659_),
    .B(_01648_),
    .X(_01695_));
 sky130_fd_sc_hd__nand2_1 _25635_ (.A(_01695_),
    .B(_01660_),
    .Y(_01696_));
 sky130_fd_sc_hd__clkinvlp_2 _25636_ (.A(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__nand3_1 _25637_ (.A(_01586_),
    .B(net119),
    .C(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hd__nand2_1 _25638_ (.A(_01693_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_2 _25639_ (.A(_01699_),
    .B(_11105_),
    .Y(_01700_));
 sky130_fd_sc_hd__nand3_2 _25640_ (.A(_01693_),
    .B(_12261_),
    .C(_01698_),
    .Y(_01701_));
 sky130_fd_sc_hd__nand2_2 _25641_ (.A(_01700_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__inv_2 _25642_ (.A(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__nand2_1 _25643_ (.A(_01589_),
    .B(_01657_),
    .Y(_01704_));
 sky130_fd_sc_hd__nand2_1 _25644_ (.A(_01658_),
    .B(_01655_),
    .Y(_01706_));
 sky130_fd_sc_hd__xnor2_1 _25645_ (.A(_01651_),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__nand3_1 _25646_ (.A(_01586_),
    .B(_01588_),
    .C(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand2_1 _25647_ (.A(_01704_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__nand2_2 _25648_ (.A(_01709_),
    .B(_12270_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand3_1 _25649_ (.A(_01704_),
    .B(_11117_),
    .C(_01708_),
    .Y(_01711_));
 sky130_fd_sc_hd__nand2_1 _25650_ (.A(_01710_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__inv_2 _25651_ (.A(_01712_),
    .Y(_01713_));
 sky130_fd_sc_hd__nand2_2 _25652_ (.A(_01703_),
    .B(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__nor2_1 _25653_ (.A(_01691_),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__nand2_1 _25654_ (.A(_01626_),
    .B(_01715_),
    .Y(_01717_));
 sky130_fd_sc_hd__inv_2 _25655_ (.A(_01701_),
    .Y(_01718_));
 sky130_fd_sc_hd__o21ai_2 _25656_ (.A1(_01710_),
    .A2(_01718_),
    .B1(_01700_),
    .Y(_01719_));
 sky130_fd_sc_hd__nor2_1 _25657_ (.A(_01679_),
    .B(_01689_),
    .Y(_01720_));
 sky130_fd_sc_hd__inv_2 _25658_ (.A(_01678_),
    .Y(_01721_));
 sky130_fd_sc_hd__o21ai_1 _25659_ (.A1(_01687_),
    .A2(_01721_),
    .B1(_01677_),
    .Y(_01722_));
 sky130_fd_sc_hd__a21oi_1 _25660_ (.A1(_01719_),
    .A2(_01720_),
    .B1(_01722_),
    .Y(_01723_));
 sky130_fd_sc_hd__nand2_2 _25661_ (.A(_01717_),
    .B(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__inv_6 _25662_ (.A(_01589_),
    .Y(_01725_));
 sky130_fd_sc_hd__nand2_1 _25663_ (.A(_01632_),
    .B(_01291_),
    .Y(_01726_));
 sky130_fd_sc_hd__nand2_1 _25664_ (.A(_01726_),
    .B(_01283_),
    .Y(_01728_));
 sky130_fd_sc_hd__nand3_1 _25665_ (.A(_01632_),
    .B(_01282_),
    .C(_01291_),
    .Y(_01729_));
 sky130_fd_sc_hd__nand2_1 _25666_ (.A(_01728_),
    .B(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hd__o21ai_1 _25667_ (.A1(_13197_),
    .A2(_01730_),
    .B1(_01637_),
    .Y(_01731_));
 sky130_fd_sc_hd__inv_2 _25668_ (.A(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__nand2_1 _25669_ (.A(_01671_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand2_1 _25670_ (.A(_01730_),
    .B(_13197_),
    .Y(_01734_));
 sky130_fd_sc_hd__inv_2 _25671_ (.A(_01364_),
    .Y(_01735_));
 sky130_fd_sc_hd__or2_1 _25672_ (.A(_01735_),
    .B(_01327_),
    .X(_01736_));
 sky130_fd_sc_hd__nand2_1 _25673_ (.A(_01327_),
    .B(_01735_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_1 _25674_ (.A(_01736_),
    .B(_01737_),
    .Y(_01739_));
 sky130_fd_sc_hd__nand2_1 _25675_ (.A(_01739_),
    .B(_12101_),
    .Y(_01740_));
 sky130_fd_sc_hd__nand3_2 _25676_ (.A(_01736_),
    .B(_12008_),
    .C(_01737_),
    .Y(_01741_));
 sky130_fd_sc_hd__nand2_1 _25677_ (.A(_01740_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__inv_2 _25678_ (.A(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand3_1 _25679_ (.A(_01733_),
    .B(_01734_),
    .C(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__a21o_1 _25680_ (.A1(_01733_),
    .A2(_01734_),
    .B1(_01743_),
    .X(_01745_));
 sky130_fd_sc_hd__nand3_1 _25681_ (.A(_01725_),
    .B(_01744_),
    .C(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__a21o_1 _25682_ (.A1(net129),
    .A2(net119),
    .B1(_01739_),
    .X(_01747_));
 sky130_fd_sc_hd__nand2_1 _25683_ (.A(_01746_),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nand2_1 _25684_ (.A(_01748_),
    .B(_11614_),
    .Y(_01750_));
 sky130_fd_sc_hd__nand3_1 _25685_ (.A(_01746_),
    .B(_11616_),
    .C(_01747_),
    .Y(_01751_));
 sky130_fd_sc_hd__nand2_2 _25686_ (.A(_01750_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__or2_1 _25687_ (.A(_13197_),
    .B(_01730_),
    .X(_01753_));
 sky130_fd_sc_hd__nand2_1 _25688_ (.A(_01753_),
    .B(_01734_),
    .Y(_01754_));
 sky130_fd_sc_hd__nand2_1 _25689_ (.A(_01671_),
    .B(_01637_),
    .Y(_01755_));
 sky130_fd_sc_hd__xor2_1 _25690_ (.A(_01754_),
    .B(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__nand2_1 _25691_ (.A(_01725_),
    .B(_01756_),
    .Y(_01757_));
 sky130_fd_sc_hd__nand2_1 _25692_ (.A(_01590_),
    .B(_01730_),
    .Y(_01758_));
 sky130_fd_sc_hd__nand2_1 _25693_ (.A(_01757_),
    .B(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__or2_1 _25694_ (.A(_12771_),
    .B(_01759_),
    .X(_01761_));
 sky130_fd_sc_hd__nand2_1 _25695_ (.A(_01759_),
    .B(_12771_),
    .Y(_01762_));
 sky130_fd_sc_hd__nand2_1 _25696_ (.A(_01761_),
    .B(_01762_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _25697_ (.A(_01752_),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__nand2_2 _25698_ (.A(_01737_),
    .B(_01363_),
    .Y(_01765_));
 sky130_fd_sc_hd__xor2_1 _25699_ (.A(_01356_),
    .B(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__nand2_1 _25700_ (.A(_01766_),
    .B(_12002_),
    .Y(_01767_));
 sky130_fd_sc_hd__inv_2 _25701_ (.A(_01356_),
    .Y(_01768_));
 sky130_fd_sc_hd__or2_1 _25702_ (.A(_01768_),
    .B(_01765_),
    .X(_01769_));
 sky130_fd_sc_hd__nand2_1 _25703_ (.A(_01765_),
    .B(_01768_),
    .Y(_01770_));
 sky130_fd_sc_hd__nand3_2 _25704_ (.A(_01769_),
    .B(_12012_),
    .C(_01770_),
    .Y(_01772_));
 sky130_fd_sc_hd__nand3_1 _25705_ (.A(_01767_),
    .B(_01772_),
    .C(_01743_),
    .Y(_01773_));
 sky130_fd_sc_hd__inv_2 _25706_ (.A(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hd__nand3_2 _25707_ (.A(_01733_),
    .B(_01774_),
    .C(_01734_),
    .Y(_01775_));
 sky130_fd_sc_hd__inv_2 _25708_ (.A(_01741_),
    .Y(_01776_));
 sky130_fd_sc_hd__inv_2 _25709_ (.A(_01772_),
    .Y(_01777_));
 sky130_fd_sc_hd__a21oi_1 _25710_ (.A1(_01767_),
    .A2(_01776_),
    .B1(_01777_),
    .Y(_01778_));
 sky130_fd_sc_hd__nand2_1 _25711_ (.A(_01775_),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hd__nand2_1 _25712_ (.A(_01327_),
    .B(_01366_),
    .Y(_01780_));
 sky130_fd_sc_hd__inv_2 _25713_ (.A(_01370_),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _25714_ (.A(_01780_),
    .B(_01781_),
    .Y(_01783_));
 sky130_fd_sc_hd__clkinvlp_2 _25715_ (.A(_01339_),
    .Y(_01784_));
 sky130_fd_sc_hd__nand2_1 _25716_ (.A(_01783_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__nand3_1 _25717_ (.A(_01780_),
    .B(_01339_),
    .C(_01781_),
    .Y(_01786_));
 sky130_fd_sc_hd__nand2_1 _25718_ (.A(_01785_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__nand2_1 _25719_ (.A(_01787_),
    .B(_12017_),
    .Y(_01788_));
 sky130_fd_sc_hd__nand3_1 _25720_ (.A(_01785_),
    .B(_11986_),
    .C(_01786_),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_1 _25721_ (.A(_01788_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__or2b_1 _25722_ (.A(_01779_),
    .B_N(_01790_),
    .X(_01791_));
 sky130_fd_sc_hd__inv_2 _25723_ (.A(_01790_),
    .Y(_01792_));
 sky130_fd_sc_hd__nand2_1 _25724_ (.A(_01779_),
    .B(_01792_),
    .Y(_01794_));
 sky130_fd_sc_hd__nand3_1 _25725_ (.A(_01791_),
    .B(_01725_),
    .C(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__a21o_1 _25726_ (.A1(net129),
    .A2(net119),
    .B1(_01787_),
    .X(_01796_));
 sky130_fd_sc_hd__nand2_1 _25727_ (.A(_01795_),
    .B(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__nand2_1 _25728_ (.A(_01797_),
    .B(_11586_),
    .Y(_01798_));
 sky130_fd_sc_hd__nand3_1 _25729_ (.A(_01795_),
    .B(_11588_),
    .C(_01796_),
    .Y(_01799_));
 sky130_fd_sc_hd__nand2_2 _25730_ (.A(_01798_),
    .B(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2_1 _25731_ (.A(_01767_),
    .B(_01772_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_1 _25732_ (.A(_01744_),
    .B(_01741_),
    .Y(_01802_));
 sky130_fd_sc_hd__xor2_1 _25733_ (.A(_01801_),
    .B(_01802_),
    .X(_01803_));
 sky130_fd_sc_hd__nand2_1 _25734_ (.A(_01803_),
    .B(_01725_),
    .Y(_01805_));
 sky130_fd_sc_hd__nand2_2 _25735_ (.A(net233),
    .B(_01766_),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2_1 _25736_ (.A(_01805_),
    .B(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__nand2_1 _25737_ (.A(_01807_),
    .B(_11600_),
    .Y(_01808_));
 sky130_fd_sc_hd__nand3_4 _25738_ (.A(_01805_),
    .B(_11603_),
    .C(_01806_),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_2 _25739_ (.A(_01808_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_2 _25740_ (.A(_01800_),
    .B(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__nand2_1 _25741_ (.A(_01764_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__inv_2 _25742_ (.A(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__nand2_1 _25743_ (.A(_01724_),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__o21ai_1 _25744_ (.A1(_01761_),
    .A2(_01752_),
    .B1(_01750_),
    .Y(_01816_));
 sky130_fd_sc_hd__o21ai_1 _25745_ (.A1(_01809_),
    .A2(_01800_),
    .B1(_01798_),
    .Y(_01817_));
 sky130_fd_sc_hd__a21oi_1 _25746_ (.A1(_01816_),
    .A2(_01811_),
    .B1(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_2 _25747_ (.A(_01814_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__nand2_1 _25748_ (.A(_01785_),
    .B(_01338_),
    .Y(_01820_));
 sky130_fd_sc_hd__inv_2 _25749_ (.A(_01347_),
    .Y(_01821_));
 sky130_fd_sc_hd__nand2_1 _25750_ (.A(_01820_),
    .B(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__nand3_1 _25751_ (.A(_01785_),
    .B(_01347_),
    .C(_01338_),
    .Y(_01823_));
 sky130_fd_sc_hd__nand2_1 _25752_ (.A(_01822_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__nand2_1 _25753_ (.A(_01824_),
    .B(_11983_),
    .Y(_01825_));
 sky130_fd_sc_hd__nand3_2 _25754_ (.A(_01822_),
    .B(_11990_),
    .C(_01823_),
    .Y(_01827_));
 sky130_fd_sc_hd__nand3_1 _25755_ (.A(_01825_),
    .B(_01827_),
    .C(_01792_),
    .Y(_01828_));
 sky130_fd_sc_hd__inv_2 _25756_ (.A(_01789_),
    .Y(_01829_));
 sky130_fd_sc_hd__inv_2 _25757_ (.A(_01827_),
    .Y(_01830_));
 sky130_fd_sc_hd__a21o_1 _25758_ (.A1(_01825_),
    .A2(_01829_),
    .B1(_01830_),
    .X(_01831_));
 sky130_fd_sc_hd__nor2_1 _25759_ (.A(_01778_),
    .B(_01828_),
    .Y(_01832_));
 sky130_fd_sc_hd__nor2_1 _25760_ (.A(_01831_),
    .B(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__o21ai_2 _25761_ (.A1(_01828_),
    .A2(_01775_),
    .B1(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__inv_2 _25762_ (.A(_01379_),
    .Y(_01835_));
 sky130_fd_sc_hd__inv_2 _25763_ (.A(_01378_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _25764_ (.A(_01374_),
    .B(_01836_),
    .Y(_01838_));
 sky130_fd_sc_hd__nand2_1 _25765_ (.A(_01838_),
    .B(_01234_),
    .Y(_01839_));
 sky130_fd_sc_hd__or2_1 _25766_ (.A(_01835_),
    .B(_01839_),
    .X(_01840_));
 sky130_fd_sc_hd__nand2_1 _25767_ (.A(_01839_),
    .B(_01835_),
    .Y(_01841_));
 sky130_fd_sc_hd__nand2_1 _25768_ (.A(_01840_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__nand2_1 _25769_ (.A(_01842_),
    .B(_12118_),
    .Y(_01843_));
 sky130_fd_sc_hd__nand3_1 _25770_ (.A(_01840_),
    .B(_12120_),
    .C(_01841_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2_1 _25771_ (.A(_01843_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__inv_2 _25772_ (.A(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__or2_1 _25773_ (.A(_01836_),
    .B(_01374_),
    .X(_01847_));
 sky130_fd_sc_hd__nand2_1 _25774_ (.A(_01847_),
    .B(_01838_),
    .Y(_01849_));
 sky130_fd_sc_hd__inv_2 _25775_ (.A(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hd__nand2_1 _25776_ (.A(_01850_),
    .B(_11671_),
    .Y(_01851_));
 sky130_fd_sc_hd__nand2_1 _25777_ (.A(_01849_),
    .B(_12817_),
    .Y(_01852_));
 sky130_fd_sc_hd__nand2_1 _25778_ (.A(_01851_),
    .B(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__inv_4 _25779_ (.A(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__nand2_1 _25780_ (.A(_01846_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__inv_2 _25781_ (.A(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nand2_1 _25782_ (.A(_01834_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__inv_2 _25783_ (.A(_01851_),
    .Y(_01858_));
 sky130_fd_sc_hd__a21boi_2 _25784_ (.A1(_01843_),
    .A2(_01858_),
    .B1_N(_01844_),
    .Y(_01860_));
 sky130_fd_sc_hd__nand2_1 _25785_ (.A(_01857_),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__nand2_1 _25786_ (.A(_01374_),
    .B(_01380_),
    .Y(_01862_));
 sky130_fd_sc_hd__inv_2 _25787_ (.A(_01241_),
    .Y(_01863_));
 sky130_fd_sc_hd__nand2_1 _25788_ (.A(_01862_),
    .B(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__inv_2 _25789_ (.A(_01220_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _25790_ (.A(_01864_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand3_1 _25791_ (.A(_01862_),
    .B(_01863_),
    .C(_01220_),
    .Y(_01867_));
 sky130_fd_sc_hd__nand2_1 _25792_ (.A(_01866_),
    .B(_01867_),
    .Y(_01868_));
 sky130_fd_sc_hd__nand2_1 _25793_ (.A(_01868_),
    .B(_12149_),
    .Y(_01869_));
 sky130_fd_sc_hd__nand3_2 _25794_ (.A(_01866_),
    .B(_01867_),
    .C(_12147_),
    .Y(_01871_));
 sky130_fd_sc_hd__nand2_1 _25795_ (.A(_01869_),
    .B(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__inv_2 _25796_ (.A(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__nand2_1 _25797_ (.A(_01861_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__nand3_1 _25798_ (.A(_01857_),
    .B(_01872_),
    .C(_01860_),
    .Y(_01875_));
 sky130_fd_sc_hd__nand3_1 _25799_ (.A(_01874_),
    .B(_01725_),
    .C(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__or2_1 _25800_ (.A(_01868_),
    .B(_01725_),
    .X(_01877_));
 sky130_fd_sc_hd__nand2_1 _25801_ (.A(_01876_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__nand2_1 _25802_ (.A(_01878_),
    .B(_11701_),
    .Y(_01879_));
 sky130_fd_sc_hd__nand3_1 _25803_ (.A(_01876_),
    .B(_11703_),
    .C(_01877_),
    .Y(_01880_));
 sky130_fd_sc_hd__nand2_1 _25804_ (.A(_01879_),
    .B(_01880_),
    .Y(_01882_));
 sky130_fd_sc_hd__nand2_1 _25805_ (.A(_01834_),
    .B(_01854_),
    .Y(_01883_));
 sky130_fd_sc_hd__nand2_1 _25806_ (.A(_01883_),
    .B(_01851_),
    .Y(_01884_));
 sky130_fd_sc_hd__nand2_1 _25807_ (.A(_01884_),
    .B(_01846_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand3_1 _25808_ (.A(_01883_),
    .B(_01845_),
    .C(_01851_),
    .Y(_01886_));
 sky130_fd_sc_hd__nand2_1 _25809_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__nand2_1 _25810_ (.A(_01887_),
    .B(_01725_),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_1 _25811_ (.A(net233),
    .B(_01842_),
    .Y(_01889_));
 sky130_fd_sc_hd__nand2_1 _25812_ (.A(_01888_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hd__nand2_1 _25813_ (.A(_01890_),
    .B(_11715_),
    .Y(_01891_));
 sky130_fd_sc_hd__nand3_1 _25814_ (.A(_01888_),
    .B(_11717_),
    .C(_01889_),
    .Y(_01893_));
 sky130_fd_sc_hd__nand2_1 _25815_ (.A(_01891_),
    .B(_01893_),
    .Y(_01894_));
 sky130_fd_sc_hd__nor2_2 _25816_ (.A(_01882_),
    .B(_01894_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _25817_ (.A(_01854_),
    .B(_01834_),
    .Y(_01896_));
 sky130_fd_sc_hd__nand2_1 _25818_ (.A(_01883_),
    .B(_01725_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_1 _25819_ (.A(net233),
    .B(_01850_),
    .Y(_01898_));
 sky130_fd_sc_hd__o211ai_1 _25820_ (.A1(_01896_),
    .A2(_01897_),
    .B1(_13304_),
    .C1(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__o21ai_1 _25821_ (.A1(_01896_),
    .A2(_01897_),
    .B1(_01898_),
    .Y(_01900_));
 sky130_fd_sc_hd__nand2_1 _25822_ (.A(_01900_),
    .B(_06149_),
    .Y(_01901_));
 sky130_fd_sc_hd__nand2_1 _25823_ (.A(_01899_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__nand2_1 _25824_ (.A(_01825_),
    .B(_01827_),
    .Y(_01904_));
 sky130_fd_sc_hd__nand2_1 _25825_ (.A(_01794_),
    .B(_01789_),
    .Y(_01905_));
 sky130_fd_sc_hd__xor2_1 _25826_ (.A(_01904_),
    .B(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__buf_6 _25827_ (.A(_01725_),
    .X(_01907_));
 sky130_fd_sc_hd__nand2_1 _25828_ (.A(_01906_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__nand2_1 _25829_ (.A(\div1i.quot[1] ),
    .B(_01824_),
    .Y(_01909_));
 sky130_fd_sc_hd__nand2_1 _25830_ (.A(_01908_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__nand2_1 _25831_ (.A(_01910_),
    .B(_11185_),
    .Y(_01911_));
 sky130_fd_sc_hd__nand3_1 _25832_ (.A(_01908_),
    .B(_12187_),
    .C(_01909_),
    .Y(_01912_));
 sky130_fd_sc_hd__nand2_2 _25833_ (.A(_01911_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_2 _25834_ (.A(_01902_),
    .B(_01913_),
    .Y(_01915_));
 sky130_fd_sc_hd__nand2_1 _25835_ (.A(_01895_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__inv_2 _25836_ (.A(_01916_),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_2 _25837_ (.A(_01819_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__o21ai_1 _25838_ (.A1(_01912_),
    .A2(_01902_),
    .B1(_01901_),
    .Y(_01919_));
 sky130_fd_sc_hd__o21ai_1 _25839_ (.A1(_01893_),
    .A2(_01882_),
    .B1(_01879_),
    .Y(_01920_));
 sky130_fd_sc_hd__a21oi_2 _25840_ (.A1(_01895_),
    .A2(_01919_),
    .B1(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__nand2_4 _25841_ (.A(_01918_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__nand2_1 _25842_ (.A(_01866_),
    .B(_01219_),
    .Y(_01923_));
 sky130_fd_sc_hd__inv_2 _25843_ (.A(_01208_),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_1 _25844_ (.A(_01923_),
    .B(_01924_),
    .Y(_01926_));
 sky130_fd_sc_hd__nand3_1 _25845_ (.A(_01866_),
    .B(_01208_),
    .C(_01219_),
    .Y(_01927_));
 sky130_fd_sc_hd__nand2_1 _25846_ (.A(_01926_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_1 _25847_ (.A(_01928_),
    .B(_12894_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand3_1 _25848_ (.A(_01926_),
    .B(_11754_),
    .C(_01927_),
    .Y(_01930_));
 sky130_fd_sc_hd__nand3_1 _25849_ (.A(_01929_),
    .B(_01930_),
    .C(_01873_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _25850_ (.A(_01931_),
    .B(_01855_),
    .Y(_01932_));
 sky130_fd_sc_hd__nand2_2 _25851_ (.A(_01834_),
    .B(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__nor2_1 _25852_ (.A(_01931_),
    .B(_01860_),
    .Y(_01934_));
 sky130_fd_sc_hd__nand2_1 _25853_ (.A(_01929_),
    .B(_01930_),
    .Y(_01935_));
 sky130_fd_sc_hd__o21ai_1 _25854_ (.A1(_01871_),
    .A2(_01935_),
    .B1(_01930_),
    .Y(_01937_));
 sky130_fd_sc_hd__nor2_1 _25855_ (.A(_01934_),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__nand2_1 _25856_ (.A(_01933_),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__clkinvlp_2 _25857_ (.A(_01417_),
    .Y(_01940_));
 sky130_fd_sc_hd__inv_2 _25858_ (.A(_01427_),
    .Y(_01941_));
 sky130_fd_sc_hd__nand2_1 _25859_ (.A(_01382_),
    .B(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__nand2_1 _25860_ (.A(_01942_),
    .B(_01426_),
    .Y(_01943_));
 sky130_fd_sc_hd__or2_1 _25861_ (.A(_01940_),
    .B(_01943_),
    .X(_01944_));
 sky130_fd_sc_hd__nand2_1 _25862_ (.A(_01943_),
    .B(_01940_),
    .Y(_01945_));
 sky130_fd_sc_hd__nand2_1 _25863_ (.A(_01944_),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__nand2_1 _25864_ (.A(_01946_),
    .B(_12914_),
    .Y(_01948_));
 sky130_fd_sc_hd__nand3_1 _25865_ (.A(_01944_),
    .B(_11774_),
    .C(_01945_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_1 _25866_ (.A(_01948_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__inv_2 _25867_ (.A(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__or2_1 _25868_ (.A(_01941_),
    .B(_01382_),
    .X(_01952_));
 sky130_fd_sc_hd__nand2_1 _25869_ (.A(_01952_),
    .B(_01942_),
    .Y(_01953_));
 sky130_fd_sc_hd__inv_2 _25870_ (.A(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__nand2_2 _25871_ (.A(_01954_),
    .B(_11199_),
    .Y(_01955_));
 sky130_fd_sc_hd__nand2_1 _25872_ (.A(_01953_),
    .B(_13461_),
    .Y(_01956_));
 sky130_fd_sc_hd__nand2_1 _25873_ (.A(_01955_),
    .B(_01956_),
    .Y(_01957_));
 sky130_fd_sc_hd__inv_2 _25874_ (.A(_01957_),
    .Y(_01959_));
 sky130_fd_sc_hd__nand2_1 _25875_ (.A(_01951_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__inv_2 _25876_ (.A(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_1 _25877_ (.A(_01939_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__inv_2 _25878_ (.A(_01955_),
    .Y(_01963_));
 sky130_fd_sc_hd__a21boi_2 _25879_ (.A1(_01948_),
    .A2(_01963_),
    .B1_N(_01949_),
    .Y(_01964_));
 sky130_fd_sc_hd__nand2_1 _25880_ (.A(_01962_),
    .B(_01964_),
    .Y(_01965_));
 sky130_fd_sc_hd__inv_2 _25881_ (.A(_01472_),
    .Y(_01966_));
 sky130_fd_sc_hd__nand2_1 _25882_ (.A(_01433_),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__nand3_1 _25883_ (.A(_01429_),
    .B(_01432_),
    .C(_01472_),
    .Y(_01968_));
 sky130_fd_sc_hd__nand2_1 _25884_ (.A(_01967_),
    .B(_01968_),
    .Y(_01970_));
 sky130_fd_sc_hd__inv_2 _25885_ (.A(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__nand2_1 _25886_ (.A(_01971_),
    .B(_11797_),
    .Y(_01972_));
 sky130_fd_sc_hd__nand2_1 _25887_ (.A(_01970_),
    .B(_12939_),
    .Y(_01973_));
 sky130_fd_sc_hd__nand2_1 _25888_ (.A(_01972_),
    .B(_01973_),
    .Y(_01974_));
 sky130_fd_sc_hd__inv_2 _25889_ (.A(_01974_),
    .Y(_01975_));
 sky130_fd_sc_hd__nand2_1 _25890_ (.A(_01965_),
    .B(_01975_),
    .Y(_01976_));
 sky130_fd_sc_hd__nand3_1 _25891_ (.A(_01962_),
    .B(_01974_),
    .C(_01964_),
    .Y(_01977_));
 sky130_fd_sc_hd__nand3_1 _25892_ (.A(_01976_),
    .B(_01907_),
    .C(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__nand2_1 _25893_ (.A(\div1i.quot[1] ),
    .B(_01971_),
    .Y(_01979_));
 sky130_fd_sc_hd__nand2_1 _25894_ (.A(_01978_),
    .B(_01979_),
    .Y(_01981_));
 sky130_fd_sc_hd__nand2_1 _25895_ (.A(_01981_),
    .B(_11808_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand3_1 _25896_ (.A(_01978_),
    .B(_11811_),
    .C(_01979_),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _25897_ (.A(_01982_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__nand2_1 _25898_ (.A(_01939_),
    .B(_01959_),
    .Y(_01985_));
 sky130_fd_sc_hd__nand2_1 _25899_ (.A(_01985_),
    .B(_01955_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_1 _25900_ (.A(_01986_),
    .B(_01951_),
    .Y(_01987_));
 sky130_fd_sc_hd__nand3_1 _25901_ (.A(_01985_),
    .B(_01950_),
    .C(_01955_),
    .Y(_01988_));
 sky130_fd_sc_hd__a21o_1 _25902_ (.A1(_01987_),
    .A2(_01988_),
    .B1(\div1i.quot[1] ),
    .X(_01989_));
 sky130_fd_sc_hd__nand2_1 _25903_ (.A(\div1i.quot[1] ),
    .B(_01946_),
    .Y(_01990_));
 sky130_fd_sc_hd__nand2_1 _25904_ (.A(_01989_),
    .B(_01990_),
    .Y(_01992_));
 sky130_fd_sc_hd__nand2_1 _25905_ (.A(_01992_),
    .B(_13537_),
    .Y(_01993_));
 sky130_fd_sc_hd__nand3_1 _25906_ (.A(_01989_),
    .B(_07400_),
    .C(_01990_),
    .Y(_01994_));
 sky130_fd_sc_hd__nand2_1 _25907_ (.A(_01993_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_2 _25908_ (.A(_01984_),
    .B(_01995_),
    .Y(_01996_));
 sky130_fd_sc_hd__nand3_1 _25909_ (.A(_01933_),
    .B(_01938_),
    .C(_01957_),
    .Y(_01997_));
 sky130_fd_sc_hd__nand3_1 _25910_ (.A(_01985_),
    .B(_01725_),
    .C(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__nand2_1 _25911_ (.A(net233),
    .B(_01954_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand2_1 _25912_ (.A(_01998_),
    .B(_01999_),
    .Y(_02000_));
 sky130_fd_sc_hd__or2_1 _25913_ (.A(_13502_),
    .B(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__nand2_1 _25914_ (.A(_02000_),
    .B(_13502_),
    .Y(_02003_));
 sky130_fd_sc_hd__nand2_1 _25915_ (.A(_02001_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__a21o_1 _25916_ (.A1(_01874_),
    .A2(_01871_),
    .B1(_01935_),
    .X(_02005_));
 sky130_fd_sc_hd__nand3_1 _25917_ (.A(_01874_),
    .B(_01935_),
    .C(_01871_),
    .Y(_02006_));
 sky130_fd_sc_hd__nand2_1 _25918_ (.A(_02005_),
    .B(_02006_),
    .Y(_02007_));
 sky130_fd_sc_hd__nand2_1 _25919_ (.A(_02007_),
    .B(_01907_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2_1 _25920_ (.A(\div1i.quot[1] ),
    .B(_01928_),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _25921_ (.A(_02008_),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__nand2_1 _25922_ (.A(_02010_),
    .B(_11838_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand3_2 _25923_ (.A(_02008_),
    .B(_11840_),
    .C(_02009_),
    .Y(_02012_));
 sky130_fd_sc_hd__nand3b_1 _25924_ (.A_N(_02004_),
    .B(_02011_),
    .C(_02012_),
    .Y(_02014_));
 sky130_fd_sc_hd__inv_2 _25925_ (.A(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__nand3_4 _25926_ (.A(_01922_),
    .B(_01996_),
    .C(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__o21ai_1 _25927_ (.A1(_02004_),
    .A2(_02012_),
    .B1(_02003_),
    .Y(_02017_));
 sky130_fd_sc_hd__o21ai_1 _25928_ (.A1(_01994_),
    .A2(_01984_),
    .B1(_01982_),
    .Y(_02018_));
 sky130_fd_sc_hd__a21oi_2 _25929_ (.A1(_01996_),
    .A2(_02017_),
    .B1(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__nand2_4 _25930_ (.A(_02016_),
    .B(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__nand2_1 _25931_ (.A(_01967_),
    .B(_01470_),
    .Y(_02021_));
 sky130_fd_sc_hd__inv_2 _25932_ (.A(_01463_),
    .Y(_02022_));
 sky130_fd_sc_hd__nand2_1 _25933_ (.A(_02021_),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__nand3_1 _25934_ (.A(_01967_),
    .B(_01463_),
    .C(_01470_),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_1 _25935_ (.A(_02023_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__nand2_1 _25936_ (.A(_02026_),
    .B(_12992_),
    .Y(_02027_));
 sky130_fd_sc_hd__nand3_1 _25937_ (.A(_02023_),
    .B(_11858_),
    .C(_02025_),
    .Y(_02028_));
 sky130_fd_sc_hd__nand3_1 _25938_ (.A(_01975_),
    .B(_02027_),
    .C(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__inv_2 _25939_ (.A(_02029_),
    .Y(_02030_));
 sky130_fd_sc_hd__nand3_1 _25940_ (.A(_01939_),
    .B(_01961_),
    .C(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__inv_2 _25941_ (.A(_02027_),
    .Y(_02032_));
 sky130_fd_sc_hd__o21ai_1 _25942_ (.A1(_01972_),
    .A2(_02032_),
    .B1(_02028_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_1 _25943_ (.A(_01964_),
    .B(_02029_),
    .Y(_02034_));
 sky130_fd_sc_hd__nor2_1 _25944_ (.A(_02033_),
    .B(_02034_),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2_1 _25945_ (.A(_02031_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__inv_2 _25946_ (.A(_01478_),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2_1 _25947_ (.A(_01523_),
    .B(_01524_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2_1 _25948_ (.A(_02038_),
    .B(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__inv_2 _25949_ (.A(_02039_),
    .Y(_02041_));
 sky130_fd_sc_hd__nand2_1 _25950_ (.A(_01478_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_1 _25951_ (.A(_02040_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__nand2_1 _25952_ (.A(_02043_),
    .B(_14113_),
    .Y(_02044_));
 sky130_fd_sc_hd__nand3_2 _25953_ (.A(_02040_),
    .B(_08554_),
    .C(_02042_),
    .Y(_02045_));
 sky130_fd_sc_hd__nand2_1 _25954_ (.A(_02044_),
    .B(_02045_),
    .Y(_02047_));
 sky130_fd_sc_hd__inv_2 _25955_ (.A(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__nand2_1 _25956_ (.A(_02037_),
    .B(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__nand3_1 _25957_ (.A(_02031_),
    .B(_02036_),
    .C(_02047_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand3_1 _25958_ (.A(_02049_),
    .B(_02050_),
    .C(_01907_),
    .Y(_02051_));
 sky130_fd_sc_hd__or2_1 _25959_ (.A(_02043_),
    .B(_01907_),
    .X(_02052_));
 sky130_fd_sc_hd__nand2_1 _25960_ (.A(_02051_),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_1 _25961_ (.A(_02053_),
    .B(_13022_),
    .Y(_02054_));
 sky130_fd_sc_hd__nand3_1 _25962_ (.A(_02051_),
    .B(_08020_),
    .C(_02052_),
    .Y(_02055_));
 sky130_fd_sc_hd__nand2_1 _25963_ (.A(_02054_),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hd__nand2_1 _25964_ (.A(_02027_),
    .B(_02028_),
    .Y(_02058_));
 sky130_fd_sc_hd__a21o_1 _25965_ (.A1(_01976_),
    .A2(_01972_),
    .B1(_02058_),
    .X(_02059_));
 sky130_fd_sc_hd__nand3_1 _25966_ (.A(_01976_),
    .B(_01972_),
    .C(_02058_),
    .Y(_02060_));
 sky130_fd_sc_hd__nand2_1 _25967_ (.A(_02059_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _25968_ (.A(_02061_),
    .B(_01907_),
    .Y(_02062_));
 sky130_fd_sc_hd__nand2_1 _25969_ (.A(\div1i.quot[1] ),
    .B(_02026_),
    .Y(_02063_));
 sky130_fd_sc_hd__nand2_1 _25970_ (.A(_02062_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__nand2_1 _25971_ (.A(_02064_),
    .B(_11896_),
    .Y(_02065_));
 sky130_fd_sc_hd__nand3_2 _25972_ (.A(_02062_),
    .B(_11899_),
    .C(_02063_),
    .Y(_02066_));
 sky130_fd_sc_hd__nand3b_1 _25973_ (.A_N(_02056_),
    .B(_02065_),
    .C(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__nand2_1 _25974_ (.A(_02049_),
    .B(_02045_),
    .Y(_02069_));
 sky130_fd_sc_hd__nand2_1 _25975_ (.A(_02042_),
    .B(_01524_),
    .Y(_02070_));
 sky130_fd_sc_hd__or2_1 _25976_ (.A(_01515_),
    .B(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__nand2_1 _25977_ (.A(_02070_),
    .B(_01515_),
    .Y(_02072_));
 sky130_fd_sc_hd__nand2_1 _25978_ (.A(_02071_),
    .B(_02072_),
    .Y(_02073_));
 sky130_fd_sc_hd__nand2_1 _25979_ (.A(_02073_),
    .B(_13042_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand3_1 _25980_ (.A(_02071_),
    .B(_12495_),
    .C(_02072_),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_1 _25981_ (.A(_02074_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__inv_2 _25982_ (.A(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_1 _25983_ (.A(_02069_),
    .B(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__nand3_1 _25984_ (.A(_02049_),
    .B(_02076_),
    .C(_02045_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _25985_ (.A(_02078_),
    .B(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hd__nand2_1 _25986_ (.A(_02081_),
    .B(_01907_),
    .Y(_02082_));
 sky130_fd_sc_hd__nand2_1 _25987_ (.A(_02073_),
    .B(\div1i.quot[1] ),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _25988_ (.A(_02082_),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__nand2_1 _25989_ (.A(_02084_),
    .B(_12506_),
    .Y(_02085_));
 sky130_fd_sc_hd__nand3_1 _25990_ (.A(_02082_),
    .B(_11376_),
    .C(_02083_),
    .Y(_02086_));
 sky130_fd_sc_hd__nand2_1 _25991_ (.A(_02085_),
    .B(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__inv_2 _25992_ (.A(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__nand3_1 _25993_ (.A(_02074_),
    .B(_02075_),
    .C(_02048_),
    .Y(_02089_));
 sky130_fd_sc_hd__inv_2 _25994_ (.A(_02089_),
    .Y(_02091_));
 sky130_fd_sc_hd__nand2_1 _25995_ (.A(_02037_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__clkinvlp_2 _25996_ (.A(_02045_),
    .Y(_02093_));
 sky130_fd_sc_hd__a21boi_1 _25997_ (.A1(_02074_),
    .A2(_02093_),
    .B1_N(_02075_),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_1 _25998_ (.A(_02092_),
    .B(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__o21bai_1 _25999_ (.A1(_01525_),
    .A2(_02038_),
    .B1_N(_01576_),
    .Y(_02096_));
 sky130_fd_sc_hd__or2_1 _26000_ (.A(_01546_),
    .B(_02096_),
    .X(_02097_));
 sky130_fd_sc_hd__nand2_1 _26001_ (.A(_02096_),
    .B(_01546_),
    .Y(_02098_));
 sky130_fd_sc_hd__nand2_1 _26002_ (.A(_02097_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hd__inv_2 _26003_ (.A(_02099_),
    .Y(_02100_));
 sky130_fd_sc_hd__nand2_1 _26004_ (.A(_02100_),
    .B(_11935_),
    .Y(_02102_));
 sky130_fd_sc_hd__nand2_1 _26005_ (.A(_02099_),
    .B(_13633_),
    .Y(_02103_));
 sky130_fd_sc_hd__nand2_1 _26006_ (.A(_02102_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__inv_2 _26007_ (.A(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__nand2_1 _26008_ (.A(_02095_),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__nand3_1 _26009_ (.A(_02092_),
    .B(_02094_),
    .C(_02104_),
    .Y(_02107_));
 sky130_fd_sc_hd__nand3_1 _26010_ (.A(_02106_),
    .B(_01907_),
    .C(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__nand2_1 _26011_ (.A(_02100_),
    .B(\div1i.quot[1] ),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _26012_ (.A(_02108_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__nand2_1 _26013_ (.A(_02110_),
    .B(_11946_),
    .Y(_02111_));
 sky130_fd_sc_hd__nand3_1 _26014_ (.A(_02108_),
    .B(_11948_),
    .C(_02109_),
    .Y(_02113_));
 sky130_fd_sc_hd__nand2_2 _26015_ (.A(_02111_),
    .B(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__inv_2 _26016_ (.A(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2_1 _26017_ (.A(_02088_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__nor2_1 _26018_ (.A(_02067_),
    .B(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__nand2_2 _26019_ (.A(_02020_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_1 _26020_ (.A(_02114_),
    .B(_02087_),
    .Y(_02119_));
 sky130_fd_sc_hd__o21ai_1 _26021_ (.A1(_02056_),
    .A2(_02066_),
    .B1(_02054_),
    .Y(_02120_));
 sky130_fd_sc_hd__o21ai_1 _26022_ (.A1(_02086_),
    .A2(_02114_),
    .B1(_02111_),
    .Y(_02121_));
 sky130_fd_sc_hd__a21oi_2 _26023_ (.A1(_02119_),
    .A2(_02120_),
    .B1(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__nand2_2 _26024_ (.A(_02118_),
    .B(_02122_),
    .Y(_02123_));
 sky130_fd_sc_hd__nand2_1 _26025_ (.A(_02098_),
    .B(_01544_),
    .Y(_02124_));
 sky130_fd_sc_hd__xor2_2 _26026_ (.A(_01570_),
    .B(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__nand3_1 _26027_ (.A(_02106_),
    .B(_01907_),
    .C(_02102_),
    .Y(_02126_));
 sky130_fd_sc_hd__xnor2_2 _26028_ (.A(_02125_),
    .B(_02126_),
    .Y(_02127_));
 sky130_fd_sc_hd__nand2_4 _26029_ (.A(_02123_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__clkinvlp_2 _26030_ (.A(_02127_),
    .Y(_02129_));
 sky130_fd_sc_hd__nand3_4 _26031_ (.A(_02118_),
    .B(_02122_),
    .C(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__nand2_8 _26032_ (.A(_02128_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__buf_8 _26033_ (.A(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__buf_6 _26034_ (.A(_02132_),
    .X(\div1i.quot[0] ));
 sky130_fd_sc_hd__buf_6 _26035_ (.A(net160),
    .X(_02134_));
 sky130_fd_sc_hd__xnor2_4 _26036_ (.A(net57),
    .B(net25),
    .Y(_02135_));
 sky130_fd_sc_hd__nand2_1 _26037_ (.A(net150),
    .B(_02134_),
    .Y(_02136_));
 sky130_fd_sc_hd__o21ai_1 _26038_ (.A1(_02134_),
    .A2(net107),
    .B1(net151),
    .Y(_00027_));
 sky130_fd_sc_hd__nor2_2 _26039_ (.A(net185),
    .B(net200),
    .Y(_02137_));
 sky130_fd_sc_hd__inv_2 _26040_ (.A(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__mux2_1 _26041_ (.A0(\M00r[20] ),
    .A1(\M00r[21] ),
    .S(net185),
    .X(_02139_));
 sky130_fd_sc_hd__inv_2 _26042_ (.A(net177),
    .Y(_02140_));
 sky130_fd_sc_hd__nand2_1 _26043_ (.A(net178),
    .B(net185),
    .Y(_02141_));
 sky130_fd_sc_hd__o21ai_1 _26044_ (.A1(net185),
    .A2(net214),
    .B1(_02141_),
    .Y(_02143_));
 sky130_fd_sc_hd__nand2_1 _26045_ (.A(_02143_),
    .B(_02138_),
    .Y(_02144_));
 sky130_fd_sc_hd__o21ai_1 _26046_ (.A1(_02138_),
    .A2(_02139_),
    .B1(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__inv_2 _26047_ (.A(net185),
    .Y(_02146_));
 sky130_fd_sc_hd__nand2_1 _26048_ (.A(_02146_),
    .B(net178),
    .Y(_02147_));
 sky130_fd_sc_hd__o21ai_1 _26049_ (.A1(net200),
    .A2(_02146_),
    .B1(net179),
    .Y(_02148_));
 sky130_fd_sc_hd__mux2_1 _26050_ (.A0(net180),
    .A1(_02143_),
    .S(_02137_),
    .X(_02149_));
 sky130_fd_sc_hd__nand2_1 _26051_ (.A(net180),
    .B(_02137_),
    .Y(_02150_));
 sky130_fd_sc_hd__mux2_1 _26052_ (.A0(_02145_),
    .A1(_02149_),
    .S(net181),
    .X(_02151_));
 sky130_fd_sc_hd__inv_2 _26053_ (.A(net181),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_4 _26054_ (.A(_02149_),
    .B(_02152_),
    .Y(_02154_));
 sky130_fd_sc_hd__clkinv_4 _26055_ (.A(_02154_),
    .Y(_02155_));
 sky130_fd_sc_hd__nand2_1 _26056_ (.A(net182),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__clkbuf_4 _26057_ (.A(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__mux2_1 _26058_ (.A0(\M00r[18] ),
    .A1(net201),
    .S(net185),
    .X(_02158_));
 sky130_fd_sc_hd__mux2_1 _26059_ (.A0(\M00r[17] ),
    .A1(\M00r[18] ),
    .S(\M00r[24] ),
    .X(_02159_));
 sky130_fd_sc_hd__mux2_1 _26060_ (.A0(_02158_),
    .A1(_02159_),
    .S(_02137_),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_1 _26061_ (.A0(net201),
    .A1(\M00r[20] ),
    .S(net185),
    .X(_02161_));
 sky130_fd_sc_hd__buf_6 _26062_ (.A(_02138_),
    .X(_02162_));
 sky130_fd_sc_hd__mux2_1 _26063_ (.A0(_02158_),
    .A1(net202),
    .S(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__clkbuf_4 _26064_ (.A(net181),
    .X(_02165_));
 sky130_fd_sc_hd__mux2_1 _26065_ (.A0(_02160_),
    .A1(_02163_),
    .S(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__mux2_1 _26066_ (.A0(_02139_),
    .A1(net202),
    .S(_02137_),
    .X(_02167_));
 sky130_fd_sc_hd__mux2_1 _26067_ (.A0(_02163_),
    .A1(net203),
    .S(net181),
    .X(_02168_));
 sky130_fd_sc_hd__mux2_1 _26068_ (.A0(_02166_),
    .A1(_02168_),
    .S(_02154_),
    .X(_02169_));
 sky130_fd_sc_hd__inv_2 _26069_ (.A(net183),
    .Y(_02170_));
 sky130_fd_sc_hd__nand2_1 _26070_ (.A(_02145_),
    .B(_02165_),
    .Y(_02171_));
 sky130_fd_sc_hd__o21ai_1 _26071_ (.A1(_02165_),
    .A2(net203),
    .B1(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_1 _26072_ (.A(_02168_),
    .B(_02155_),
    .Y(_02173_));
 sky130_fd_sc_hd__o21ai_1 _26073_ (.A1(_02155_),
    .A2(net204),
    .B1(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__or2_1 _26074_ (.A(_02170_),
    .B(_02174_),
    .X(_02176_));
 sky130_fd_sc_hd__o21ai_1 _26075_ (.A1(_02157_),
    .A2(_02169_),
    .B1(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__mux2_1 _26076_ (.A0(net204),
    .A1(net182),
    .S(_02154_),
    .X(_02178_));
 sky130_fd_sc_hd__nand2_1 _26077_ (.A(_02178_),
    .B(_02157_),
    .Y(_02179_));
 sky130_fd_sc_hd__o21ai_2 _26078_ (.A1(_02157_),
    .A2(net205),
    .B1(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_1 _26079_ (.A(_02178_),
    .B(_02170_),
    .Y(_02181_));
 sky130_fd_sc_hd__clkbuf_4 _26080_ (.A(_02181_),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_1 _26081_ (.A0(_02177_),
    .A1(_02180_),
    .S(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__clkbuf_4 _26082_ (.A(net185),
    .X(_02184_));
 sky130_fd_sc_hd__mux2_1 _26083_ (.A0(\M00r[16] ),
    .A1(\M00r[17] ),
    .S(_02184_),
    .X(_02185_));
 sky130_fd_sc_hd__mux2_1 _26084_ (.A0(_02185_),
    .A1(_02159_),
    .S(_02162_),
    .X(_02187_));
 sky130_fd_sc_hd__mux2_1 _26085_ (.A0(_02187_),
    .A1(_02160_),
    .S(_02165_),
    .X(_02188_));
 sky130_fd_sc_hd__mux2_1 _26086_ (.A0(_02188_),
    .A1(_02166_),
    .S(_02154_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _26087_ (.A0(_02189_),
    .A1(_02169_),
    .S(_02157_),
    .X(_02190_));
 sky130_fd_sc_hd__nand2_1 _26088_ (.A(_02177_),
    .B(_02182_),
    .Y(_02191_));
 sky130_fd_sc_hd__o21ai_1 _26089_ (.A1(_02182_),
    .A2(_02190_),
    .B1(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hd__inv_2 _26090_ (.A(_02181_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand2_4 _26091_ (.A(_02180_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__inv_2 _26092_ (.A(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hd__mux2_1 _26093_ (.A0(_02183_),
    .A1(_02192_),
    .S(_02195_),
    .X(_02196_));
 sky130_fd_sc_hd__nand2_4 _26094_ (.A(_02183_),
    .B(_02195_),
    .Y(_02198_));
 sky130_fd_sc_hd__inv_2 _26095_ (.A(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__nand2_4 _26096_ (.A(_02196_),
    .B(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__mux2_1 _26097_ (.A0(\M00r[14] ),
    .A1(\M00r[15] ),
    .S(_02184_),
    .X(_02201_));
 sky130_fd_sc_hd__mux2_1 _26098_ (.A0(\M00r[13] ),
    .A1(\M00r[14] ),
    .S(_02184_),
    .X(_02202_));
 sky130_fd_sc_hd__buf_6 _26099_ (.A(_02137_),
    .X(_02203_));
 sky130_fd_sc_hd__mux2_1 _26100_ (.A0(_02201_),
    .A1(_02202_),
    .S(_02203_),
    .X(_02204_));
 sky130_fd_sc_hd__mux2_1 _26101_ (.A0(\M00r[15] ),
    .A1(\M00r[16] ),
    .S(_02184_),
    .X(_02205_));
 sky130_fd_sc_hd__mux2_1 _26102_ (.A0(_02201_),
    .A1(_02205_),
    .S(_02162_),
    .X(_02206_));
 sky130_fd_sc_hd__mux2_1 _26103_ (.A0(_02204_),
    .A1(_02206_),
    .S(_02165_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _26104_ (.A0(_02185_),
    .A1(_02205_),
    .S(_02203_),
    .X(_02209_));
 sky130_fd_sc_hd__mux2_1 _26105_ (.A0(_02206_),
    .A1(_02209_),
    .S(_02165_),
    .X(_02210_));
 sky130_fd_sc_hd__mux2_1 _26106_ (.A0(_02207_),
    .A1(_02210_),
    .S(_02154_),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _26107_ (.A0(_02209_),
    .A1(_02187_),
    .S(_02165_),
    .X(_02212_));
 sky130_fd_sc_hd__mux2_1 _26108_ (.A0(_02210_),
    .A1(_02212_),
    .S(_02154_),
    .X(_02213_));
 sky130_fd_sc_hd__mux2_1 _26109_ (.A0(_02211_),
    .A1(_02213_),
    .S(_02157_),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _26110_ (.A0(_02212_),
    .A1(_02188_),
    .S(_02154_),
    .X(_02215_));
 sky130_fd_sc_hd__mux2_1 _26111_ (.A0(_02213_),
    .A1(_02215_),
    .S(_02157_),
    .X(_02216_));
 sky130_fd_sc_hd__mux2_1 _26112_ (.A0(_02214_),
    .A1(_02216_),
    .S(_02182_),
    .X(_02217_));
 sky130_fd_sc_hd__mux2_1 _26113_ (.A0(_02215_),
    .A1(_02189_),
    .S(_02157_),
    .X(_02218_));
 sky130_fd_sc_hd__mux2_1 _26114_ (.A0(_02216_),
    .A1(_02218_),
    .S(_02182_),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _26115_ (.A0(_02217_),
    .A1(_02220_),
    .S(_02194_),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _26116_ (.A0(_02218_),
    .A1(_02190_),
    .S(_02182_),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _26117_ (.A0(_02220_),
    .A1(_02222_),
    .S(_02194_),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _26118_ (.A0(_02221_),
    .A1(_02223_),
    .S(_02198_),
    .X(_02224_));
 sky130_fd_sc_hd__nand2_1 _26119_ (.A(_02192_),
    .B(_02194_),
    .Y(_02225_));
 sky130_fd_sc_hd__o21ai_1 _26120_ (.A1(_02194_),
    .A2(_02222_),
    .B1(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2_1 _26121_ (.A(_02226_),
    .B(_02198_),
    .Y(_02227_));
 sky130_fd_sc_hd__o21ai_1 _26122_ (.A1(_02198_),
    .A2(_02223_),
    .B1(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__nand2_1 _26123_ (.A(_02228_),
    .B(_02200_),
    .Y(_02229_));
 sky130_fd_sc_hd__o21ai_1 _26124_ (.A1(_02200_),
    .A2(_02224_),
    .B1(_02229_),
    .Y(_02231_));
 sky130_fd_sc_hd__mux2_1 _26125_ (.A0(_02196_),
    .A1(_02226_),
    .S(_02199_),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _26126_ (.A0(_02228_),
    .A1(_02232_),
    .S(_02200_),
    .X(_02233_));
 sky130_fd_sc_hd__clkinv_4 _26127_ (.A(_02200_),
    .Y(_02234_));
 sky130_fd_sc_hd__nand2_4 _26128_ (.A(_02232_),
    .B(_02234_),
    .Y(_02235_));
 sky130_fd_sc_hd__mux2_1 _26129_ (.A0(_02231_),
    .A1(_02233_),
    .S(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__clkinv_4 _26130_ (.A(_02235_),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_2 _26131_ (.A(_02233_),
    .B(_02237_),
    .Y(_02238_));
 sky130_fd_sc_hd__inv_2 _26132_ (.A(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__nand2_4 _26133_ (.A(_02236_),
    .B(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__clkbuf_4 _26134_ (.A(_02240_),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_1 _26135_ (.A0(\M00r[10] ),
    .A1(\M00r[11] ),
    .S(_02184_),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_1 _26136_ (.A0(\M00r[11] ),
    .A1(\M00r[12] ),
    .S(_02184_),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _26137_ (.A0(_02243_),
    .A1(_02244_),
    .S(_02162_),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _26138_ (.A0(\M00r[12] ),
    .A1(\M00r[13] ),
    .S(_02184_),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _26139_ (.A0(_02246_),
    .A1(_02244_),
    .S(_02203_),
    .X(_02247_));
 sky130_fd_sc_hd__clkbuf_4 _26140_ (.A(_02165_),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _26141_ (.A0(_02245_),
    .A1(_02247_),
    .S(_02248_),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _26142_ (.A0(_02246_),
    .A1(_02202_),
    .S(_02162_),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _26143_ (.A0(_02247_),
    .A1(_02250_),
    .S(_02165_),
    .X(_02251_));
 sky130_fd_sc_hd__clkbuf_4 _26144_ (.A(_02154_),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _26145_ (.A0(_02249_),
    .A1(_02251_),
    .S(_02253_),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _26146_ (.A0(_02250_),
    .A1(_02204_),
    .S(_02165_),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _26147_ (.A0(_02251_),
    .A1(_02255_),
    .S(_02154_),
    .X(_02256_));
 sky130_fd_sc_hd__clkbuf_4 _26148_ (.A(_02157_),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _26149_ (.A0(_02254_),
    .A1(_02256_),
    .S(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _26150_ (.A0(_02255_),
    .A1(_02207_),
    .S(_02154_),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _26151_ (.A0(_02256_),
    .A1(_02259_),
    .S(_02157_),
    .X(_02260_));
 sky130_fd_sc_hd__clkbuf_4 _26152_ (.A(_02182_),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _26153_ (.A0(_02258_),
    .A1(_02260_),
    .S(_02261_),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _26154_ (.A0(_02259_),
    .A1(_02211_),
    .S(_02157_),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _26155_ (.A0(_02260_),
    .A1(_02264_),
    .S(_02182_),
    .X(_02265_));
 sky130_fd_sc_hd__clkbuf_4 _26156_ (.A(_02194_),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _26157_ (.A0(_02262_),
    .A1(_02265_),
    .S(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _26158_ (.A0(_02264_),
    .A1(_02214_),
    .S(_02182_),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _26159_ (.A0(_02265_),
    .A1(_02268_),
    .S(_02194_),
    .X(_02269_));
 sky130_fd_sc_hd__clkbuf_4 _26160_ (.A(_02198_),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _26161_ (.A0(_02267_),
    .A1(_02269_),
    .S(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _26162_ (.A0(_02268_),
    .A1(_02217_),
    .S(_02194_),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _26163_ (.A0(_02269_),
    .A1(_02272_),
    .S(_02198_),
    .X(_02273_));
 sky130_fd_sc_hd__clkbuf_4 _26164_ (.A(_02200_),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _26165_ (.A0(_02271_),
    .A1(_02273_),
    .S(_02275_),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _26166_ (.A0(_02272_),
    .A1(_02221_),
    .S(_02198_),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _26167_ (.A0(_02273_),
    .A1(_02277_),
    .S(_02200_),
    .X(_02278_));
 sky130_fd_sc_hd__clkbuf_4 _26168_ (.A(_02235_),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _26169_ (.A0(_02276_),
    .A1(_02278_),
    .S(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _26170_ (.A0(_02277_),
    .A1(_02224_),
    .S(_02200_),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _26171_ (.A0(_02278_),
    .A1(_02281_),
    .S(_02235_),
    .X(_02282_));
 sky130_fd_sc_hd__clkbuf_4 _26172_ (.A(_02238_),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _26173_ (.A0(_02280_),
    .A1(_02282_),
    .S(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__nand2_1 _26174_ (.A(_02231_),
    .B(_02235_),
    .Y(_02286_));
 sky130_fd_sc_hd__o21ai_1 _26175_ (.A1(_02235_),
    .A2(_02281_),
    .B1(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand2_1 _26176_ (.A(_02287_),
    .B(_02238_),
    .Y(_02288_));
 sky130_fd_sc_hd__o21ai_1 _26177_ (.A1(_02238_),
    .A2(_02282_),
    .B1(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__nand2_1 _26178_ (.A(_02289_),
    .B(_02240_),
    .Y(_02290_));
 sky130_fd_sc_hd__o21ai_1 _26179_ (.A1(_02242_),
    .A2(_02284_),
    .B1(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__mux2_1 _26180_ (.A0(_02287_),
    .A1(_02236_),
    .S(_02238_),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _26181_ (.A0(_02289_),
    .A1(_02292_),
    .S(_02240_),
    .X(_02293_));
 sky130_fd_sc_hd__clkinv_4 _26182_ (.A(_02240_),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_2 _26183_ (.A(_02292_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__mux2_1 _26184_ (.A0(_02291_),
    .A1(_02293_),
    .S(_02295_),
    .X(_02297_));
 sky130_fd_sc_hd__inv_4 _26185_ (.A(_02295_),
    .Y(_02298_));
 sky130_fd_sc_hd__nand2_1 _26186_ (.A(_02293_),
    .B(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__clkbuf_4 _26187_ (.A(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__inv_2 _26188_ (.A(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hd__nand2_1 _26189_ (.A(_02297_),
    .B(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hd__clkbuf_4 _26190_ (.A(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__buf_6 _26191_ (.A(_02184_),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _26192_ (.A0(\M00r[8] ),
    .A1(\M00r[9] ),
    .S(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _26193_ (.A0(net206),
    .A1(\M00r[8] ),
    .S(_02304_),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _26194_ (.A0(_02305_),
    .A1(_02306_),
    .S(_02203_),
    .X(_02308_));
 sky130_fd_sc_hd__mux2_1 _26195_ (.A0(\M00r[9] ),
    .A1(\M00r[10] ),
    .S(_02184_),
    .X(_02309_));
 sky130_fd_sc_hd__mux2_1 _26196_ (.A0(_02305_),
    .A1(_02309_),
    .S(_02162_),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _26197_ (.A0(_02308_),
    .A1(_02310_),
    .S(_02248_),
    .X(_02311_));
 sky130_fd_sc_hd__mux2_1 _26198_ (.A0(_02243_),
    .A1(_02309_),
    .S(_02203_),
    .X(_02312_));
 sky130_fd_sc_hd__mux2_1 _26199_ (.A0(_02310_),
    .A1(_02312_),
    .S(_02248_),
    .X(_02313_));
 sky130_fd_sc_hd__mux2_1 _26200_ (.A0(_02311_),
    .A1(_02313_),
    .S(_02253_),
    .X(_02314_));
 sky130_fd_sc_hd__mux2_1 _26201_ (.A0(_02312_),
    .A1(_02245_),
    .S(_02248_),
    .X(_02315_));
 sky130_fd_sc_hd__mux2_1 _26202_ (.A0(_02313_),
    .A1(_02315_),
    .S(_02253_),
    .X(_02316_));
 sky130_fd_sc_hd__mux2_1 _26203_ (.A0(_02314_),
    .A1(_02316_),
    .S(_02257_),
    .X(_02317_));
 sky130_fd_sc_hd__mux2_1 _26204_ (.A0(_02315_),
    .A1(_02249_),
    .S(_02253_),
    .X(_02319_));
 sky130_fd_sc_hd__mux2_1 _26205_ (.A0(_02316_),
    .A1(_02319_),
    .S(_02257_),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _26206_ (.A0(_02317_),
    .A1(_02320_),
    .S(_02261_),
    .X(_02321_));
 sky130_fd_sc_hd__mux2_1 _26207_ (.A0(_02319_),
    .A1(_02254_),
    .S(_02257_),
    .X(_02322_));
 sky130_fd_sc_hd__mux2_1 _26208_ (.A0(_02320_),
    .A1(_02322_),
    .S(_02261_),
    .X(_02323_));
 sky130_fd_sc_hd__mux2_1 _26209_ (.A0(_02321_),
    .A1(_02323_),
    .S(_02266_),
    .X(_02324_));
 sky130_fd_sc_hd__mux2_1 _26210_ (.A0(_02322_),
    .A1(_02258_),
    .S(_02261_),
    .X(_02325_));
 sky130_fd_sc_hd__mux2_1 _26211_ (.A0(_02323_),
    .A1(_02325_),
    .S(_02266_),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_1 _26212_ (.A0(_02324_),
    .A1(_02326_),
    .S(_02270_),
    .X(_02327_));
 sky130_fd_sc_hd__mux2_1 _26213_ (.A0(_02325_),
    .A1(_02262_),
    .S(_02266_),
    .X(_02328_));
 sky130_fd_sc_hd__mux2_1 _26214_ (.A0(_02326_),
    .A1(_02328_),
    .S(_02270_),
    .X(_02330_));
 sky130_fd_sc_hd__mux2_1 _26215_ (.A0(_02327_),
    .A1(_02330_),
    .S(_02275_),
    .X(_02331_));
 sky130_fd_sc_hd__mux2_1 _26216_ (.A0(_02328_),
    .A1(_02267_),
    .S(_02270_),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _26217_ (.A0(_02330_),
    .A1(_02332_),
    .S(_02275_),
    .X(_02333_));
 sky130_fd_sc_hd__mux2_1 _26218_ (.A0(_02331_),
    .A1(_02333_),
    .S(_02279_),
    .X(_02334_));
 sky130_fd_sc_hd__mux2_1 _26219_ (.A0(_02332_),
    .A1(_02271_),
    .S(_02275_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _26220_ (.A0(_02333_),
    .A1(_02335_),
    .S(_02279_),
    .X(_02336_));
 sky130_fd_sc_hd__mux2_1 _26221_ (.A0(_02334_),
    .A1(_02336_),
    .S(_02283_),
    .X(_02337_));
 sky130_fd_sc_hd__mux2_1 _26222_ (.A0(_02335_),
    .A1(_02276_),
    .S(_02279_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _26223_ (.A0(_02336_),
    .A1(_02338_),
    .S(_02283_),
    .X(_02339_));
 sky130_fd_sc_hd__mux2_1 _26224_ (.A0(_02337_),
    .A1(_02339_),
    .S(_02242_),
    .X(_02341_));
 sky130_fd_sc_hd__mux2_1 _26225_ (.A0(_02338_),
    .A1(_02280_),
    .S(_02283_),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _26226_ (.A0(_02339_),
    .A1(_02342_),
    .S(_02242_),
    .X(_02343_));
 sky130_fd_sc_hd__clkbuf_4 _26227_ (.A(_02295_),
    .X(_02344_));
 sky130_fd_sc_hd__mux2_1 _26228_ (.A0(_02341_),
    .A1(_02343_),
    .S(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__mux2_1 _26229_ (.A0(_02342_),
    .A1(_02284_),
    .S(_02240_),
    .X(_02346_));
 sky130_fd_sc_hd__mux2_1 _26230_ (.A0(_02343_),
    .A1(_02346_),
    .S(_02344_),
    .X(_02347_));
 sky130_fd_sc_hd__mux2_1 _26231_ (.A0(_02345_),
    .A1(_02347_),
    .S(_02300_),
    .X(_02348_));
 sky130_fd_sc_hd__inv_4 _26232_ (.A(_02302_),
    .Y(_02349_));
 sky130_fd_sc_hd__nand2_1 _26233_ (.A(_02291_),
    .B(_02295_),
    .Y(_02350_));
 sky130_fd_sc_hd__o21ai_1 _26234_ (.A1(_02344_),
    .A2(_02346_),
    .B1(_02350_),
    .Y(_02352_));
 sky130_fd_sc_hd__nand2_1 _26235_ (.A(_02347_),
    .B(_02301_),
    .Y(_02353_));
 sky130_fd_sc_hd__o21ai_1 _26236_ (.A1(_02301_),
    .A2(_02352_),
    .B1(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__or2_1 _26237_ (.A(_02349_),
    .B(_02354_),
    .X(_02355_));
 sky130_fd_sc_hd__o21ai_1 _26238_ (.A1(_02303_),
    .A2(_02348_),
    .B1(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__mux2_1 _26239_ (.A0(_02352_),
    .A1(_02297_),
    .S(_02300_),
    .X(_02357_));
 sky130_fd_sc_hd__nand2_1 _26240_ (.A(_02357_),
    .B(_02303_),
    .Y(_02358_));
 sky130_fd_sc_hd__o21ai_1 _26241_ (.A1(_02303_),
    .A2(_02354_),
    .B1(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hd__nand2_1 _26242_ (.A(_02357_),
    .B(_02349_),
    .Y(_02360_));
 sky130_fd_sc_hd__mux2_1 _26243_ (.A0(_02356_),
    .A1(_02359_),
    .S(_02360_),
    .X(_02361_));
 sky130_fd_sc_hd__inv_1 _26244_ (.A(_02360_),
    .Y(_02363_));
 sky130_fd_sc_hd__nand2_1 _26245_ (.A(_02359_),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hd__inv_2 _26246_ (.A(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__nand2_1 _26247_ (.A(_02361_),
    .B(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__buf_6 _26248_ (.A(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__mux2_1 _26249_ (.A0(\M00r[4] ),
    .A1(net191),
    .S(_02304_),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _26250_ (.A0(net191),
    .A1(\M00r[6] ),
    .S(_02304_),
    .X(_02369_));
 sky130_fd_sc_hd__mux2_1 _26251_ (.A0(net192),
    .A1(_02369_),
    .S(_02162_),
    .X(_02370_));
 sky130_fd_sc_hd__mux2_1 _26252_ (.A0(\M00r[6] ),
    .A1(net206),
    .S(_02304_),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _26253_ (.A0(net207),
    .A1(_02369_),
    .S(_02203_),
    .X(_02372_));
 sky130_fd_sc_hd__mux2_1 _26254_ (.A0(_02370_),
    .A1(net208),
    .S(_02248_),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _26255_ (.A0(_02371_),
    .A1(_02306_),
    .S(_02162_),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _26256_ (.A0(_02372_),
    .A1(_02375_),
    .S(_02248_),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _26257_ (.A0(_02374_),
    .A1(_02376_),
    .S(_02253_),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _26258_ (.A0(_02375_),
    .A1(_02308_),
    .S(_02248_),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _26259_ (.A0(_02376_),
    .A1(_02378_),
    .S(_02253_),
    .X(_02379_));
 sky130_fd_sc_hd__mux2_1 _26260_ (.A0(_02377_),
    .A1(_02379_),
    .S(_02257_),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _26261_ (.A0(_02378_),
    .A1(_02311_),
    .S(_02253_),
    .X(_02381_));
 sky130_fd_sc_hd__mux2_1 _26262_ (.A0(_02379_),
    .A1(_02381_),
    .S(_02257_),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _26263_ (.A0(_02380_),
    .A1(_02382_),
    .S(_02261_),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _26264_ (.A0(_02381_),
    .A1(_02314_),
    .S(_02257_),
    .X(_02385_));
 sky130_fd_sc_hd__mux2_1 _26265_ (.A0(_02382_),
    .A1(_02385_),
    .S(_02261_),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _26266_ (.A0(_02383_),
    .A1(_02386_),
    .S(_02266_),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_1 _26267_ (.A0(_02385_),
    .A1(_02317_),
    .S(_02261_),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _26268_ (.A0(_02386_),
    .A1(_02388_),
    .S(_02266_),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _26269_ (.A0(_02387_),
    .A1(_02389_),
    .S(_02270_),
    .X(_02390_));
 sky130_fd_sc_hd__mux2_1 _26270_ (.A0(_02388_),
    .A1(_02321_),
    .S(_02266_),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _26271_ (.A0(_02389_),
    .A1(_02391_),
    .S(_02270_),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _26272_ (.A0(_02390_),
    .A1(_02392_),
    .S(_02275_),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _26273_ (.A0(_02391_),
    .A1(_02324_),
    .S(_02270_),
    .X(_02394_));
 sky130_fd_sc_hd__mux2_1 _26274_ (.A0(_02392_),
    .A1(_02394_),
    .S(_02275_),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _26275_ (.A0(_02393_),
    .A1(_02396_),
    .S(_02279_),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _26276_ (.A0(_02394_),
    .A1(_02327_),
    .S(_02275_),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _26277_ (.A0(_02396_),
    .A1(_02398_),
    .S(_02279_),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _26278_ (.A0(_02397_),
    .A1(_02399_),
    .S(_02283_),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _26279_ (.A0(_02398_),
    .A1(_02331_),
    .S(_02279_),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _26280_ (.A0(_02399_),
    .A1(_02401_),
    .S(_02283_),
    .X(_02402_));
 sky130_fd_sc_hd__mux2_1 _26281_ (.A0(_02400_),
    .A1(_02402_),
    .S(_02242_),
    .X(_02403_));
 sky130_fd_sc_hd__mux2_1 _26282_ (.A0(_02401_),
    .A1(_02334_),
    .S(_02283_),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _26283_ (.A0(_02402_),
    .A1(_02404_),
    .S(_02242_),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _26284_ (.A0(_02403_),
    .A1(_02405_),
    .S(_02344_),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _26285_ (.A0(_02404_),
    .A1(_02337_),
    .S(_02242_),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _26286_ (.A0(_02405_),
    .A1(_02408_),
    .S(_02344_),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _26287_ (.A0(_02407_),
    .A1(_02409_),
    .S(_02300_),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _26288_ (.A0(_02408_),
    .A1(_02341_),
    .S(_02344_),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _26289_ (.A0(_02409_),
    .A1(_02411_),
    .S(_02300_),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _26290_ (.A0(_02410_),
    .A1(_02412_),
    .S(_02303_),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _26291_ (.A0(_02411_),
    .A1(_02345_),
    .S(_02300_),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _26292_ (.A0(_02412_),
    .A1(_02414_),
    .S(_02303_),
    .X(_02415_));
 sky130_fd_sc_hd__clkbuf_4 _26293_ (.A(_02360_),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _26294_ (.A0(_02413_),
    .A1(_02415_),
    .S(_02416_),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _26295_ (.A0(_02414_),
    .A1(_02348_),
    .S(_02303_),
    .X(_02419_));
 sky130_fd_sc_hd__mux2_1 _26296_ (.A0(_02415_),
    .A1(_02419_),
    .S(_02416_),
    .X(_02420_));
 sky130_fd_sc_hd__buf_6 _26297_ (.A(_02364_),
    .X(_02421_));
 sky130_fd_sc_hd__mux2_1 _26298_ (.A0(_02418_),
    .A1(_02420_),
    .S(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__nand2_1 _26299_ (.A(_02356_),
    .B(_02416_),
    .Y(_02423_));
 sky130_fd_sc_hd__o21ai_1 _26300_ (.A1(_02416_),
    .A2(_02419_),
    .B1(_02423_),
    .Y(_02424_));
 sky130_fd_sc_hd__nand2_1 _26301_ (.A(_02424_),
    .B(_02421_),
    .Y(_02425_));
 sky130_fd_sc_hd__o21ai_1 _26302_ (.A1(_02421_),
    .A2(_02420_),
    .B1(_02425_),
    .Y(_02426_));
 sky130_fd_sc_hd__nand2_1 _26303_ (.A(_02426_),
    .B(_02367_),
    .Y(_02427_));
 sky130_fd_sc_hd__o21ai_1 _26304_ (.A1(_02367_),
    .A2(_02422_),
    .B1(_02427_),
    .Y(_02429_));
 sky130_fd_sc_hd__mux2_1 _26305_ (.A0(_02361_),
    .A1(_02424_),
    .S(_02365_),
    .X(_02430_));
 sky130_fd_sc_hd__mux2_1 _26306_ (.A0(_02426_),
    .A1(_02430_),
    .S(_02367_),
    .X(_02431_));
 sky130_fd_sc_hd__inv_2 _26307_ (.A(_02366_),
    .Y(_02432_));
 sky130_fd_sc_hd__nand2_4 _26308_ (.A(_02430_),
    .B(_02432_),
    .Y(_02433_));
 sky130_fd_sc_hd__mux2_1 _26309_ (.A0(_02429_),
    .A1(_02431_),
    .S(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__inv_2 _26310_ (.A(_02433_),
    .Y(_02435_));
 sky130_fd_sc_hd__nand2_4 _26311_ (.A(_02431_),
    .B(_02435_),
    .Y(_02436_));
 sky130_fd_sc_hd__inv_2 _26312_ (.A(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__nand2_2 _26313_ (.A(_02434_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__mux2_1 _26314_ (.A0(net171),
    .A1(net217),
    .S(_02304_),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _26315_ (.A0(net187),
    .A1(net171),
    .S(_02304_),
    .X(_02441_));
 sky130_fd_sc_hd__mux2_1 _26316_ (.A0(net218),
    .A1(net172),
    .S(_02203_),
    .X(_02442_));
 sky130_fd_sc_hd__mux2_1 _26317_ (.A0(\M00r[3] ),
    .A1(\M00r[4] ),
    .S(_02304_),
    .X(_02443_));
 sky130_fd_sc_hd__mux2_1 _26318_ (.A0(_02440_),
    .A1(_02443_),
    .S(_02162_),
    .X(_02444_));
 sky130_fd_sc_hd__mux2_1 _26319_ (.A0(_02442_),
    .A1(_02444_),
    .S(_02248_),
    .X(_02445_));
 sky130_fd_sc_hd__mux2_1 _26320_ (.A0(net192),
    .A1(_02443_),
    .S(_02203_),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _26321_ (.A0(_02444_),
    .A1(net193),
    .S(_02248_),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _26322_ (.A0(_02445_),
    .A1(net194),
    .S(_02253_),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _26323_ (.A0(net193),
    .A1(_02370_),
    .S(_02248_),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _26324_ (.A0(net194),
    .A1(_02449_),
    .S(_02253_),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _26325_ (.A0(net195),
    .A1(_02451_),
    .S(_02257_),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _26326_ (.A0(_02449_),
    .A1(net209),
    .S(_02253_),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _26327_ (.A0(_02451_),
    .A1(net210),
    .S(_02257_),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _26328_ (.A0(_02452_),
    .A1(net211),
    .S(_02261_),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _26329_ (.A0(_02453_),
    .A1(_02377_),
    .S(_02257_),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _26330_ (.A0(_02454_),
    .A1(_02456_),
    .S(_02261_),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _26331_ (.A0(_02455_),
    .A1(_02457_),
    .S(_02266_),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _26332_ (.A0(_02456_),
    .A1(_02380_),
    .S(_02261_),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _26333_ (.A0(_02457_),
    .A1(_02459_),
    .S(_02266_),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _26334_ (.A0(_02458_),
    .A1(_02460_),
    .S(_02270_),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _26335_ (.A0(_02459_),
    .A1(_02383_),
    .S(_02266_),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _26336_ (.A0(_02460_),
    .A1(_02463_),
    .S(_02270_),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _26337_ (.A0(_02462_),
    .A1(_02464_),
    .S(_02275_),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _26338_ (.A0(_02463_),
    .A1(_02387_),
    .S(_02270_),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _26339_ (.A0(_02464_),
    .A1(_02466_),
    .S(_02275_),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _26340_ (.A0(_02465_),
    .A1(_02467_),
    .S(_02279_),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _26341_ (.A0(_02466_),
    .A1(_02390_),
    .S(_02275_),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _26342_ (.A0(_02467_),
    .A1(_02469_),
    .S(_02279_),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _26343_ (.A0(_02468_),
    .A1(_02470_),
    .S(_02283_),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _26344_ (.A0(_02469_),
    .A1(_02393_),
    .S(_02279_),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _26345_ (.A0(_02470_),
    .A1(_02473_),
    .S(_02283_),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _26346_ (.A0(_02471_),
    .A1(_02474_),
    .S(_02242_),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _26347_ (.A0(_02473_),
    .A1(_02397_),
    .S(_02283_),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _26348_ (.A0(_02474_),
    .A1(_02476_),
    .S(_02242_),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _26349_ (.A0(_02475_),
    .A1(_02477_),
    .S(_02344_),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _26350_ (.A0(_02476_),
    .A1(_02400_),
    .S(_02242_),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _26351_ (.A0(_02477_),
    .A1(_02479_),
    .S(_02344_),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _26352_ (.A0(_02478_),
    .A1(_02480_),
    .S(_02300_),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _26353_ (.A0(_02479_),
    .A1(_02403_),
    .S(_02344_),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _26354_ (.A0(_02480_),
    .A1(_02482_),
    .S(_02300_),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _26355_ (.A0(_02481_),
    .A1(_02484_),
    .S(_02303_),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _26356_ (.A0(_02482_),
    .A1(_02407_),
    .S(_02300_),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _26357_ (.A0(_02484_),
    .A1(_02486_),
    .S(_02303_),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _26358_ (.A0(_02485_),
    .A1(_02487_),
    .S(_02416_),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _26359_ (.A0(_02486_),
    .A1(_02410_),
    .S(_02303_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _26360_ (.A0(_02487_),
    .A1(_02489_),
    .S(_02416_),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _26361_ (.A0(_02488_),
    .A1(_02490_),
    .S(_02421_),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _26362_ (.A0(_02489_),
    .A1(_02413_),
    .S(_02416_),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _26363_ (.A0(_02490_),
    .A1(_02492_),
    .S(_02421_),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _26364_ (.A0(_02491_),
    .A1(_02493_),
    .S(_02367_),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _26365_ (.A0(_02492_),
    .A1(_02418_),
    .S(_02421_),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _26366_ (.A0(_02493_),
    .A1(_02496_),
    .S(_02367_),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _26367_ (.A0(_02495_),
    .A1(_02497_),
    .S(_02433_),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _26368_ (.A0(_02496_),
    .A1(_02422_),
    .S(_02367_),
    .X(_02499_));
 sky130_fd_sc_hd__mux2_1 _26369_ (.A0(_02497_),
    .A1(_02499_),
    .S(_02433_),
    .X(_02500_));
 sky130_fd_sc_hd__mux2_1 _26370_ (.A0(_02498_),
    .A1(_02500_),
    .S(_02436_),
    .X(_02501_));
 sky130_fd_sc_hd__nand2_1 _26371_ (.A(_02429_),
    .B(_02433_),
    .Y(_02502_));
 sky130_fd_sc_hd__o21ai_1 _26372_ (.A1(_02433_),
    .A2(_02499_),
    .B1(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__nand2_1 _26373_ (.A(_02503_),
    .B(_02436_),
    .Y(_02504_));
 sky130_fd_sc_hd__o21ai_1 _26374_ (.A1(_02436_),
    .A2(_02500_),
    .B1(_02504_),
    .Y(_02506_));
 sky130_fd_sc_hd__nand2_1 _26375_ (.A(_02506_),
    .B(_02438_),
    .Y(_02507_));
 sky130_fd_sc_hd__o21ai_1 _26376_ (.A1(_02438_),
    .A2(_02501_),
    .B1(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hd__mux2_1 _26377_ (.A0(_02503_),
    .A1(_02434_),
    .S(_02436_),
    .X(_02509_));
 sky130_fd_sc_hd__mux2_1 _26378_ (.A0(_02506_),
    .A1(_02509_),
    .S(_02438_),
    .X(_02510_));
 sky130_fd_sc_hd__inv_2 _26379_ (.A(_02438_),
    .Y(_02511_));
 sky130_fd_sc_hd__nand2_2 _26380_ (.A(_02509_),
    .B(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__mux2_1 _26381_ (.A0(_02508_),
    .A1(_02510_),
    .S(_02512_),
    .X(_02513_));
 sky130_fd_sc_hd__inv_2 _26382_ (.A(_02512_),
    .Y(_02514_));
 sky130_fd_sc_hd__or2_1 _26383_ (.A(_02437_),
    .B(_02498_),
    .X(_02515_));
 sky130_fd_sc_hd__or2_1 _26384_ (.A(_02349_),
    .B(_02481_),
    .X(_02517_));
 sky130_fd_sc_hd__or2_1 _26385_ (.A(net187),
    .B(_02146_),
    .X(_02518_));
 sky130_fd_sc_hd__o21a_1 _26386_ (.A1(_02304_),
    .A2(net167),
    .B1(net188),
    .X(_02519_));
 sky130_fd_sc_hd__mux2_1 _26387_ (.A0(net172),
    .A1(_02519_),
    .S(_02203_),
    .X(_02520_));
 sky130_fd_sc_hd__mux2_1 _26388_ (.A0(_02442_),
    .A1(net173),
    .S(_02152_),
    .X(_02521_));
 sky130_fd_sc_hd__inv_2 _26389_ (.A(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__nand2_1 _26390_ (.A(_02522_),
    .B(_02155_),
    .Y(_02523_));
 sky130_fd_sc_hd__o21ai_1 _26391_ (.A1(_02155_),
    .A2(_02445_),
    .B1(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__nand2_1 _26392_ (.A(_02524_),
    .B(_02170_),
    .Y(_02525_));
 sky130_fd_sc_hd__o21ai_1 _26393_ (.A1(_02170_),
    .A2(net195),
    .B1(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__nand2_1 _26394_ (.A(net196),
    .B(_02193_),
    .Y(_02528_));
 sky130_fd_sc_hd__o21ai_1 _26395_ (.A1(_02193_),
    .A2(_02452_),
    .B1(net197),
    .Y(_02529_));
 sky130_fd_sc_hd__nand2_1 _26396_ (.A(net198),
    .B(_02195_),
    .Y(_02530_));
 sky130_fd_sc_hd__o21ai_2 _26397_ (.A1(_02195_),
    .A2(net212),
    .B1(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__nand2_1 _26398_ (.A(_02531_),
    .B(_02199_),
    .Y(_02532_));
 sky130_fd_sc_hd__o21ai_1 _26399_ (.A1(_02199_),
    .A2(_02458_),
    .B1(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__nand2_1 _26400_ (.A(_02533_),
    .B(_02234_),
    .Y(_02534_));
 sky130_fd_sc_hd__o21ai_2 _26401_ (.A1(_02234_),
    .A2(_02462_),
    .B1(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__nand2_1 _26402_ (.A(_02535_),
    .B(_02237_),
    .Y(_02536_));
 sky130_fd_sc_hd__o21ai_2 _26403_ (.A1(_02237_),
    .A2(_02465_),
    .B1(_02536_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2_1 _26404_ (.A(_02537_),
    .B(_02239_),
    .Y(_02539_));
 sky130_fd_sc_hd__o21ai_2 _26405_ (.A1(_02239_),
    .A2(_02468_),
    .B1(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__nand2_1 _26406_ (.A(_02540_),
    .B(_02294_),
    .Y(_02541_));
 sky130_fd_sc_hd__o21ai_2 _26407_ (.A1(_02294_),
    .A2(_02471_),
    .B1(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_1 _26408_ (.A(_02542_),
    .B(_02298_),
    .Y(_02543_));
 sky130_fd_sc_hd__o21ai_2 _26409_ (.A1(_02298_),
    .A2(_02475_),
    .B1(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__nand2_1 _26410_ (.A(_02544_),
    .B(_02301_),
    .Y(_02545_));
 sky130_fd_sc_hd__o21ai_2 _26411_ (.A1(_02301_),
    .A2(_02478_),
    .B1(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__nand2_1 _26412_ (.A(_02546_),
    .B(_02349_),
    .Y(_02547_));
 sky130_fd_sc_hd__nand2_2 _26413_ (.A(_02517_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__nand2_1 _26414_ (.A(_02485_),
    .B(_02416_),
    .Y(_02550_));
 sky130_fd_sc_hd__o21ai_2 _26415_ (.A1(_02416_),
    .A2(_02548_),
    .B1(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__mux2_1 _26416_ (.A0(_02488_),
    .A1(_02551_),
    .S(_02365_),
    .X(_02552_));
 sky130_fd_sc_hd__mux2_1 _26417_ (.A0(_02491_),
    .A1(_02552_),
    .S(_02432_),
    .X(_02553_));
 sky130_fd_sc_hd__mux2_1 _26418_ (.A0(_02495_),
    .A1(_02553_),
    .S(_02435_),
    .X(_02554_));
 sky130_fd_sc_hd__or2_1 _26419_ (.A(_02436_),
    .B(_02554_),
    .X(_02555_));
 sky130_fd_sc_hd__nand2_1 _26420_ (.A(_02515_),
    .B(_02555_),
    .Y(_02556_));
 sky130_fd_sc_hd__nand2_1 _26421_ (.A(_02501_),
    .B(_02438_),
    .Y(_02557_));
 sky130_fd_sc_hd__o21ai_1 _26422_ (.A1(_02438_),
    .A2(_02556_),
    .B1(_02557_),
    .Y(_02558_));
 sky130_fd_sc_hd__nand2_1 _26423_ (.A(_02558_),
    .B(_02514_),
    .Y(_02559_));
 sky130_fd_sc_hd__o21ai_1 _26424_ (.A1(_02514_),
    .A2(_02508_),
    .B1(_02559_),
    .Y(_02561_));
 sky130_fd_sc_hd__inv_2 _26425_ (.A(_02561_),
    .Y(_02562_));
 sky130_fd_sc_hd__nand2_1 _26426_ (.A(_02510_),
    .B(_02514_),
    .Y(_02563_));
 sky130_fd_sc_hd__clkinvlp_2 _26427_ (.A(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__mux2_1 _26428_ (.A0(_02513_),
    .A1(_02562_),
    .S(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__nand2_1 _26429_ (.A(_02513_),
    .B(_02564_),
    .Y(_02566_));
 sky130_fd_sc_hd__clkinvlp_2 _26430_ (.A(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__nand2_1 _26431_ (.A(_02565_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__inv_2 _26432_ (.A(net16),
    .Y(_02569_));
 sky130_fd_sc_hd__nand2_1 _26433_ (.A(_07088_),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__nand2_1 _26434_ (.A(_08790_),
    .B(net16),
    .Y(_02572_));
 sky130_fd_sc_hd__nand2_1 _26435_ (.A(_02570_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__or2_2 _26436_ (.A(net48),
    .B(_02573_),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_1 _26437_ (.A(_02573_),
    .B(net48),
    .Y(_02575_));
 sky130_fd_sc_hd__nand2_4 _26438_ (.A(_02574_),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__inv_2 _26439_ (.A(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_1 _26440_ (.A(_02577_),
    .B(\M00r[24] ),
    .Y(_02578_));
 sky130_fd_sc_hd__nand2_1 _26441_ (.A(_02576_),
    .B(_02146_),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _26442_ (.A(_02578_),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__xor2_1 _26443_ (.A(_02138_),
    .B(_02580_),
    .X(_02581_));
 sky130_fd_sc_hd__or2_1 _26444_ (.A(_02150_),
    .B(_02581_),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_1 _26445_ (.A(_02581_),
    .B(_02150_),
    .Y(_02584_));
 sky130_fd_sc_hd__and2_1 _26446_ (.A(_02583_),
    .B(_02584_),
    .X(_02585_));
 sky130_fd_sc_hd__or2_1 _26447_ (.A(_02155_),
    .B(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__nand2_1 _26448_ (.A(_02585_),
    .B(_02155_),
    .Y(_02587_));
 sky130_fd_sc_hd__nand2_1 _26449_ (.A(_02586_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__inv_2 _26450_ (.A(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__nand2_1 _26451_ (.A(_02589_),
    .B(_02156_),
    .Y(_02590_));
 sky130_fd_sc_hd__nand2_1 _26452_ (.A(_02588_),
    .B(_02170_),
    .Y(_02591_));
 sky130_fd_sc_hd__nand2_1 _26453_ (.A(_02590_),
    .B(_02591_),
    .Y(_02592_));
 sky130_fd_sc_hd__xor2_1 _26454_ (.A(_02193_),
    .B(_02592_),
    .X(_02594_));
 sky130_fd_sc_hd__xor2_1 _26455_ (.A(_02194_),
    .B(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__inv_2 _26456_ (.A(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__nand2_1 _26457_ (.A(_02596_),
    .B(_02199_),
    .Y(_02597_));
 sky130_fd_sc_hd__nand2_1 _26458_ (.A(_02595_),
    .B(_02198_),
    .Y(_02598_));
 sky130_fd_sc_hd__nand2_1 _26459_ (.A(_02597_),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__or2_1 _26460_ (.A(_02200_),
    .B(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__nand2_1 _26461_ (.A(_02599_),
    .B(_02200_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand2_1 _26462_ (.A(_02600_),
    .B(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__or2_1 _26463_ (.A(_02235_),
    .B(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__nand2_1 _26464_ (.A(_02602_),
    .B(_02235_),
    .Y(_02605_));
 sky130_fd_sc_hd__and2_1 _26465_ (.A(_02603_),
    .B(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__or2_1 _26466_ (.A(_02239_),
    .B(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__nand2_1 _26467_ (.A(_02606_),
    .B(_02239_),
    .Y(_02608_));
 sky130_fd_sc_hd__nand2_1 _26468_ (.A(_02607_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__or2_1 _26469_ (.A(_02240_),
    .B(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__nand2_1 _26470_ (.A(_02609_),
    .B(_02240_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand2_1 _26471_ (.A(_02610_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__or2_1 _26472_ (.A(_02295_),
    .B(_02612_),
    .X(_02613_));
 sky130_fd_sc_hd__nand2_1 _26473_ (.A(_02612_),
    .B(_02295_),
    .Y(_02614_));
 sky130_fd_sc_hd__nand2_1 _26474_ (.A(_02613_),
    .B(_02614_),
    .Y(_02616_));
 sky130_fd_sc_hd__or2_1 _26475_ (.A(_02299_),
    .B(_02616_),
    .X(_02617_));
 sky130_fd_sc_hd__nand2_1 _26476_ (.A(_02616_),
    .B(_02300_),
    .Y(_02618_));
 sky130_fd_sc_hd__nand2_1 _26477_ (.A(_02617_),
    .B(_02618_),
    .Y(_02619_));
 sky130_fd_sc_hd__or2_1 _26478_ (.A(_02302_),
    .B(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__nand2_1 _26479_ (.A(_02619_),
    .B(_02303_),
    .Y(_02621_));
 sky130_fd_sc_hd__nand2_1 _26480_ (.A(_02620_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__xor2_1 _26481_ (.A(_02416_),
    .B(_02622_),
    .X(_02623_));
 sky130_fd_sc_hd__xor2_1 _26482_ (.A(_02421_),
    .B(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__or2_1 _26483_ (.A(_02367_),
    .B(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__nand2_1 _26484_ (.A(_02624_),
    .B(_02367_),
    .Y(_02627_));
 sky130_fd_sc_hd__nand2_1 _26485_ (.A(_02625_),
    .B(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__or2_1 _26486_ (.A(_02433_),
    .B(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__nand2_1 _26487_ (.A(_02628_),
    .B(_02433_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2_1 _26488_ (.A(_02629_),
    .B(_02630_),
    .Y(_02631_));
 sky130_fd_sc_hd__or2_1 _26489_ (.A(_02436_),
    .B(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__nand2_1 _26490_ (.A(_02631_),
    .B(_02436_),
    .Y(_02633_));
 sky130_fd_sc_hd__nand2_1 _26491_ (.A(_02632_),
    .B(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__or2_1 _26492_ (.A(_02438_),
    .B(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__nand2_1 _26493_ (.A(_02634_),
    .B(_02438_),
    .Y(_02636_));
 sky130_fd_sc_hd__nand2_1 _26494_ (.A(_02635_),
    .B(_02636_),
    .Y(_02638_));
 sky130_fd_sc_hd__or2_1 _26495_ (.A(_02512_),
    .B(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__nand2_1 _26496_ (.A(_02638_),
    .B(_02512_),
    .Y(_02640_));
 sky130_fd_sc_hd__nand2_1 _26497_ (.A(_02639_),
    .B(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__or2_1 _26498_ (.A(_02563_),
    .B(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__nand2_1 _26499_ (.A(_02641_),
    .B(_02563_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_1 _26500_ (.A(_02642_),
    .B(_02643_),
    .Y(_02644_));
 sky130_fd_sc_hd__or2_1 _26501_ (.A(_02566_),
    .B(_02644_),
    .X(_02645_));
 sky130_fd_sc_hd__nand2_1 _26502_ (.A(_02644_),
    .B(_02566_),
    .Y(_02646_));
 sky130_fd_sc_hd__nand2_1 _26503_ (.A(_02645_),
    .B(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__or2_1 _26504_ (.A(_02568_),
    .B(_02647_),
    .X(_02649_));
 sky130_fd_sc_hd__nand2_1 _26505_ (.A(_02647_),
    .B(_02568_),
    .Y(_02650_));
 sky130_fd_sc_hd__nand2_1 _26506_ (.A(_02649_),
    .B(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__buf_6 _26507_ (.A(net160),
    .X(_02652_));
 sky130_fd_sc_hd__inv_2 _26508_ (.A(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__nand2_1 _26509_ (.A(net160),
    .B(net153),
    .Y(_02654_));
 sky130_fd_sc_hd__inv_2 _26510_ (.A(net154),
    .Y(_02655_));
 sky130_fd_sc_hd__a21o_1 _26511_ (.A1(_02651_),
    .A2(_02653_),
    .B1(_02655_),
    .X(_00018_));
 sky130_fd_sc_hd__inv_2 _26512_ (.A(_02622_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2_1 _26513_ (.A(_02619_),
    .B(_02363_),
    .Y(_02657_));
 sky130_fd_sc_hd__inv_2 _26514_ (.A(_02597_),
    .Y(_02659_));
 sky130_fd_sc_hd__inv_2 _26515_ (.A(_02592_),
    .Y(_02660_));
 sky130_fd_sc_hd__nand2_1 _26516_ (.A(_02660_),
    .B(_02195_),
    .Y(_02661_));
 sky130_fd_sc_hd__inv_2 _26517_ (.A(net17),
    .Y(_02662_));
 sky130_fd_sc_hd__or2_1 _26518_ (.A(_02662_),
    .B(_02572_),
    .X(_02663_));
 sky130_fd_sc_hd__nand2_1 _26519_ (.A(_02572_),
    .B(_02662_),
    .Y(_02664_));
 sky130_fd_sc_hd__nand2_1 _26520_ (.A(_02663_),
    .B(_02664_),
    .Y(_02665_));
 sky130_fd_sc_hd__or2_1 _26521_ (.A(net49),
    .B(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__nand2_1 _26522_ (.A(_02665_),
    .B(net49),
    .Y(_02667_));
 sky130_fd_sc_hd__nand2_1 _26523_ (.A(_02666_),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__or2_2 _26524_ (.A(_02574_),
    .B(_02668_),
    .X(_02670_));
 sky130_fd_sc_hd__nand2_1 _26525_ (.A(_02668_),
    .B(_02574_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand2_4 _26526_ (.A(_02670_),
    .B(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__nor2_1 _26527_ (.A(_02576_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__nor2_1 _26528_ (.A(_02138_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__nand2_1 _26529_ (.A(_02672_),
    .B(_02576_),
    .Y(_02675_));
 sky130_fd_sc_hd__or2_1 _26530_ (.A(_02578_),
    .B(_02672_),
    .X(_02676_));
 sky130_fd_sc_hd__nand2_1 _26531_ (.A(_02672_),
    .B(_02578_),
    .Y(_02677_));
 sky130_fd_sc_hd__nand2_1 _26532_ (.A(_02676_),
    .B(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hd__a22o_1 _26533_ (.A1(_02674_),
    .A2(_02675_),
    .B1(_02678_),
    .B2(_02138_),
    .X(_02679_));
 sky130_fd_sc_hd__or2_1 _26534_ (.A(_02583_),
    .B(_02679_),
    .X(_02681_));
 sky130_fd_sc_hd__nand2_1 _26535_ (.A(_02679_),
    .B(_02583_),
    .Y(_02682_));
 sky130_fd_sc_hd__nand2_1 _26536_ (.A(_02681_),
    .B(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__nor2_1 _26537_ (.A(_02587_),
    .B(_02679_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21o_1 _26538_ (.A1(_02683_),
    .A2(_02587_),
    .B1(_02684_),
    .X(_02685_));
 sky130_fd_sc_hd__nand2_1 _26539_ (.A(_02589_),
    .B(_02170_),
    .Y(_02686_));
 sky130_fd_sc_hd__a21oi_1 _26540_ (.A1(_02683_),
    .A2(_02587_),
    .B1(_02686_),
    .Y(_02687_));
 sky130_fd_sc_hd__a21oi_1 _26541_ (.A1(_02685_),
    .A2(_02686_),
    .B1(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__inv_2 _26542_ (.A(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__or3_1 _26543_ (.A(_02181_),
    .B(_02589_),
    .C(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__o21ai_1 _26544_ (.A1(_02182_),
    .A2(_02589_),
    .B1(_02689_),
    .Y(_02692_));
 sky130_fd_sc_hd__nand2_1 _26545_ (.A(_02690_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__or2_1 _26546_ (.A(_02661_),
    .B(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__nand2_1 _26547_ (.A(_02693_),
    .B(_02661_),
    .Y(_02695_));
 sky130_fd_sc_hd__and2_1 _26548_ (.A(_02694_),
    .B(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__or2_1 _26549_ (.A(_02659_),
    .B(_02696_),
    .X(_02697_));
 sky130_fd_sc_hd__nand2_1 _26550_ (.A(_02696_),
    .B(_02659_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_1 _26551_ (.A(_02697_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__xor2_1 _26552_ (.A(_02600_),
    .B(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__inv_2 _26553_ (.A(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__nor3_1 _26554_ (.A(_02235_),
    .B(_02602_),
    .C(_02701_),
    .Y(_02703_));
 sky130_fd_sc_hd__a21oi_1 _26555_ (.A1(_02603_),
    .A2(_02701_),
    .B1(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__or2b_1 _26556_ (.A(_02704_),
    .B_N(_02608_),
    .X(_02705_));
 sky130_fd_sc_hd__nand3_1 _26557_ (.A(_02704_),
    .B(_02239_),
    .C(_02606_),
    .Y(_02706_));
 sky130_fd_sc_hd__nand2_1 _26558_ (.A(_02705_),
    .B(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__nor2_1 _26559_ (.A(_02610_),
    .B(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__inv_2 _26560_ (.A(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__nand2_1 _26561_ (.A(_02707_),
    .B(_02610_),
    .Y(_02710_));
 sky130_fd_sc_hd__nand2_1 _26562_ (.A(_02709_),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__inv_2 _26563_ (.A(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__inv_2 _26564_ (.A(_02613_),
    .Y(_02714_));
 sky130_fd_sc_hd__nand2_1 _26565_ (.A(_02712_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand2_1 _26566_ (.A(_02711_),
    .B(_02613_),
    .Y(_02716_));
 sky130_fd_sc_hd__nand2_1 _26567_ (.A(_02715_),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__or2_1 _26568_ (.A(_02617_),
    .B(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__nand2_1 _26569_ (.A(_02717_),
    .B(_02617_),
    .Y(_02719_));
 sky130_fd_sc_hd__nand2_1 _26570_ (.A(_02718_),
    .B(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__or2_1 _26571_ (.A(_02620_),
    .B(_02720_),
    .X(_02721_));
 sky130_fd_sc_hd__nand2_1 _26572_ (.A(_02720_),
    .B(_02620_),
    .Y(_02722_));
 sky130_fd_sc_hd__nand2_1 _26573_ (.A(_02721_),
    .B(_02722_),
    .Y(_02723_));
 sky130_fd_sc_hd__or2_1 _26574_ (.A(_02657_),
    .B(_02723_),
    .X(_02725_));
 sky130_fd_sc_hd__nand2_1 _26575_ (.A(_02723_),
    .B(_02657_),
    .Y(_02726_));
 sky130_fd_sc_hd__nand2_1 _26576_ (.A(_02725_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__or3_1 _26577_ (.A(_02364_),
    .B(_02656_),
    .C(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__o21ai_1 _26578_ (.A1(_02421_),
    .A2(_02656_),
    .B1(_02727_),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_1 _26579_ (.A(_02728_),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__or2_1 _26580_ (.A(_02625_),
    .B(_02730_),
    .X(_02731_));
 sky130_fd_sc_hd__nand2_1 _26581_ (.A(_02730_),
    .B(_02625_),
    .Y(_02732_));
 sky130_fd_sc_hd__nand2_1 _26582_ (.A(_02731_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__or2_1 _26583_ (.A(_02629_),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__nand2_1 _26584_ (.A(_02733_),
    .B(_02629_),
    .Y(_02736_));
 sky130_fd_sc_hd__nand2_1 _26585_ (.A(_02734_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__or2_1 _26586_ (.A(_02632_),
    .B(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__nand2_1 _26587_ (.A(_02737_),
    .B(_02632_),
    .Y(_02739_));
 sky130_fd_sc_hd__nand2_1 _26588_ (.A(_02738_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__or2_1 _26589_ (.A(_02635_),
    .B(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__nand2_1 _26590_ (.A(_02740_),
    .B(_02635_),
    .Y(_02742_));
 sky130_fd_sc_hd__nand2_1 _26591_ (.A(_02741_),
    .B(_02742_),
    .Y(_02743_));
 sky130_fd_sc_hd__or2_1 _26592_ (.A(_02639_),
    .B(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__nand2_1 _26593_ (.A(_02743_),
    .B(_02639_),
    .Y(_02745_));
 sky130_fd_sc_hd__nand2_1 _26594_ (.A(_02744_),
    .B(_02745_),
    .Y(_02747_));
 sky130_fd_sc_hd__or2_1 _26595_ (.A(_02642_),
    .B(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__nand2_1 _26596_ (.A(_02747_),
    .B(_02642_),
    .Y(_02749_));
 sky130_fd_sc_hd__nand2_1 _26597_ (.A(_02748_),
    .B(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__or2_1 _26598_ (.A(_02645_),
    .B(_02750_),
    .X(_02751_));
 sky130_fd_sc_hd__nand2_1 _26599_ (.A(_02750_),
    .B(_02645_),
    .Y(_02752_));
 sky130_fd_sc_hd__nand2_1 _26600_ (.A(_02751_),
    .B(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__or2_1 _26601_ (.A(_02649_),
    .B(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__nand2_1 _26602_ (.A(_02753_),
    .B(_02649_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_1 _26603_ (.A(_02754_),
    .B(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__a21o_1 _26604_ (.A1(_02756_),
    .A2(_02653_),
    .B1(_02655_),
    .X(_00019_));
 sky130_fd_sc_hd__nor2_1 _26605_ (.A(_02600_),
    .B(_02699_),
    .Y(_02758_));
 sky130_fd_sc_hd__and3_1 _26606_ (.A(_02676_),
    .B(_02580_),
    .C(_02677_),
    .X(_02759_));
 sky130_fd_sc_hd__inv_2 _26607_ (.A(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__nand2_1 _26608_ (.A(net18),
    .B(net17),
    .Y(_02761_));
 sky130_fd_sc_hd__or2_1 _26609_ (.A(_02569_),
    .B(_02761_),
    .X(_02762_));
 sky130_fd_sc_hd__a31o_1 _26610_ (.A1(_08790_),
    .A2(net16),
    .A3(net17),
    .B1(net18),
    .X(_02763_));
 sky130_fd_sc_hd__o21ai_1 _26611_ (.A1(_07088_),
    .A2(_02762_),
    .B1(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__or2_1 _26612_ (.A(net50),
    .B(_02764_),
    .X(_02765_));
 sky130_fd_sc_hd__nand2_1 _26613_ (.A(_02764_),
    .B(net50),
    .Y(_02766_));
 sky130_fd_sc_hd__nand2_1 _26614_ (.A(_02765_),
    .B(_02766_),
    .Y(_02768_));
 sky130_fd_sc_hd__or2_1 _26615_ (.A(_02666_),
    .B(_02768_),
    .X(_02769_));
 sky130_fd_sc_hd__nand2_1 _26616_ (.A(_02768_),
    .B(_02666_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _26617_ (.A(_02769_),
    .B(_02770_),
    .Y(_02771_));
 sky130_fd_sc_hd__or2_1 _26618_ (.A(_02670_),
    .B(_02771_),
    .X(_02772_));
 sky130_fd_sc_hd__nand2_1 _26619_ (.A(_02771_),
    .B(_02670_),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_2 _26620_ (.A(_02772_),
    .B(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hd__and2_1 _26621_ (.A(_02774_),
    .B(_02672_),
    .X(_02775_));
 sky130_fd_sc_hd__nand2_1 _26622_ (.A(_02775_),
    .B(_02578_),
    .Y(_02776_));
 sky130_fd_sc_hd__or2b_1 _26623_ (.A(_02774_),
    .B_N(_02677_),
    .X(_02777_));
 sky130_fd_sc_hd__nand2_1 _26624_ (.A(_02776_),
    .B(_02777_),
    .Y(_02779_));
 sky130_fd_sc_hd__or3_1 _26625_ (.A(_02138_),
    .B(_02760_),
    .C(_02779_),
    .X(_02780_));
 sky130_fd_sc_hd__o21ai_1 _26626_ (.A1(_02138_),
    .A2(_02760_),
    .B1(_02779_),
    .Y(_02781_));
 sky130_fd_sc_hd__nand2_1 _26627_ (.A(_02780_),
    .B(_02781_),
    .Y(_02782_));
 sky130_fd_sc_hd__or2_1 _26628_ (.A(_02681_),
    .B(_02782_),
    .X(_02783_));
 sky130_fd_sc_hd__nand2_1 _26629_ (.A(_02782_),
    .B(_02681_),
    .Y(_02784_));
 sky130_fd_sc_hd__nand2_1 _26630_ (.A(_02783_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__inv_2 _26631_ (.A(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__or2_1 _26632_ (.A(_02684_),
    .B(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__nand2_1 _26633_ (.A(_02786_),
    .B(_02684_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _26634_ (.A(_02787_),
    .B(_02788_),
    .Y(_02790_));
 sky130_fd_sc_hd__inv_2 _26635_ (.A(_02790_),
    .Y(_02791_));
 sky130_fd_sc_hd__or2_1 _26636_ (.A(_02687_),
    .B(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__nand2_1 _26637_ (.A(_02791_),
    .B(_02687_),
    .Y(_02793_));
 sky130_fd_sc_hd__nand2_1 _26638_ (.A(_02792_),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hd__inv_2 _26639_ (.A(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__inv_2 _26640_ (.A(_02690_),
    .Y(_02796_));
 sky130_fd_sc_hd__nand2_1 _26641_ (.A(_02795_),
    .B(_02796_),
    .Y(_02797_));
 sky130_fd_sc_hd__nand2_1 _26642_ (.A(_02794_),
    .B(_02690_),
    .Y(_02798_));
 sky130_fd_sc_hd__nand2_1 _26643_ (.A(_02797_),
    .B(_02798_),
    .Y(_02799_));
 sky130_fd_sc_hd__or2_1 _26644_ (.A(_02694_),
    .B(_02799_),
    .X(_02801_));
 sky130_fd_sc_hd__nand2_1 _26645_ (.A(_02799_),
    .B(_02694_),
    .Y(_02802_));
 sky130_fd_sc_hd__nand2_1 _26646_ (.A(_02801_),
    .B(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__inv_2 _26647_ (.A(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__inv_2 _26648_ (.A(_02698_),
    .Y(_02805_));
 sky130_fd_sc_hd__nand2_1 _26649_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__nand2_1 _26650_ (.A(_02803_),
    .B(_02698_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand2_1 _26651_ (.A(_02806_),
    .B(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__inv_2 _26652_ (.A(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__or2_1 _26653_ (.A(_02758_),
    .B(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__nand2_1 _26654_ (.A(_02809_),
    .B(_02758_),
    .Y(_02812_));
 sky130_fd_sc_hd__nand2_1 _26655_ (.A(_02810_),
    .B(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hd__inv_2 _26656_ (.A(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__or2_1 _26657_ (.A(_02703_),
    .B(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__nand2_1 _26658_ (.A(_02814_),
    .B(_02703_),
    .Y(_02816_));
 sky130_fd_sc_hd__nand2_1 _26659_ (.A(_02815_),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__or2_1 _26660_ (.A(_02706_),
    .B(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__nand2_1 _26661_ (.A(_02817_),
    .B(_02706_),
    .Y(_02819_));
 sky130_fd_sc_hd__nand2_1 _26662_ (.A(_02818_),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__or2_1 _26663_ (.A(_02709_),
    .B(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__nand2_1 _26664_ (.A(_02820_),
    .B(_02709_),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _26665_ (.A(_02821_),
    .B(_02823_),
    .Y(_02824_));
 sky130_fd_sc_hd__or2_1 _26666_ (.A(_02715_),
    .B(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__nand2_1 _26667_ (.A(_02824_),
    .B(_02715_),
    .Y(_02826_));
 sky130_fd_sc_hd__nand2_1 _26668_ (.A(_02825_),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__or2_1 _26669_ (.A(_02718_),
    .B(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__nand2_1 _26670_ (.A(_02827_),
    .B(_02718_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2_1 _26671_ (.A(_02828_),
    .B(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__or2_1 _26672_ (.A(_02721_),
    .B(_02830_),
    .X(_02831_));
 sky130_fd_sc_hd__nand2_1 _26673_ (.A(_02830_),
    .B(_02721_),
    .Y(_02832_));
 sky130_fd_sc_hd__nand2_1 _26674_ (.A(_02831_),
    .B(_02832_),
    .Y(_02834_));
 sky130_fd_sc_hd__or2_1 _26675_ (.A(_02725_),
    .B(_02834_),
    .X(_02835_));
 sky130_fd_sc_hd__nand2_1 _26676_ (.A(_02834_),
    .B(_02725_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand2_1 _26677_ (.A(_02835_),
    .B(_02836_),
    .Y(_02837_));
 sky130_fd_sc_hd__or2_1 _26678_ (.A(_02728_),
    .B(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__nand2_1 _26679_ (.A(_02837_),
    .B(_02728_),
    .Y(_02839_));
 sky130_fd_sc_hd__nand2_1 _26680_ (.A(_02838_),
    .B(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__or2_1 _26681_ (.A(_02731_),
    .B(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__nand2_1 _26682_ (.A(_02840_),
    .B(_02731_),
    .Y(_02842_));
 sky130_fd_sc_hd__nand2_1 _26683_ (.A(_02841_),
    .B(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__or2_1 _26684_ (.A(_02734_),
    .B(_02843_),
    .X(_02845_));
 sky130_fd_sc_hd__nand2_1 _26685_ (.A(_02843_),
    .B(_02734_),
    .Y(_02846_));
 sky130_fd_sc_hd__nand2_1 _26686_ (.A(_02845_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__or2_1 _26687_ (.A(_02738_),
    .B(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__nand2_1 _26688_ (.A(_02847_),
    .B(_02738_),
    .Y(_02849_));
 sky130_fd_sc_hd__nand2_1 _26689_ (.A(_02848_),
    .B(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__or2_1 _26690_ (.A(_02741_),
    .B(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__nand2_1 _26691_ (.A(_02850_),
    .B(_02741_),
    .Y(_02852_));
 sky130_fd_sc_hd__nand2_1 _26692_ (.A(_02851_),
    .B(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__or2_1 _26693_ (.A(_02744_),
    .B(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__nand2_1 _26694_ (.A(_02853_),
    .B(_02744_),
    .Y(_02856_));
 sky130_fd_sc_hd__nand2_1 _26695_ (.A(_02854_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__or2_1 _26696_ (.A(_02748_),
    .B(_02857_),
    .X(_02858_));
 sky130_fd_sc_hd__nand2_1 _26697_ (.A(_02857_),
    .B(_02748_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_1 _26698_ (.A(_02858_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__or2_1 _26699_ (.A(_02751_),
    .B(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__nand2_1 _26700_ (.A(_02860_),
    .B(_02751_),
    .Y(_02862_));
 sky130_fd_sc_hd__nand2_1 _26701_ (.A(_02861_),
    .B(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__or2_1 _26702_ (.A(_02754_),
    .B(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__nand2_1 _26703_ (.A(_02863_),
    .B(_02754_),
    .Y(_02865_));
 sky130_fd_sc_hd__and2_1 _26704_ (.A(_02864_),
    .B(_02865_),
    .X(_02867_));
 sky130_fd_sc_hd__o21ai_1 _26705_ (.A1(_02134_),
    .A2(_02867_),
    .B1(net154),
    .Y(_00020_));
 sky130_fd_sc_hd__inv_2 _26706_ (.A(_02816_),
    .Y(_02868_));
 sky130_fd_sc_hd__inv_2 _26707_ (.A(_02806_),
    .Y(_02869_));
 sky130_fd_sc_hd__nor2_1 _26708_ (.A(_02762_),
    .B(_07088_),
    .Y(_02870_));
 sky130_fd_sc_hd__or2_1 _26709_ (.A(net19),
    .B(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__nand2_1 _26710_ (.A(_02870_),
    .B(net19),
    .Y(_02872_));
 sky130_fd_sc_hd__nand2_1 _26711_ (.A(_02871_),
    .B(_02872_),
    .Y(_02873_));
 sky130_fd_sc_hd__or2_1 _26712_ (.A(net51),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__nand2_1 _26713_ (.A(_02873_),
    .B(net51),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _26714_ (.A(_02874_),
    .B(_02875_),
    .Y(_02877_));
 sky130_fd_sc_hd__or2_1 _26715_ (.A(_02765_),
    .B(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__nand2_1 _26716_ (.A(_02877_),
    .B(_02765_),
    .Y(_02879_));
 sky130_fd_sc_hd__nand2_1 _26717_ (.A(_02878_),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__inv_2 _26718_ (.A(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__nand2_1 _26719_ (.A(_02772_),
    .B(_02769_),
    .Y(_02882_));
 sky130_fd_sc_hd__or2_1 _26720_ (.A(_02881_),
    .B(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__nand2_1 _26721_ (.A(_02882_),
    .B(_02881_),
    .Y(_02884_));
 sky130_fd_sc_hd__nand2_4 _26722_ (.A(_02883_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__xor2_1 _26723_ (.A(_02776_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__or2_1 _26724_ (.A(_02886_),
    .B(_02780_),
    .X(_02888_));
 sky130_fd_sc_hd__nand2_1 _26725_ (.A(_02780_),
    .B(_02886_),
    .Y(_02889_));
 sky130_fd_sc_hd__nand2_1 _26726_ (.A(_02888_),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__or2_1 _26727_ (.A(_02783_),
    .B(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__nand2_1 _26728_ (.A(_02783_),
    .B(_02890_),
    .Y(_02892_));
 sky130_fd_sc_hd__nand2_1 _26729_ (.A(_02891_),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__or2_1 _26730_ (.A(_02788_),
    .B(_02893_),
    .X(_02894_));
 sky130_fd_sc_hd__nand2_1 _26731_ (.A(_02893_),
    .B(_02788_),
    .Y(_02895_));
 sky130_fd_sc_hd__nand2_1 _26732_ (.A(_02894_),
    .B(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__or2_1 _26733_ (.A(_02793_),
    .B(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__nand2_1 _26734_ (.A(_02896_),
    .B(_02793_),
    .Y(_02899_));
 sky130_fd_sc_hd__and2_1 _26735_ (.A(_02897_),
    .B(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__inv_2 _26736_ (.A(_02797_),
    .Y(_02901_));
 sky130_fd_sc_hd__or2_1 _26737_ (.A(_02900_),
    .B(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__nand2_1 _26738_ (.A(_02901_),
    .B(_02900_),
    .Y(_02903_));
 sky130_fd_sc_hd__nand2_1 _26739_ (.A(_02902_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__nor2_1 _26740_ (.A(_02801_),
    .B(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__and2_1 _26741_ (.A(_02904_),
    .B(_02801_),
    .X(_02906_));
 sky130_fd_sc_hd__nor2_1 _26742_ (.A(_02905_),
    .B(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hd__or2_1 _26743_ (.A(_02869_),
    .B(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__nand2_1 _26744_ (.A(_02907_),
    .B(_02869_),
    .Y(_02910_));
 sky130_fd_sc_hd__nand2_1 _26745_ (.A(_02908_),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__nor2_1 _26746_ (.A(_02812_),
    .B(_02911_),
    .Y(_02912_));
 sky130_fd_sc_hd__and2_1 _26747_ (.A(_02911_),
    .B(_02812_),
    .X(_02913_));
 sky130_fd_sc_hd__nor2_1 _26748_ (.A(_02912_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__or2_1 _26749_ (.A(_02868_),
    .B(_02914_),
    .X(_02915_));
 sky130_fd_sc_hd__nand2_1 _26750_ (.A(_02914_),
    .B(_02868_),
    .Y(_02916_));
 sky130_fd_sc_hd__nand2_2 _26751_ (.A(_02915_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__a21bo_1 _26752_ (.A1(_02708_),
    .A2(_02819_),
    .B1_N(_02818_),
    .X(_02918_));
 sky130_fd_sc_hd__xnor2_1 _26753_ (.A(_02917_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__or2b_1 _26754_ (.A(_02919_),
    .B_N(_02825_),
    .X(_02921_));
 sky130_fd_sc_hd__or2b_1 _26755_ (.A(_02825_),
    .B_N(_02919_),
    .X(_02922_));
 sky130_fd_sc_hd__nand2_1 _26756_ (.A(_02921_),
    .B(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__nor2_1 _26757_ (.A(_02828_),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_1 _26758_ (.A(_02923_),
    .B(_02828_),
    .Y(_02925_));
 sky130_fd_sc_hd__or2b_1 _26759_ (.A(_02924_),
    .B_N(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__nor2_1 _26760_ (.A(_02831_),
    .B(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__inv_2 _26761_ (.A(_02927_),
    .Y(_02928_));
 sky130_fd_sc_hd__nand2_1 _26762_ (.A(_02926_),
    .B(_02831_),
    .Y(_02929_));
 sky130_fd_sc_hd__nand2_1 _26763_ (.A(_02928_),
    .B(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hd__or2_1 _26764_ (.A(_02930_),
    .B(_02835_),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_1 _26765_ (.A(_02835_),
    .B(_02930_),
    .Y(_02933_));
 sky130_fd_sc_hd__nand2_1 _26766_ (.A(_02932_),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__or2_1 _26767_ (.A(_02838_),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__nand2_1 _26768_ (.A(_02934_),
    .B(_02838_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand2_1 _26769_ (.A(_02935_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hd__or2_1 _26770_ (.A(_02841_),
    .B(_02937_),
    .X(_02938_));
 sky130_fd_sc_hd__nand2_1 _26771_ (.A(_02937_),
    .B(_02841_),
    .Y(_02939_));
 sky130_fd_sc_hd__nand2_1 _26772_ (.A(_02938_),
    .B(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__or2_1 _26773_ (.A(_02845_),
    .B(_02940_),
    .X(_02941_));
 sky130_fd_sc_hd__nand2_1 _26774_ (.A(_02940_),
    .B(_02845_),
    .Y(_02943_));
 sky130_fd_sc_hd__nand2_1 _26775_ (.A(_02941_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__or2_1 _26776_ (.A(_02848_),
    .B(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__nand2_1 _26777_ (.A(_02944_),
    .B(_02848_),
    .Y(_02946_));
 sky130_fd_sc_hd__nand2_1 _26778_ (.A(_02945_),
    .B(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__or2_1 _26779_ (.A(_02851_),
    .B(_02947_),
    .X(_02948_));
 sky130_fd_sc_hd__nand2_1 _26780_ (.A(_02947_),
    .B(_02851_),
    .Y(_02949_));
 sky130_fd_sc_hd__nand2_1 _26781_ (.A(_02948_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__or2_1 _26782_ (.A(_02854_),
    .B(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__nand2_1 _26783_ (.A(_02950_),
    .B(_02854_),
    .Y(_02952_));
 sky130_fd_sc_hd__nand2_1 _26784_ (.A(_02951_),
    .B(_02952_),
    .Y(_02954_));
 sky130_fd_sc_hd__or2_1 _26785_ (.A(_02858_),
    .B(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__nand2_1 _26786_ (.A(_02954_),
    .B(_02858_),
    .Y(_02956_));
 sky130_fd_sc_hd__nand2_1 _26787_ (.A(_02955_),
    .B(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__or2_1 _26788_ (.A(_02861_),
    .B(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__nand2_1 _26789_ (.A(_02957_),
    .B(_02861_),
    .Y(_02959_));
 sky130_fd_sc_hd__nand2_1 _26790_ (.A(_02958_),
    .B(_02959_),
    .Y(_02960_));
 sky130_fd_sc_hd__or4_1 _26791_ (.A(_02647_),
    .B(_02753_),
    .C(_02863_),
    .D(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__nor2_1 _26792_ (.A(_02568_),
    .B(_02961_),
    .Y(_02962_));
 sky130_fd_sc_hd__inv_2 _26793_ (.A(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__nand2_1 _26794_ (.A(_02960_),
    .B(_02864_),
    .Y(_02965_));
 sky130_fd_sc_hd__nand2_1 _26795_ (.A(_02963_),
    .B(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__a21o_1 _26796_ (.A1(_02966_),
    .A2(_02653_),
    .B1(_02655_),
    .X(_00021_));
 sky130_fd_sc_hd__or4_1 _26797_ (.A(_02644_),
    .B(_02750_),
    .C(_02860_),
    .D(_02957_),
    .X(_02967_));
 sky130_fd_sc_hd__or4_1 _26798_ (.A(_02433_),
    .B(_02628_),
    .C(_02733_),
    .D(_02843_),
    .X(_02968_));
 sky130_fd_sc_hd__or3_1 _26799_ (.A(_02624_),
    .B(_02730_),
    .C(_02840_),
    .X(_02969_));
 sky130_fd_sc_hd__nor2_1 _26800_ (.A(_02917_),
    .B(_02821_),
    .Y(_02970_));
 sky130_fd_sc_hd__nor2_1 _26801_ (.A(_02917_),
    .B(_02818_),
    .Y(_02971_));
 sky130_fd_sc_hd__nand2_1 _26802_ (.A(_02885_),
    .B(_02775_),
    .Y(_02972_));
 sky130_fd_sc_hd__nor3_1 _26803_ (.A(_02184_),
    .B(_02576_),
    .C(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hd__inv_2 _26804_ (.A(net20),
    .Y(_02975_));
 sky130_fd_sc_hd__or2_1 _26805_ (.A(_02975_),
    .B(_02872_),
    .X(_02976_));
 sky130_fd_sc_hd__nand2_1 _26806_ (.A(_02872_),
    .B(_02975_),
    .Y(_02977_));
 sky130_fd_sc_hd__nand2_1 _26807_ (.A(_02976_),
    .B(_02977_),
    .Y(_02978_));
 sky130_fd_sc_hd__or2_1 _26808_ (.A(net52),
    .B(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__nand2_1 _26809_ (.A(_02978_),
    .B(net52),
    .Y(_02980_));
 sky130_fd_sc_hd__nand2_1 _26810_ (.A(_02979_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__or2_1 _26811_ (.A(_02874_),
    .B(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__nand2_1 _26812_ (.A(_02981_),
    .B(_02874_),
    .Y(_02983_));
 sky130_fd_sc_hd__nand2_1 _26813_ (.A(_02982_),
    .B(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__inv_2 _26814_ (.A(_02984_),
    .Y(_02986_));
 sky130_fd_sc_hd__nand2_1 _26815_ (.A(_02884_),
    .B(_02878_),
    .Y(_02987_));
 sky130_fd_sc_hd__or2_1 _26816_ (.A(_02986_),
    .B(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__nand2_1 _26817_ (.A(_02987_),
    .B(_02986_),
    .Y(_02989_));
 sky130_fd_sc_hd__nand2_4 _26818_ (.A(_02988_),
    .B(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__inv_2 _26819_ (.A(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__or2_1 _26820_ (.A(_02577_),
    .B(_02972_),
    .X(_02992_));
 sky130_fd_sc_hd__nor2_1 _26821_ (.A(_02991_),
    .B(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__and2_1 _26822_ (.A(_02992_),
    .B(_02991_),
    .X(_02994_));
 sky130_fd_sc_hd__nor2_1 _26823_ (.A(_02993_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__or2_1 _26824_ (.A(_02973_),
    .B(_02995_),
    .X(_02997_));
 sky130_fd_sc_hd__nand2_1 _26825_ (.A(_02995_),
    .B(_02973_),
    .Y(_02998_));
 sky130_fd_sc_hd__nand2_1 _26826_ (.A(_02997_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__or2_1 _26827_ (.A(_02888_),
    .B(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__nand2_1 _26828_ (.A(_02999_),
    .B(_02888_),
    .Y(_03001_));
 sky130_fd_sc_hd__nand2_1 _26829_ (.A(_03000_),
    .B(_03001_),
    .Y(_03002_));
 sky130_fd_sc_hd__or2_1 _26830_ (.A(_02891_),
    .B(_03002_),
    .X(_03003_));
 sky130_fd_sc_hd__nand2_1 _26831_ (.A(_03002_),
    .B(_02891_),
    .Y(_03004_));
 sky130_fd_sc_hd__nand2_1 _26832_ (.A(_03003_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__or2_1 _26833_ (.A(_02894_),
    .B(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__nand2_1 _26834_ (.A(_03005_),
    .B(_02894_),
    .Y(_03008_));
 sky130_fd_sc_hd__nand2_1 _26835_ (.A(_03006_),
    .B(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__or2_1 _26836_ (.A(_02897_),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__nand2_1 _26837_ (.A(_03009_),
    .B(_02897_),
    .Y(_03011_));
 sky130_fd_sc_hd__nand2_1 _26838_ (.A(_03010_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__or2_1 _26839_ (.A(_02903_),
    .B(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__nand2_1 _26840_ (.A(_03012_),
    .B(_02903_),
    .Y(_03014_));
 sky130_fd_sc_hd__nand2_1 _26841_ (.A(_03013_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__inv_2 _26842_ (.A(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__or2_1 _26843_ (.A(_02905_),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__nand2_1 _26844_ (.A(_03016_),
    .B(_02905_),
    .Y(_03019_));
 sky130_fd_sc_hd__nand2_1 _26845_ (.A(_03017_),
    .B(_03019_),
    .Y(_03020_));
 sky130_fd_sc_hd__or2_1 _26846_ (.A(_02910_),
    .B(_03020_),
    .X(_03021_));
 sky130_fd_sc_hd__nand2_1 _26847_ (.A(_03020_),
    .B(_02910_),
    .Y(_03022_));
 sky130_fd_sc_hd__nand2_1 _26848_ (.A(_03021_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__inv_2 _26849_ (.A(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__or2_1 _26850_ (.A(_02912_),
    .B(_03024_),
    .X(_03025_));
 sky130_fd_sc_hd__nand2_1 _26851_ (.A(_03024_),
    .B(_02912_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand2_1 _26852_ (.A(_03025_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__or2_1 _26853_ (.A(_02916_),
    .B(_03027_),
    .X(_03028_));
 sky130_fd_sc_hd__nand2_1 _26854_ (.A(_03027_),
    .B(_02916_),
    .Y(_03030_));
 sky130_fd_sc_hd__nand2_1 _26855_ (.A(_03028_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__inv_2 _26856_ (.A(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__or2_1 _26857_ (.A(_02971_),
    .B(_03032_),
    .X(_03033_));
 sky130_fd_sc_hd__nand2_1 _26858_ (.A(_03032_),
    .B(_02971_),
    .Y(_03034_));
 sky130_fd_sc_hd__nand2_1 _26859_ (.A(_03033_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__inv_2 _26860_ (.A(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__or2_1 _26861_ (.A(_02970_),
    .B(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__nand2_1 _26862_ (.A(_03036_),
    .B(_02970_),
    .Y(_03038_));
 sky130_fd_sc_hd__nand2_1 _26863_ (.A(_03037_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hd__or4b_1 _26864_ (.A(_02612_),
    .B(_02711_),
    .C(_02824_),
    .D_N(_02919_),
    .X(_03041_));
 sky130_fd_sc_hd__or3_1 _26865_ (.A(_02344_),
    .B(_03039_),
    .C(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__nand2_1 _26866_ (.A(_03039_),
    .B(_02922_),
    .Y(_03043_));
 sky130_fd_sc_hd__nand2_1 _26867_ (.A(_03042_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__inv_2 _26868_ (.A(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__or2_1 _26869_ (.A(_02924_),
    .B(_03045_),
    .X(_03046_));
 sky130_fd_sc_hd__nand2_1 _26870_ (.A(_03045_),
    .B(_02924_),
    .Y(_03047_));
 sky130_fd_sc_hd__nand2_1 _26871_ (.A(_03046_),
    .B(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__or2_1 _26872_ (.A(_02928_),
    .B(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__nand2_1 _26873_ (.A(_03048_),
    .B(_02928_),
    .Y(_03050_));
 sky130_fd_sc_hd__nand2_1 _26874_ (.A(_03049_),
    .B(_03050_),
    .Y(_03052_));
 sky130_fd_sc_hd__or2_1 _26875_ (.A(_02932_),
    .B(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__nand2_1 _26876_ (.A(_03052_),
    .B(_02932_),
    .Y(_03054_));
 sky130_fd_sc_hd__nand2_1 _26877_ (.A(_03053_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hd__or2_1 _26878_ (.A(_02935_),
    .B(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__nand2_1 _26879_ (.A(_03055_),
    .B(_02935_),
    .Y(_03057_));
 sky130_fd_sc_hd__nand2_1 _26880_ (.A(_03056_),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__or4_1 _26881_ (.A(_02367_),
    .B(_02937_),
    .C(_02969_),
    .D(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__nand2_1 _26882_ (.A(_03058_),
    .B(_02938_),
    .Y(_03060_));
 sky130_fd_sc_hd__nand2_1 _26883_ (.A(_03059_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__or3_1 _26884_ (.A(_02968_),
    .B(_02940_),
    .C(_03061_),
    .X(_03063_));
 sky130_fd_sc_hd__nand2_1 _26885_ (.A(_03061_),
    .B(_02941_),
    .Y(_03064_));
 sky130_fd_sc_hd__nand2_1 _26886_ (.A(_03063_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__or2_1 _26887_ (.A(_02945_),
    .B(_03065_),
    .X(_03066_));
 sky130_fd_sc_hd__nand2_1 _26888_ (.A(_03065_),
    .B(_02945_),
    .Y(_03067_));
 sky130_fd_sc_hd__nand2_1 _26889_ (.A(_03066_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__or2_1 _26890_ (.A(_02948_),
    .B(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__nand2_1 _26891_ (.A(_03068_),
    .B(_02948_),
    .Y(_03070_));
 sky130_fd_sc_hd__nand2_1 _26892_ (.A(_03069_),
    .B(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__or2_1 _26893_ (.A(_02951_),
    .B(_03071_),
    .X(_03072_));
 sky130_fd_sc_hd__nand2_1 _26894_ (.A(_03071_),
    .B(_02951_),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2_1 _26895_ (.A(_03072_),
    .B(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hd__or2_1 _26896_ (.A(_02955_),
    .B(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__nand2_1 _26897_ (.A(_03075_),
    .B(_02955_),
    .Y(_03077_));
 sky130_fd_sc_hd__nand2_1 _26898_ (.A(_03076_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hd__or3_1 _26899_ (.A(_02566_),
    .B(_02967_),
    .C(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__nand2_1 _26900_ (.A(_03078_),
    .B(_02958_),
    .Y(_03080_));
 sky130_fd_sc_hd__nand2_1 _26901_ (.A(_03079_),
    .B(_03080_),
    .Y(_03081_));
 sky130_fd_sc_hd__inv_2 _26902_ (.A(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__nor2_1 _26903_ (.A(_02864_),
    .B(_02960_),
    .Y(_03083_));
 sky130_fd_sc_hd__nand2_2 _26904_ (.A(_03082_),
    .B(_03083_),
    .Y(_03085_));
 sky130_fd_sc_hd__nand2_1 _26905_ (.A(_03081_),
    .B(_02963_),
    .Y(_03086_));
 sky130_fd_sc_hd__nand2_1 _26906_ (.A(_03085_),
    .B(_03086_),
    .Y(_03087_));
 sky130_fd_sc_hd__a21o_1 _26907_ (.A1(_03087_),
    .A2(_02653_),
    .B1(_02655_),
    .X(_00022_));
 sky130_fd_sc_hd__inv_2 _26908_ (.A(_03028_),
    .Y(_03088_));
 sky130_fd_sc_hd__inv_2 _26909_ (.A(_03021_),
    .Y(_03089_));
 sky130_fd_sc_hd__inv_2 _26910_ (.A(net21),
    .Y(_03090_));
 sky130_fd_sc_hd__nor2_1 _26911_ (.A(_03090_),
    .B(_02976_),
    .Y(_03091_));
 sky130_fd_sc_hd__nand2_1 _26912_ (.A(_02976_),
    .B(_03090_),
    .Y(_03092_));
 sky130_fd_sc_hd__or2b_1 _26913_ (.A(_03091_),
    .B_N(_03092_),
    .X(_03093_));
 sky130_fd_sc_hd__or2_1 _26914_ (.A(net53),
    .B(_03093_),
    .X(_03095_));
 sky130_fd_sc_hd__nand2_1 _26915_ (.A(_03093_),
    .B(net53),
    .Y(_03096_));
 sky130_fd_sc_hd__nand2_1 _26916_ (.A(_03095_),
    .B(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__or2_1 _26917_ (.A(_02979_),
    .B(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__nand2_1 _26918_ (.A(_03097_),
    .B(_02979_),
    .Y(_03099_));
 sky130_fd_sc_hd__nand2_1 _26919_ (.A(_03098_),
    .B(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__inv_2 _26920_ (.A(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_1 _26921_ (.A(_02989_),
    .B(_02982_),
    .Y(_03102_));
 sky130_fd_sc_hd__or2_1 _26922_ (.A(_03101_),
    .B(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__nand2_1 _26923_ (.A(_03102_),
    .B(_03101_),
    .Y(_03104_));
 sky130_fd_sc_hd__nand2_4 _26924_ (.A(_03103_),
    .B(_03104_),
    .Y(_03106_));
 sky130_fd_sc_hd__or2_1 _26925_ (.A(_03106_),
    .B(_02993_),
    .X(_03107_));
 sky130_fd_sc_hd__nand2_1 _26926_ (.A(_02993_),
    .B(_03106_),
    .Y(_03108_));
 sky130_fd_sc_hd__a22o_1 _26927_ (.A1(_02995_),
    .A2(_02973_),
    .B1(_03107_),
    .B2(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__or2b_1 _26928_ (.A(_02998_),
    .B_N(_03106_),
    .X(_03110_));
 sky130_fd_sc_hd__nand2_1 _26929_ (.A(_03109_),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__or2_1 _26930_ (.A(_03111_),
    .B(_03000_),
    .X(_03112_));
 sky130_fd_sc_hd__nand2_1 _26931_ (.A(_03000_),
    .B(_03111_),
    .Y(_03113_));
 sky130_fd_sc_hd__nand2_1 _26932_ (.A(_03112_),
    .B(_03113_),
    .Y(_03114_));
 sky130_fd_sc_hd__or2_1 _26933_ (.A(_03114_),
    .B(_03006_),
    .X(_03115_));
 sky130_fd_sc_hd__or2_1 _26934_ (.A(_03003_),
    .B(_03114_),
    .X(_03117_));
 sky130_fd_sc_hd__nand2_1 _26935_ (.A(_03114_),
    .B(_03003_),
    .Y(_03118_));
 sky130_fd_sc_hd__nand2_1 _26936_ (.A(_03117_),
    .B(_03118_),
    .Y(_03119_));
 sky130_fd_sc_hd__nand2_1 _26937_ (.A(_03119_),
    .B(_03006_),
    .Y(_03120_));
 sky130_fd_sc_hd__nand2_1 _26938_ (.A(_03115_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__or2_1 _26939_ (.A(_03121_),
    .B(_03013_),
    .X(_03122_));
 sky130_fd_sc_hd__nand2_1 _26940_ (.A(_03013_),
    .B(_03121_),
    .Y(_03123_));
 sky130_fd_sc_hd__nand2_1 _26941_ (.A(_03122_),
    .B(_03123_),
    .Y(_03124_));
 sky130_fd_sc_hd__xnor2_1 _26942_ (.A(_03010_),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__or2_1 _26943_ (.A(_03019_),
    .B(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__nand2_1 _26944_ (.A(_03125_),
    .B(_03019_),
    .Y(_03128_));
 sky130_fd_sc_hd__and2_1 _26945_ (.A(_03126_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__or2_1 _26946_ (.A(_03089_),
    .B(_03129_),
    .X(_03130_));
 sky130_fd_sc_hd__nand2_1 _26947_ (.A(_03129_),
    .B(_03089_),
    .Y(_03131_));
 sky130_fd_sc_hd__nand2_1 _26948_ (.A(_03130_),
    .B(_03131_),
    .Y(_03132_));
 sky130_fd_sc_hd__or2_1 _26949_ (.A(_03026_),
    .B(_03132_),
    .X(_03133_));
 sky130_fd_sc_hd__nand2_1 _26950_ (.A(_03132_),
    .B(_03026_),
    .Y(_03134_));
 sky130_fd_sc_hd__and2_1 _26951_ (.A(_03133_),
    .B(_03134_),
    .X(_03135_));
 sky130_fd_sc_hd__or2_1 _26952_ (.A(_03088_),
    .B(_03135_),
    .X(_03136_));
 sky130_fd_sc_hd__nand2_1 _26953_ (.A(_03135_),
    .B(_03088_),
    .Y(_03137_));
 sky130_fd_sc_hd__nand2_1 _26954_ (.A(_03136_),
    .B(_03137_),
    .Y(_03139_));
 sky130_fd_sc_hd__or2_1 _26955_ (.A(_03034_),
    .B(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__nand2_1 _26956_ (.A(_03139_),
    .B(_03034_),
    .Y(_03141_));
 sky130_fd_sc_hd__nand2_1 _26957_ (.A(_03140_),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__or2_1 _26958_ (.A(_03038_),
    .B(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__nand2_1 _26959_ (.A(_03142_),
    .B(_03038_),
    .Y(_03144_));
 sky130_fd_sc_hd__nand2_1 _26960_ (.A(_03143_),
    .B(_03144_),
    .Y(_03145_));
 sky130_fd_sc_hd__or2_1 _26961_ (.A(_03145_),
    .B(_03042_),
    .X(_03146_));
 sky130_fd_sc_hd__nand2_1 _26962_ (.A(_03042_),
    .B(_03145_),
    .Y(_03147_));
 sky130_fd_sc_hd__nand2_1 _26963_ (.A(_03146_),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__or2_1 _26964_ (.A(_03047_),
    .B(_03148_),
    .X(_03150_));
 sky130_fd_sc_hd__nand2_1 _26965_ (.A(_03148_),
    .B(_03047_),
    .Y(_03151_));
 sky130_fd_sc_hd__nand2_1 _26966_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__or2_1 _26967_ (.A(_03152_),
    .B(_03049_),
    .X(_03153_));
 sky130_fd_sc_hd__nand2_1 _26968_ (.A(_03049_),
    .B(_03152_),
    .Y(_03154_));
 sky130_fd_sc_hd__nand2_1 _26969_ (.A(_03153_),
    .B(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__or2_1 _26970_ (.A(_03053_),
    .B(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__nand2_1 _26971_ (.A(_03155_),
    .B(_03053_),
    .Y(_03157_));
 sky130_fd_sc_hd__nand2_1 _26972_ (.A(_03156_),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__or2_1 _26973_ (.A(_03056_),
    .B(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__nand2_1 _26974_ (.A(_03158_),
    .B(_03056_),
    .Y(_03161_));
 sky130_fd_sc_hd__nand2_1 _26975_ (.A(_03159_),
    .B(_03161_),
    .Y(_03162_));
 sky130_fd_sc_hd__or2_1 _26976_ (.A(_03162_),
    .B(_03059_),
    .X(_03163_));
 sky130_fd_sc_hd__nand2_1 _26977_ (.A(_03059_),
    .B(_03162_),
    .Y(_03164_));
 sky130_fd_sc_hd__nand2_1 _26978_ (.A(_03163_),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__or2_1 _26979_ (.A(_03165_),
    .B(_03063_),
    .X(_03166_));
 sky130_fd_sc_hd__nand2_1 _26980_ (.A(_03063_),
    .B(_03165_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand2_1 _26981_ (.A(_03166_),
    .B(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__or2_1 _26982_ (.A(_03066_),
    .B(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__nand2_1 _26983_ (.A(_03168_),
    .B(_03066_),
    .Y(_03170_));
 sky130_fd_sc_hd__nand2_1 _26984_ (.A(_03169_),
    .B(_03170_),
    .Y(_03172_));
 sky130_fd_sc_hd__nor2_1 _26985_ (.A(_03069_),
    .B(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__and2_1 _26986_ (.A(_03172_),
    .B(_03069_),
    .X(_03174_));
 sky130_fd_sc_hd__or2_1 _26987_ (.A(_03173_),
    .B(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__and2_1 _26988_ (.A(_03175_),
    .B(_03072_),
    .X(_03176_));
 sky130_fd_sc_hd__or4_1 _26989_ (.A(_02512_),
    .B(_02638_),
    .C(_02743_),
    .D(_02853_),
    .X(_03177_));
 sky130_fd_sc_hd__or3_1 _26990_ (.A(_03177_),
    .B(_02950_),
    .C(_03071_),
    .X(_03178_));
 sky130_fd_sc_hd__nor2_1 _26991_ (.A(_03175_),
    .B(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__or2_1 _26992_ (.A(_03176_),
    .B(_03179_),
    .X(_03180_));
 sky130_fd_sc_hd__or2_1 _26993_ (.A(_03076_),
    .B(_03180_),
    .X(_03181_));
 sky130_fd_sc_hd__nand2_1 _26994_ (.A(_03180_),
    .B(_03076_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2_1 _26995_ (.A(_03181_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__or2_1 _26996_ (.A(_03079_),
    .B(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__nand2_1 _26997_ (.A(_03184_),
    .B(_03079_),
    .Y(_03186_));
 sky130_fd_sc_hd__nand2_1 _26998_ (.A(_03185_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__xor2_2 _26999_ (.A(_03085_),
    .B(_03187_),
    .X(_03188_));
 sky130_fd_sc_hd__o21ai_1 _27000_ (.A1(_02134_),
    .A2(_03188_),
    .B1(net154),
    .Y(_00023_));
 sky130_fd_sc_hd__or3b_1 _27001_ (.A(_02727_),
    .B(_02837_),
    .C_N(_02623_),
    .X(_03189_));
 sky130_fd_sc_hd__or4_1 _27002_ (.A(_02421_),
    .B(_03189_),
    .C(_02934_),
    .D(_03055_),
    .X(_03190_));
 sky130_fd_sc_hd__nor2_1 _27003_ (.A(_03119_),
    .B(_03010_),
    .Y(_03191_));
 sky130_fd_sc_hd__nor2_1 _27004_ (.A(net22),
    .B(_03091_),
    .Y(_03193_));
 sky130_fd_sc_hd__and2_1 _27005_ (.A(_03091_),
    .B(net22),
    .X(_03194_));
 sky130_fd_sc_hd__or2_1 _27006_ (.A(_03193_),
    .B(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__or2_2 _27007_ (.A(net54),
    .B(_03195_),
    .X(_03196_));
 sky130_fd_sc_hd__nand2_1 _27008_ (.A(_03195_),
    .B(net54),
    .Y(_03197_));
 sky130_fd_sc_hd__nand2_1 _27009_ (.A(_03196_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__or2_1 _27010_ (.A(_03095_),
    .B(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__nand2_1 _27011_ (.A(_03198_),
    .B(_03095_),
    .Y(_03200_));
 sky130_fd_sc_hd__and2_1 _27012_ (.A(_03199_),
    .B(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__nand2_1 _27013_ (.A(_03104_),
    .B(_03098_),
    .Y(_03202_));
 sky130_fd_sc_hd__or2_1 _27014_ (.A(_03201_),
    .B(_03202_),
    .X(_03204_));
 sky130_fd_sc_hd__nand2_1 _27015_ (.A(_03202_),
    .B(_03201_),
    .Y(_03205_));
 sky130_fd_sc_hd__nand2_4 _27016_ (.A(_03204_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__inv_2 _27017_ (.A(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__or2_1 _27018_ (.A(_03108_),
    .B(_03207_),
    .X(_03208_));
 sky130_fd_sc_hd__nand2_1 _27019_ (.A(_03207_),
    .B(_03108_),
    .Y(_03209_));
 sky130_fd_sc_hd__nand2_1 _27020_ (.A(_03208_),
    .B(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__or2_1 _27021_ (.A(_03110_),
    .B(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__nand2_1 _27022_ (.A(_03210_),
    .B(_03110_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _27023_ (.A(_03211_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_1 _27024_ (.A(_03213_),
    .B(_03112_),
    .Y(_03215_));
 sky130_fd_sc_hd__xnor2_1 _27025_ (.A(_03117_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__or2_1 _27026_ (.A(_03115_),
    .B(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__nand2_1 _27027_ (.A(_03216_),
    .B(_03115_),
    .Y(_03218_));
 sky130_fd_sc_hd__and2_1 _27028_ (.A(_03217_),
    .B(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__or2_1 _27029_ (.A(_03191_),
    .B(_03219_),
    .X(_03220_));
 sky130_fd_sc_hd__nand2_1 _27030_ (.A(_03219_),
    .B(_03191_),
    .Y(_03221_));
 sky130_fd_sc_hd__nand2_1 _27031_ (.A(_03220_),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__or2_1 _27032_ (.A(_03122_),
    .B(_03222_),
    .X(_03223_));
 sky130_fd_sc_hd__nand2_1 _27033_ (.A(_03222_),
    .B(_03122_),
    .Y(_03224_));
 sky130_fd_sc_hd__nand2_1 _27034_ (.A(_03223_),
    .B(_03224_),
    .Y(_03226_));
 sky130_fd_sc_hd__or2_1 _27035_ (.A(_03226_),
    .B(_03126_),
    .X(_03227_));
 sky130_fd_sc_hd__nand2_1 _27036_ (.A(_03126_),
    .B(_03226_),
    .Y(_03228_));
 sky130_fd_sc_hd__nand2_1 _27037_ (.A(_03227_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__or2_1 _27038_ (.A(_03131_),
    .B(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__nand2_1 _27039_ (.A(_03229_),
    .B(_03131_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _27040_ (.A(_03230_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__or2_1 _27041_ (.A(_03232_),
    .B(_03133_),
    .X(_03233_));
 sky130_fd_sc_hd__nand2_1 _27042_ (.A(_03133_),
    .B(_03232_),
    .Y(_03234_));
 sky130_fd_sc_hd__nand2_1 _27043_ (.A(_03233_),
    .B(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__or2_1 _27044_ (.A(_03137_),
    .B(_03235_),
    .X(_03237_));
 sky130_fd_sc_hd__nand2_1 _27045_ (.A(_03235_),
    .B(_03137_),
    .Y(_03238_));
 sky130_fd_sc_hd__nand2_1 _27046_ (.A(_03237_),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__or2_1 _27047_ (.A(_03239_),
    .B(_03140_),
    .X(_03240_));
 sky130_fd_sc_hd__nand2_1 _27048_ (.A(_03140_),
    .B(_03239_),
    .Y(_03241_));
 sky130_fd_sc_hd__nand2_1 _27049_ (.A(_03240_),
    .B(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__and2_1 _27050_ (.A(_03143_),
    .B(_03242_),
    .X(_03243_));
 sky130_fd_sc_hd__or2_1 _27051_ (.A(_02609_),
    .B(_02707_),
    .X(_03244_));
 sky130_fd_sc_hd__or4_1 _27052_ (.A(_03244_),
    .B(_02820_),
    .C(_02917_),
    .D(_03035_),
    .X(_03245_));
 sky130_fd_sc_hd__or3_1 _27053_ (.A(_02242_),
    .B(_03245_),
    .C(_03142_),
    .X(_03246_));
 sky130_fd_sc_hd__nor2_1 _27054_ (.A(_03242_),
    .B(_03246_),
    .Y(_03248_));
 sky130_fd_sc_hd__or2_1 _27055_ (.A(_03243_),
    .B(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__or4_1 _27056_ (.A(_02922_),
    .B(_03039_),
    .C(_03145_),
    .D(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__nand2_1 _27057_ (.A(_03249_),
    .B(_03146_),
    .Y(_03251_));
 sky130_fd_sc_hd__nand2_1 _27058_ (.A(_03250_),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__or2_1 _27059_ (.A(_03150_),
    .B(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__nand2_1 _27060_ (.A(_03252_),
    .B(_03150_),
    .Y(_03254_));
 sky130_fd_sc_hd__nand2_1 _27061_ (.A(_03253_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__xnor2_1 _27062_ (.A(_03153_),
    .B(_03255_),
    .Y(_03256_));
 sky130_fd_sc_hd__or2_1 _27063_ (.A(_03156_),
    .B(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__nand2_1 _27064_ (.A(_03256_),
    .B(_03156_),
    .Y(_03259_));
 sky130_fd_sc_hd__nand2_1 _27065_ (.A(_03257_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__or3_1 _27066_ (.A(_03190_),
    .B(_03158_),
    .C(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__nand2_1 _27067_ (.A(_03260_),
    .B(_03159_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _27068_ (.A(_03261_),
    .B(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__or2_1 _27069_ (.A(_03163_),
    .B(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__nand2_1 _27070_ (.A(_03263_),
    .B(_03163_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_1 _27071_ (.A(_03264_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__or2_1 _27072_ (.A(_03166_),
    .B(_03266_),
    .X(_03267_));
 sky130_fd_sc_hd__nand2_1 _27073_ (.A(_03266_),
    .B(_03166_),
    .Y(_03268_));
 sky130_fd_sc_hd__nand2_1 _27074_ (.A(_03267_),
    .B(_03268_),
    .Y(_03270_));
 sky130_fd_sc_hd__or2_1 _27075_ (.A(_03169_),
    .B(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__nand2_1 _27076_ (.A(_03270_),
    .B(_03169_),
    .Y(_03272_));
 sky130_fd_sc_hd__a21o_1 _27077_ (.A1(_03271_),
    .A2(_03272_),
    .B1(_03173_),
    .X(_03273_));
 sky130_fd_sc_hd__nand2_1 _27078_ (.A(_03173_),
    .B(_03272_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_1 _27079_ (.A(_03273_),
    .B(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__o21a_1 _27080_ (.A1(_03072_),
    .A2(_03175_),
    .B1(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__or3_1 _27081_ (.A(_03072_),
    .B(_03175_),
    .C(_03275_),
    .X(_03277_));
 sky130_fd_sc_hd__or2b_1 _27082_ (.A(_03276_),
    .B_N(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__xnor2_1 _27083_ (.A(_03181_),
    .B(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__or4_1 _27084_ (.A(_02958_),
    .B(_03078_),
    .C(_03184_),
    .D(_03279_),
    .X(_03281_));
 sky130_fd_sc_hd__nand2_1 _27085_ (.A(_03279_),
    .B(_03185_),
    .Y(_03282_));
 sky130_fd_sc_hd__nor2_1 _27086_ (.A(_03184_),
    .B(_03085_),
    .Y(_03283_));
 sky130_fd_sc_hd__a21o_1 _27087_ (.A1(_03281_),
    .A2(_03282_),
    .B1(_03283_),
    .X(_03284_));
 sky130_fd_sc_hd__nand2_1 _27088_ (.A(_03282_),
    .B(_03283_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _27089_ (.A(_03284_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__a21o_1 _27090_ (.A1(_03286_),
    .A2(_02653_),
    .B1(_02655_),
    .X(_00024_));
 sky130_fd_sc_hd__inv_2 _27091_ (.A(net56),
    .Y(_03287_));
 sky130_fd_sc_hd__inv_2 _27092_ (.A(net24),
    .Y(_03288_));
 sky130_fd_sc_hd__xor2_1 _27093_ (.A(_03288_),
    .B(_03194_),
    .X(_03289_));
 sky130_fd_sc_hd__xor2_2 _27094_ (.A(_03287_),
    .B(_03289_),
    .X(_03291_));
 sky130_fd_sc_hd__xor2_4 _27095_ (.A(_03196_),
    .B(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__nand2_2 _27096_ (.A(_03205_),
    .B(_03199_),
    .Y(_03293_));
 sky130_fd_sc_hd__xor2_4 _27097_ (.A(_03292_),
    .B(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__and2b_1 _27098_ (.A_N(_03294_),
    .B(_03208_),
    .X(_03295_));
 sky130_fd_sc_hd__and2b_4 _27099_ (.A_N(_03208_),
    .B(_03294_),
    .X(_03296_));
 sky130_fd_sc_hd__or2_1 _27100_ (.A(_03295_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__o21ai_1 _27101_ (.A1(_03213_),
    .A2(_03112_),
    .B1(_03211_),
    .Y(_03298_));
 sky130_fd_sc_hd__xor2_1 _27102_ (.A(_03297_),
    .B(_03298_),
    .X(_03299_));
 sky130_fd_sc_hd__o21ai_1 _27103_ (.A1(_03117_),
    .A2(_03215_),
    .B1(_03217_),
    .Y(_03300_));
 sky130_fd_sc_hd__xor2_1 _27104_ (.A(_03299_),
    .B(_03300_),
    .X(_03302_));
 sky130_fd_sc_hd__xnor2_1 _27105_ (.A(_03221_),
    .B(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__nand2_1 _27106_ (.A(_03227_),
    .B(_03223_),
    .Y(_03304_));
 sky130_fd_sc_hd__xor2_1 _27107_ (.A(_03303_),
    .B(_03304_),
    .X(_03305_));
 sky130_fd_sc_hd__nand2_1 _27108_ (.A(_03233_),
    .B(_03230_),
    .Y(_03306_));
 sky130_fd_sc_hd__xnor2_1 _27109_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__xor2_1 _27110_ (.A(_03237_),
    .B(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__xor2_1 _27111_ (.A(_03308_),
    .B(_03240_),
    .X(_03309_));
 sky130_fd_sc_hd__xor2_1 _27112_ (.A(_03309_),
    .B(_03248_),
    .X(_03310_));
 sky130_fd_sc_hd__nand2_1 _27113_ (.A(_03253_),
    .B(_03250_),
    .Y(_03311_));
 sky130_fd_sc_hd__xnor2_1 _27114_ (.A(_03310_),
    .B(_03311_),
    .Y(_03313_));
 sky130_fd_sc_hd__o21ai_1 _27115_ (.A1(_03153_),
    .A2(_03255_),
    .B1(_03257_),
    .Y(_03314_));
 sky130_fd_sc_hd__xor2_1 _27116_ (.A(_03313_),
    .B(_03314_),
    .X(_03315_));
 sky130_fd_sc_hd__xor2_1 _27117_ (.A(_03315_),
    .B(_03261_),
    .X(_03316_));
 sky130_fd_sc_hd__nand2_1 _27118_ (.A(_03267_),
    .B(_03264_),
    .Y(_03317_));
 sky130_fd_sc_hd__xnor2_1 _27119_ (.A(_03316_),
    .B(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__nand2_1 _27120_ (.A(_03274_),
    .B(_03271_),
    .Y(_03319_));
 sky130_fd_sc_hd__xnor2_1 _27121_ (.A(_03318_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__o21ai_1 _27122_ (.A1(_03276_),
    .A2(_03181_),
    .B1(_03277_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_2 _27123_ (.A(_03320_),
    .B(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _27124_ (.A(_03281_),
    .B(_03285_),
    .Y(_03324_));
 sky130_fd_sc_hd__xnor2_2 _27125_ (.A(_03322_),
    .B(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__o21ai_1 _27126_ (.A1(_02134_),
    .A2(_03325_),
    .B1(net154),
    .Y(_00026_));
 sky130_fd_sc_hd__nor2_1 _27127_ (.A(_00161_),
    .B(_01907_),
    .Y(_03326_));
 sky130_fd_sc_hd__or2_1 _27128_ (.A(_11412_),
    .B(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__nand2_1 _27129_ (.A(_03327_),
    .B(_01601_),
    .Y(_03328_));
 sky130_fd_sc_hd__inv_2 _27130_ (.A(_03328_),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _27131_ (.A(_02131_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand3_1 _27132_ (.A(_02128_),
    .B(_02130_),
    .C(_03326_),
    .Y(_03331_));
 sky130_fd_sc_hd__nand2_1 _27133_ (.A(_03330_),
    .B(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand2_2 _27134_ (.A(_03332_),
    .B(_11421_),
    .Y(_03334_));
 sky130_fd_sc_hd__nand3_1 _27135_ (.A(_03330_),
    .B(_11426_),
    .C(_03331_),
    .Y(_03335_));
 sky130_fd_sc_hd__nand3_1 _27136_ (.A(_02131_),
    .B(_00174_),
    .C(_12221_),
    .Y(_03336_));
 sky130_fd_sc_hd__inv_2 _27137_ (.A(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hd__nand3_2 _27138_ (.A(_03334_),
    .B(_03335_),
    .C(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__inv_2 _27139_ (.A(_03338_),
    .Y(_03339_));
 sky130_fd_sc_hd__nand2_1 _27140_ (.A(_01599_),
    .B(_01600_),
    .Y(_03340_));
 sky130_fd_sc_hd__nand2_1 _27141_ (.A(_03340_),
    .B(_01601_),
    .Y(_03341_));
 sky130_fd_sc_hd__nand2_1 _27142_ (.A(_03341_),
    .B(_01603_),
    .Y(_03342_));
 sky130_fd_sc_hd__inv_2 _27143_ (.A(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__nand2_1 _27144_ (.A(net122),
    .B(_03343_),
    .Y(_03345_));
 sky130_fd_sc_hd__o21ai_2 _27145_ (.A1(_00161_),
    .A2(\div1i.quot[1] ),
    .B1(_00174_),
    .Y(_03346_));
 sky130_fd_sc_hd__nand2_1 _27146_ (.A(_03342_),
    .B(_12030_),
    .Y(_03347_));
 sky130_fd_sc_hd__nand3_1 _27147_ (.A(_03341_),
    .B(_12035_),
    .C(_01603_),
    .Y(_03348_));
 sky130_fd_sc_hd__nand2_1 _27148_ (.A(_03347_),
    .B(_03348_),
    .Y(_03349_));
 sky130_fd_sc_hd__xor2_1 _27149_ (.A(_03346_),
    .B(_03349_),
    .X(_03350_));
 sky130_fd_sc_hd__nand3b_1 _27150_ (.A_N(_03350_),
    .B(_02128_),
    .C(_02130_),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _27151_ (.A(_03345_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__nand2_1 _27152_ (.A(_03352_),
    .B(_13679_),
    .Y(_03353_));
 sky130_fd_sc_hd__nand3_2 _27153_ (.A(_03345_),
    .B(_03351_),
    .C(_11799_),
    .Y(_03354_));
 sky130_fd_sc_hd__nand2_2 _27154_ (.A(_03353_),
    .B(_03354_),
    .Y(_03356_));
 sky130_fd_sc_hd__inv_2 _27155_ (.A(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__nand2_1 _27156_ (.A(_03339_),
    .B(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__inv_2 _27157_ (.A(_03334_),
    .Y(_03359_));
 sky130_fd_sc_hd__a21boi_2 _27158_ (.A1(_03359_),
    .A2(_03354_),
    .B1_N(_03353_),
    .Y(_03360_));
 sky130_fd_sc_hd__nand2_2 _27159_ (.A(_03358_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__nand2_1 _27160_ (.A(_01626_),
    .B(_01713_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand3_1 _27161_ (.A(_01623_),
    .B(_01625_),
    .C(_01712_),
    .Y(_03363_));
 sky130_fd_sc_hd__nand2_1 _27162_ (.A(_03362_),
    .B(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__inv_2 _27163_ (.A(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__nand2_1 _27164_ (.A(net122),
    .B(_03365_),
    .Y(_03367_));
 sky130_fd_sc_hd__nand2_1 _27165_ (.A(_01603_),
    .B(_01599_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _27166_ (.A(_03368_),
    .B(_01622_),
    .Y(_03369_));
 sky130_fd_sc_hd__nand3_1 _27167_ (.A(_01603_),
    .B(_01621_),
    .C(_01599_),
    .Y(_03370_));
 sky130_fd_sc_hd__a21oi_1 _27168_ (.A1(_03369_),
    .A2(_03370_),
    .B1(_12047_),
    .Y(_03371_));
 sky130_fd_sc_hd__a21boi_2 _27169_ (.A1(_03347_),
    .A2(_03346_),
    .B1_N(_03348_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand2_1 _27170_ (.A(_03369_),
    .B(_03370_),
    .Y(_03373_));
 sky130_fd_sc_hd__inv_2 _27171_ (.A(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__nand2_1 _27172_ (.A(_03374_),
    .B(_12047_),
    .Y(_03375_));
 sky130_fd_sc_hd__o21ai_1 _27173_ (.A1(_03371_),
    .A2(_03372_),
    .B1(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__nand2_1 _27174_ (.A(_03364_),
    .B(_12056_),
    .Y(_03378_));
 sky130_fd_sc_hd__nand3_1 _27175_ (.A(_03362_),
    .B(_03363_),
    .C(_12058_),
    .Y(_03379_));
 sky130_fd_sc_hd__nand2_1 _27176_ (.A(_03378_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hd__inv_2 _27177_ (.A(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__or2_1 _27178_ (.A(_03376_),
    .B(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__nand2_1 _27179_ (.A(_03381_),
    .B(_03376_),
    .Y(_03383_));
 sky130_fd_sc_hd__nand2_1 _27180_ (.A(_03382_),
    .B(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__nand3b_1 _27181_ (.A_N(_03384_),
    .B(_02128_),
    .C(_02130_),
    .Y(_03385_));
 sky130_fd_sc_hd__a21o_1 _27182_ (.A1(_03367_),
    .A2(_03385_),
    .B1(_12261_),
    .X(_03386_));
 sky130_fd_sc_hd__nand3_1 _27183_ (.A(_03367_),
    .B(_03385_),
    .C(_12261_),
    .Y(_03387_));
 sky130_fd_sc_hd__nand2_1 _27184_ (.A(_03386_),
    .B(_03387_),
    .Y(_03389_));
 sky130_fd_sc_hd__or2b_1 _27185_ (.A(_03371_),
    .B_N(_03375_),
    .X(_03390_));
 sky130_fd_sc_hd__xnor2_1 _27186_ (.A(_03372_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__nand2_1 _27187_ (.A(net122),
    .B(_03374_),
    .Y(_03392_));
 sky130_fd_sc_hd__o21ai_2 _27188_ (.A1(_03391_),
    .A2(_02131_),
    .B1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__or2_4 _27189_ (.A(_12270_),
    .B(_03393_),
    .X(_03394_));
 sky130_fd_sc_hd__nand2_2 _27190_ (.A(_03393_),
    .B(_12270_),
    .Y(_03395_));
 sky130_fd_sc_hd__nand2_2 _27191_ (.A(_03394_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hd__nor2_4 _27192_ (.A(_03396_),
    .B(_03389_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _27193_ (.A(_03361_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__inv_2 _27194_ (.A(_03387_),
    .Y(_03400_));
 sky130_fd_sc_hd__o21ai_2 _27195_ (.A1(_03400_),
    .A2(_03395_),
    .B1(_03386_),
    .Y(_03401_));
 sky130_fd_sc_hd__inv_2 _27196_ (.A(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__nand2_1 _27197_ (.A(_03398_),
    .B(_03402_),
    .Y(_03403_));
 sky130_fd_sc_hd__inv_6 _27198_ (.A(_02131_),
    .Y(_03404_));
 sky130_fd_sc_hd__nand2_1 _27199_ (.A(_03362_),
    .B(_01710_),
    .Y(_03405_));
 sky130_fd_sc_hd__nand2_1 _27200_ (.A(_03405_),
    .B(_01703_),
    .Y(_03406_));
 sky130_fd_sc_hd__nand3_1 _27201_ (.A(_03362_),
    .B(_01702_),
    .C(_01710_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand2_1 _27202_ (.A(_03406_),
    .B(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__nand2_1 _27203_ (.A(_03408_),
    .B(_13182_),
    .Y(_03409_));
 sky130_fd_sc_hd__nand3_1 _27204_ (.A(_03406_),
    .B(_08176_),
    .C(_03407_),
    .Y(_03411_));
 sky130_fd_sc_hd__nand2_1 _27205_ (.A(_03409_),
    .B(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__nand2_1 _27206_ (.A(_03383_),
    .B(_03379_),
    .Y(_03413_));
 sky130_fd_sc_hd__xor2_1 _27207_ (.A(_03412_),
    .B(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__nand2_1 _27208_ (.A(_03404_),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__nand2_1 _27209_ (.A(_02132_),
    .B(_03408_),
    .Y(_03416_));
 sky130_fd_sc_hd__nand2_1 _27210_ (.A(_03415_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _27211_ (.A(_03417_),
    .B(_11496_),
    .Y(_03418_));
 sky130_fd_sc_hd__nand3_2 _27212_ (.A(_03415_),
    .B(_11494_),
    .C(_03416_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_2 _27213_ (.A(_03418_),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__clkinvlp_2 _27214_ (.A(_03420_),
    .Y(_03422_));
 sky130_fd_sc_hd__nand2_2 _27215_ (.A(_03403_),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__nand2_1 _27216_ (.A(_03423_),
    .B(_03419_),
    .Y(_03424_));
 sky130_fd_sc_hd__nand3_1 _27217_ (.A(_03383_),
    .B(_03411_),
    .C(_03379_),
    .Y(_03425_));
 sky130_fd_sc_hd__inv_2 _27218_ (.A(_01714_),
    .Y(_03426_));
 sky130_fd_sc_hd__nand2_1 _27219_ (.A(_01626_),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__inv_2 _27220_ (.A(_01719_),
    .Y(_03428_));
 sky130_fd_sc_hd__nand2_1 _27221_ (.A(_03427_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__nand2_1 _27222_ (.A(_03429_),
    .B(_01690_),
    .Y(_03430_));
 sky130_fd_sc_hd__nand3_1 _27223_ (.A(_03427_),
    .B(_01689_),
    .C(_03428_),
    .Y(_03431_));
 sky130_fd_sc_hd__nand2_1 _27224_ (.A(_03430_),
    .B(_03431_),
    .Y(_03433_));
 sky130_fd_sc_hd__nand2_1 _27225_ (.A(_03433_),
    .B(_12085_),
    .Y(_03434_));
 sky130_fd_sc_hd__nand3_1 _27226_ (.A(_03430_),
    .B(_12087_),
    .C(_03431_),
    .Y(_03435_));
 sky130_fd_sc_hd__nand2_1 _27227_ (.A(_03434_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__inv_4 _27228_ (.A(_03436_),
    .Y(_03437_));
 sky130_fd_sc_hd__a21o_1 _27229_ (.A1(_03425_),
    .A2(_03409_),
    .B1(_03437_),
    .X(_03438_));
 sky130_fd_sc_hd__nand3_2 _27230_ (.A(_03425_),
    .B(_03437_),
    .C(_03409_),
    .Y(_03439_));
 sky130_fd_sc_hd__nand2_1 _27231_ (.A(_03438_),
    .B(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__nand3b_1 _27232_ (.A_N(_03440_),
    .B(_02130_),
    .C(_02128_),
    .Y(_03441_));
 sky130_fd_sc_hd__inv_2 _27233_ (.A(_03433_),
    .Y(_03442_));
 sky130_fd_sc_hd__nand2_1 _27234_ (.A(_02132_),
    .B(_03442_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand2_1 _27235_ (.A(_03441_),
    .B(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__nand2_1 _27236_ (.A(_03445_),
    .B(_11482_),
    .Y(_03446_));
 sky130_fd_sc_hd__nand3_1 _27237_ (.A(_03441_),
    .B(_03444_),
    .C(_11484_),
    .Y(_03447_));
 sky130_fd_sc_hd__nand2_2 _27238_ (.A(_03446_),
    .B(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hd__clkinvlp_2 _27239_ (.A(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__nand2_1 _27240_ (.A(_03424_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hd__nand3_1 _27241_ (.A(_03423_),
    .B(_03448_),
    .C(_03419_),
    .Y(_03451_));
 sky130_fd_sc_hd__nand2_2 _27242_ (.A(_03450_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__nand2_2 _27243_ (.A(_03452_),
    .B(_13197_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand3_1 _27244_ (.A(_03450_),
    .B(_10939_),
    .C(_03451_),
    .Y(_03455_));
 sky130_fd_sc_hd__nand3_1 _27245_ (.A(_03398_),
    .B(_03420_),
    .C(_03402_),
    .Y(_03456_));
 sky130_fd_sc_hd__nand2_1 _27246_ (.A(_03423_),
    .B(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__nand2_1 _27247_ (.A(_03457_),
    .B(_12085_),
    .Y(_03458_));
 sky130_fd_sc_hd__nand3_2 _27248_ (.A(_03423_),
    .B(_12087_),
    .C(_03456_),
    .Y(_03459_));
 sky130_fd_sc_hd__nand2_1 _27249_ (.A(_03458_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hd__inv_2 _27250_ (.A(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__nand3_1 _27251_ (.A(_03453_),
    .B(_03455_),
    .C(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__inv_2 _27252_ (.A(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__nand2_1 _27253_ (.A(_03338_),
    .B(_03334_),
    .Y(_03464_));
 sky130_fd_sc_hd__xor2_1 _27254_ (.A(_03356_),
    .B(_03464_),
    .X(_03466_));
 sky130_fd_sc_hd__or2_1 _27255_ (.A(_12043_),
    .B(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__nand2_1 _27256_ (.A(_03334_),
    .B(_03335_),
    .Y(_03468_));
 sky130_fd_sc_hd__nand2_1 _27257_ (.A(_03468_),
    .B(_03336_),
    .Y(_03469_));
 sky130_fd_sc_hd__nand2_1 _27258_ (.A(_03469_),
    .B(_03338_),
    .Y(_03470_));
 sky130_fd_sc_hd__nand2_1 _27259_ (.A(_03470_),
    .B(_12030_),
    .Y(_03471_));
 sky130_fd_sc_hd__o21ai_1 _27260_ (.A1(_00161_),
    .A2(\div1i.quot[0] ),
    .B1(_00174_),
    .Y(_03472_));
 sky130_fd_sc_hd__nand3_1 _27261_ (.A(_03469_),
    .B(_12035_),
    .C(_03338_),
    .Y(_03473_));
 sky130_fd_sc_hd__inv_2 _27262_ (.A(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__a21o_1 _27263_ (.A1(_03471_),
    .A2(_03472_),
    .B1(_03474_),
    .X(_03475_));
 sky130_fd_sc_hd__nand2_1 _27264_ (.A(_03466_),
    .B(_12043_),
    .Y(_03477_));
 sky130_fd_sc_hd__nand2_1 _27265_ (.A(_03475_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__nand2_1 _27266_ (.A(_03467_),
    .B(_03478_),
    .Y(_03479_));
 sky130_fd_sc_hd__inv_2 _27267_ (.A(_03396_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2_2 _27268_ (.A(_03361_),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__nand3_1 _27269_ (.A(_03358_),
    .B(_03360_),
    .C(_03396_),
    .Y(_03482_));
 sky130_fd_sc_hd__nand2_1 _27270_ (.A(_03481_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hd__nand2_1 _27271_ (.A(_03483_),
    .B(_12056_),
    .Y(_03484_));
 sky130_fd_sc_hd__nand3_1 _27272_ (.A(_03481_),
    .B(_03482_),
    .C(_12058_),
    .Y(_03485_));
 sky130_fd_sc_hd__nand2_1 _27273_ (.A(_03484_),
    .B(_03485_),
    .Y(_03486_));
 sky130_fd_sc_hd__inv_2 _27274_ (.A(_03486_),
    .Y(_03488_));
 sky130_fd_sc_hd__nand2_1 _27275_ (.A(_03479_),
    .B(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__nand2_1 _27276_ (.A(_03489_),
    .B(_03485_),
    .Y(_03490_));
 sky130_fd_sc_hd__inv_2 _27277_ (.A(_03389_),
    .Y(_03491_));
 sky130_fd_sc_hd__nand2_1 _27278_ (.A(_03481_),
    .B(_03395_),
    .Y(_03492_));
 sky130_fd_sc_hd__or2_1 _27279_ (.A(_03491_),
    .B(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__nand2_1 _27280_ (.A(_03492_),
    .B(_03491_),
    .Y(_03494_));
 sky130_fd_sc_hd__nand2_1 _27281_ (.A(_03493_),
    .B(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__nand2_1 _27282_ (.A(_03495_),
    .B(_13182_),
    .Y(_03496_));
 sky130_fd_sc_hd__nand2_1 _27283_ (.A(_03490_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__nand3_1 _27284_ (.A(_03493_),
    .B(_08176_),
    .C(_03494_),
    .Y(_03499_));
 sky130_fd_sc_hd__nand2_1 _27285_ (.A(_03497_),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__nand2_1 _27286_ (.A(_03463_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__inv_2 _27287_ (.A(_03459_),
    .Y(_03502_));
 sky130_fd_sc_hd__a21boi_1 _27288_ (.A1(_03453_),
    .A2(_03502_),
    .B1_N(_03455_),
    .Y(_03503_));
 sky130_fd_sc_hd__nand2_1 _27289_ (.A(_03501_),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__nor2_2 _27290_ (.A(_03448_),
    .B(_03420_),
    .Y(_03505_));
 sky130_fd_sc_hd__nand3_2 _27291_ (.A(_03361_),
    .B(_03397_),
    .C(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__o21ai_1 _27292_ (.A1(_03419_),
    .A2(_03448_),
    .B1(_03446_),
    .Y(_03507_));
 sky130_fd_sc_hd__a21oi_2 _27293_ (.A1(_03401_),
    .A2(_03505_),
    .B1(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__nand2_4 _27294_ (.A(_03506_),
    .B(_03508_),
    .Y(_03510_));
 sky130_fd_sc_hd__nand2_1 _27295_ (.A(_03430_),
    .B(_01687_),
    .Y(_03511_));
 sky130_fd_sc_hd__or2_1 _27296_ (.A(_01680_),
    .B(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__nand2_1 _27297_ (.A(_03511_),
    .B(_01680_),
    .Y(_03513_));
 sky130_fd_sc_hd__nand3_1 _27298_ (.A(net122),
    .B(_03512_),
    .C(_03513_),
    .Y(_03514_));
 sky130_fd_sc_hd__nand2_1 _27299_ (.A(_03439_),
    .B(_03435_),
    .Y(_03515_));
 sky130_fd_sc_hd__nand2_1 _27300_ (.A(_03512_),
    .B(_03513_),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_1 _27301_ (.A(_03516_),
    .B(_13197_),
    .Y(_03517_));
 sky130_fd_sc_hd__nand3_2 _27302_ (.A(_03512_),
    .B(_10939_),
    .C(_03513_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2_2 _27303_ (.A(_03518_),
    .B(_03517_),
    .Y(_03519_));
 sky130_fd_sc_hd__inv_2 _27304_ (.A(_03519_),
    .Y(_03521_));
 sky130_fd_sc_hd__nand2_1 _27305_ (.A(_03515_),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__nand3_1 _27306_ (.A(_03519_),
    .B(_03439_),
    .C(_03435_),
    .Y(_03523_));
 sky130_fd_sc_hd__nand2_1 _27307_ (.A(_03522_),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__inv_2 _27308_ (.A(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__nand2_1 _27309_ (.A(_03404_),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__nand2_1 _27310_ (.A(_03514_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__nand2_1 _27311_ (.A(_03527_),
    .B(_08951_),
    .Y(_03528_));
 sky130_fd_sc_hd__nand3_1 _27312_ (.A(_03514_),
    .B(_03526_),
    .C(_12771_),
    .Y(_03529_));
 sky130_fd_sc_hd__nand2_2 _27313_ (.A(_03528_),
    .B(_03529_),
    .Y(_03530_));
 sky130_fd_sc_hd__inv_2 _27314_ (.A(_03530_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand2_1 _27315_ (.A(_03510_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__inv_2 _27316_ (.A(_01763_),
    .Y(_03534_));
 sky130_fd_sc_hd__or2_1 _27317_ (.A(_03534_),
    .B(_01724_),
    .X(_03535_));
 sky130_fd_sc_hd__nand2_1 _27318_ (.A(_01724_),
    .B(_03534_),
    .Y(_03536_));
 sky130_fd_sc_hd__nand2_1 _27319_ (.A(_03535_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hd__inv_2 _27320_ (.A(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hd__nand2_1 _27321_ (.A(_03538_),
    .B(_12008_),
    .Y(_03539_));
 sky130_fd_sc_hd__nand2_1 _27322_ (.A(_03537_),
    .B(_12101_),
    .Y(_03540_));
 sky130_fd_sc_hd__nand2_1 _27323_ (.A(_03539_),
    .B(_03540_),
    .Y(_03541_));
 sky130_fd_sc_hd__inv_2 _27324_ (.A(_03541_),
    .Y(_03543_));
 sky130_fd_sc_hd__nand2_2 _27325_ (.A(_03522_),
    .B(_03518_),
    .Y(_03544_));
 sky130_fd_sc_hd__or2_1 _27326_ (.A(_03543_),
    .B(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__nand2_1 _27327_ (.A(_03544_),
    .B(_03543_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand3_1 _27328_ (.A(_03545_),
    .B(_03404_),
    .C(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__nand2_1 _27329_ (.A(_02132_),
    .B(_03538_),
    .Y(_03548_));
 sky130_fd_sc_hd__nand2_1 _27330_ (.A(_03547_),
    .B(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__nand2_1 _27331_ (.A(_03549_),
    .B(_11614_),
    .Y(_03550_));
 sky130_fd_sc_hd__nand3_2 _27332_ (.A(_03547_),
    .B(_11616_),
    .C(_03548_),
    .Y(_03551_));
 sky130_fd_sc_hd__nand2_1 _27333_ (.A(_03550_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__a21o_1 _27334_ (.A1(_03533_),
    .A2(_03528_),
    .B1(_03552_),
    .X(_03554_));
 sky130_fd_sc_hd__nand3_1 _27335_ (.A(_03533_),
    .B(_03552_),
    .C(_03528_),
    .Y(_03555_));
 sky130_fd_sc_hd__nand2_1 _27336_ (.A(_03554_),
    .B(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__nand2_1 _27337_ (.A(_03556_),
    .B(_12002_),
    .Y(_03557_));
 sky130_fd_sc_hd__xor2_1 _27338_ (.A(_03530_),
    .B(_03510_),
    .X(_03558_));
 sky130_fd_sc_hd__nand2_1 _27339_ (.A(_03558_),
    .B(_12101_),
    .Y(_03559_));
 sky130_fd_sc_hd__or2_1 _27340_ (.A(_03532_),
    .B(_03510_),
    .X(_03560_));
 sky130_fd_sc_hd__nand3_2 _27341_ (.A(_03560_),
    .B(_12008_),
    .C(_03533_),
    .Y(_03561_));
 sky130_fd_sc_hd__nand2_1 _27342_ (.A(_03559_),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__inv_2 _27343_ (.A(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__nand3_1 _27344_ (.A(_03554_),
    .B(_12012_),
    .C(_03555_),
    .Y(_03565_));
 sky130_fd_sc_hd__nand3_1 _27345_ (.A(_03557_),
    .B(_03563_),
    .C(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hd__inv_2 _27346_ (.A(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__nand2_1 _27347_ (.A(_03504_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__inv_2 _27348_ (.A(_03561_),
    .Y(_03569_));
 sky130_fd_sc_hd__a21boi_1 _27349_ (.A1(_03557_),
    .A2(_03569_),
    .B1_N(_03565_),
    .Y(_03570_));
 sky130_fd_sc_hd__nand2_1 _27350_ (.A(_03568_),
    .B(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hd__nand2_1 _27351_ (.A(_03536_),
    .B(_01761_),
    .Y(_03572_));
 sky130_fd_sc_hd__xor2_1 _27352_ (.A(_01752_),
    .B(_03572_),
    .X(_03573_));
 sky130_fd_sc_hd__nand2_1 _27353_ (.A(_03573_),
    .B(_12002_),
    .Y(_03574_));
 sky130_fd_sc_hd__inv_2 _27354_ (.A(_01752_),
    .Y(_03576_));
 sky130_fd_sc_hd__or2_1 _27355_ (.A(_03576_),
    .B(_03572_),
    .X(_03577_));
 sky130_fd_sc_hd__nand2_1 _27356_ (.A(_03572_),
    .B(_03576_),
    .Y(_03578_));
 sky130_fd_sc_hd__nand3_1 _27357_ (.A(_03577_),
    .B(_12012_),
    .C(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__nand2_1 _27358_ (.A(_03574_),
    .B(_03579_),
    .Y(_03580_));
 sky130_fd_sc_hd__inv_2 _27359_ (.A(_03580_),
    .Y(_03581_));
 sky130_fd_sc_hd__nand2_1 _27360_ (.A(_03581_),
    .B(_03543_),
    .Y(_03582_));
 sky130_fd_sc_hd__inv_2 _27361_ (.A(_03582_),
    .Y(_03583_));
 sky130_fd_sc_hd__nand2_1 _27362_ (.A(_03544_),
    .B(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__inv_2 _27363_ (.A(_03539_),
    .Y(_03585_));
 sky130_fd_sc_hd__inv_2 _27364_ (.A(_03579_),
    .Y(_03587_));
 sky130_fd_sc_hd__a21oi_2 _27365_ (.A1(_03574_),
    .A2(_03585_),
    .B1(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__nand2_1 _27366_ (.A(_03584_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__nand2_1 _27367_ (.A(_01724_),
    .B(_01764_),
    .Y(_03590_));
 sky130_fd_sc_hd__inv_2 _27368_ (.A(_01816_),
    .Y(_03591_));
 sky130_fd_sc_hd__nand2_1 _27369_ (.A(_03590_),
    .B(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__clkinvlp_2 _27370_ (.A(_01810_),
    .Y(_03593_));
 sky130_fd_sc_hd__nand2_1 _27371_ (.A(_03592_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__nand3_1 _27372_ (.A(_03590_),
    .B(_01810_),
    .C(_03591_),
    .Y(_03595_));
 sky130_fd_sc_hd__nand2_1 _27373_ (.A(_03594_),
    .B(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__nand2_1 _27374_ (.A(_03596_),
    .B(_12017_),
    .Y(_03598_));
 sky130_fd_sc_hd__nand3_2 _27375_ (.A(_03594_),
    .B(_11986_),
    .C(_03595_),
    .Y(_03599_));
 sky130_fd_sc_hd__nand2_1 _27376_ (.A(_03598_),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__inv_2 _27377_ (.A(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__nand2_1 _27378_ (.A(_03589_),
    .B(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__nand3_1 _27379_ (.A(_03584_),
    .B(_03600_),
    .C(_03588_),
    .Y(_03603_));
 sky130_fd_sc_hd__nand3_1 _27380_ (.A(_03602_),
    .B(_03404_),
    .C(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__or2_1 _27381_ (.A(_03596_),
    .B(_03404_),
    .X(_03605_));
 sky130_fd_sc_hd__nand2_1 _27382_ (.A(_03604_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__nand2_1 _27383_ (.A(_03606_),
    .B(_11586_),
    .Y(_03607_));
 sky130_fd_sc_hd__nand3_1 _27384_ (.A(_03604_),
    .B(_11588_),
    .C(_03605_),
    .Y(_03609_));
 sky130_fd_sc_hd__nand2_2 _27385_ (.A(_03607_),
    .B(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__nand3_1 _27386_ (.A(_03532_),
    .B(_03550_),
    .C(_03551_),
    .Y(_03611_));
 sky130_fd_sc_hd__inv_2 _27387_ (.A(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__nand2_1 _27388_ (.A(_03510_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__inv_2 _27389_ (.A(_03551_),
    .Y(_03614_));
 sky130_fd_sc_hd__o21ai_1 _27390_ (.A1(_03528_),
    .A2(_03614_),
    .B1(_03550_),
    .Y(_03615_));
 sky130_fd_sc_hd__inv_2 _27391_ (.A(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_2 _27392_ (.A(_03613_),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2_1 _27393_ (.A(_03546_),
    .B(_03539_),
    .Y(_03618_));
 sky130_fd_sc_hd__nand2_1 _27394_ (.A(_03618_),
    .B(_03581_),
    .Y(_03620_));
 sky130_fd_sc_hd__nand3_1 _27395_ (.A(_03546_),
    .B(_03580_),
    .C(_03539_),
    .Y(_03621_));
 sky130_fd_sc_hd__nand2_1 _27396_ (.A(_03620_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__nand2_1 _27397_ (.A(_03622_),
    .B(_03404_),
    .Y(_03623_));
 sky130_fd_sc_hd__nand2_1 _27398_ (.A(_02132_),
    .B(_03573_),
    .Y(_03624_));
 sky130_fd_sc_hd__nand2_1 _27399_ (.A(_03623_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__nand2_1 _27400_ (.A(_03625_),
    .B(_11600_),
    .Y(_03626_));
 sky130_fd_sc_hd__nand3_2 _27401_ (.A(_03623_),
    .B(_11603_),
    .C(_03624_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand2_2 _27402_ (.A(_03626_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__inv_2 _27403_ (.A(_03628_),
    .Y(_03629_));
 sky130_fd_sc_hd__nand2_2 _27404_ (.A(_03617_),
    .B(_03629_),
    .Y(_03631_));
 sky130_fd_sc_hd__nand2_1 _27405_ (.A(_03631_),
    .B(_03627_),
    .Y(_03632_));
 sky130_fd_sc_hd__xor2_1 _27406_ (.A(_03610_),
    .B(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__nand2_2 _27407_ (.A(_03633_),
    .B(_11983_),
    .Y(_03634_));
 sky130_fd_sc_hd__inv_2 _27408_ (.A(_03610_),
    .Y(_03635_));
 sky130_fd_sc_hd__or2_1 _27409_ (.A(_03635_),
    .B(_03632_),
    .X(_03636_));
 sky130_fd_sc_hd__nand2_1 _27410_ (.A(_03632_),
    .B(_03635_),
    .Y(_03637_));
 sky130_fd_sc_hd__nand3_2 _27411_ (.A(_03636_),
    .B(_11990_),
    .C(_03637_),
    .Y(_03638_));
 sky130_fd_sc_hd__xor2_1 _27412_ (.A(_03628_),
    .B(_03617_),
    .X(_03639_));
 sky130_fd_sc_hd__nand2_1 _27413_ (.A(_03639_),
    .B(_12017_),
    .Y(_03640_));
 sky130_fd_sc_hd__or2_1 _27414_ (.A(_03629_),
    .B(_03617_),
    .X(_03642_));
 sky130_fd_sc_hd__nand3_2 _27415_ (.A(_03642_),
    .B(_11986_),
    .C(_03631_),
    .Y(_03643_));
 sky130_fd_sc_hd__nand2_1 _27416_ (.A(_03640_),
    .B(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__inv_2 _27417_ (.A(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hd__nand3_2 _27418_ (.A(_03634_),
    .B(_03638_),
    .C(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__inv_2 _27419_ (.A(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__nand2_1 _27420_ (.A(_03571_),
    .B(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__inv_2 _27421_ (.A(_03643_),
    .Y(_03649_));
 sky130_fd_sc_hd__a21boi_2 _27422_ (.A1(_03634_),
    .A2(_03649_),
    .B1_N(_03638_),
    .Y(_03650_));
 sky130_fd_sc_hd__nand2_1 _27423_ (.A(_03648_),
    .B(_03650_),
    .Y(_03651_));
 sky130_fd_sc_hd__nand2_1 _27424_ (.A(_03602_),
    .B(_03599_),
    .Y(_03653_));
 sky130_fd_sc_hd__nand2_1 _27425_ (.A(_03594_),
    .B(_01809_),
    .Y(_03654_));
 sky130_fd_sc_hd__clkinvlp_2 _27426_ (.A(_01800_),
    .Y(_03655_));
 sky130_fd_sc_hd__nand2_1 _27427_ (.A(_03654_),
    .B(_03655_),
    .Y(_03656_));
 sky130_fd_sc_hd__nand3_1 _27428_ (.A(_03594_),
    .B(_01800_),
    .C(_01809_),
    .Y(_03657_));
 sky130_fd_sc_hd__nand2_1 _27429_ (.A(_03656_),
    .B(_03657_),
    .Y(_03658_));
 sky130_fd_sc_hd__nand2_1 _27430_ (.A(_03658_),
    .B(_11983_),
    .Y(_03659_));
 sky130_fd_sc_hd__nand3_1 _27431_ (.A(_03656_),
    .B(_11990_),
    .C(_03657_),
    .Y(_03660_));
 sky130_fd_sc_hd__nand2_1 _27432_ (.A(_03659_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__inv_2 _27433_ (.A(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__nand2_1 _27434_ (.A(_03653_),
    .B(_03662_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand3_1 _27435_ (.A(_03602_),
    .B(_03661_),
    .C(_03599_),
    .Y(_03665_));
 sky130_fd_sc_hd__nand2_1 _27436_ (.A(_03664_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__nand2_1 _27437_ (.A(_03666_),
    .B(_03404_),
    .Y(_03667_));
 sky130_fd_sc_hd__nand2_1 _27438_ (.A(net239),
    .B(_03658_),
    .Y(_03668_));
 sky130_fd_sc_hd__a21o_1 _27439_ (.A1(_03667_),
    .A2(_03668_),
    .B1(_12187_),
    .X(_03669_));
 sky130_fd_sc_hd__nand3_2 _27440_ (.A(_03667_),
    .B(_12187_),
    .C(_03668_),
    .Y(_03670_));
 sky130_fd_sc_hd__nand2_1 _27441_ (.A(_03669_),
    .B(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hd__inv_2 _27442_ (.A(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__nor3_1 _27443_ (.A(_03610_),
    .B(_03611_),
    .C(_03628_),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2_1 _27444_ (.A(_03673_),
    .B(_03510_),
    .Y(_03675_));
 sky130_fd_sc_hd__nor2_1 _27445_ (.A(_03610_),
    .B(_03628_),
    .Y(_03676_));
 sky130_fd_sc_hd__inv_2 _27446_ (.A(_03609_),
    .Y(_03677_));
 sky130_fd_sc_hd__o21ai_1 _27447_ (.A1(_03627_),
    .A2(_03677_),
    .B1(_03607_),
    .Y(_03678_));
 sky130_fd_sc_hd__a21oi_1 _27448_ (.A1(_03676_),
    .A2(_03615_),
    .B1(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__nand2_2 _27449_ (.A(_03675_),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__or2_1 _27450_ (.A(_03672_),
    .B(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__nand2_2 _27451_ (.A(_03680_),
    .B(_03672_),
    .Y(_03682_));
 sky130_fd_sc_hd__nand2_1 _27452_ (.A(_03681_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__nor2_1 _27453_ (.A(_12817_),
    .B(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__inv_2 _27454_ (.A(_03684_),
    .Y(_03686_));
 sky130_fd_sc_hd__nand2_1 _27455_ (.A(_03683_),
    .B(_12817_),
    .Y(_03687_));
 sky130_fd_sc_hd__nand2_1 _27456_ (.A(_03686_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__inv_2 _27457_ (.A(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__nand2_1 _27458_ (.A(_03682_),
    .B(_03670_),
    .Y(_03690_));
 sky130_fd_sc_hd__clkinvlp_2 _27459_ (.A(_01913_),
    .Y(_03691_));
 sky130_fd_sc_hd__or2_1 _27460_ (.A(_03691_),
    .B(_01819_),
    .X(_03692_));
 sky130_fd_sc_hd__nand2_1 _27461_ (.A(_01819_),
    .B(_03691_),
    .Y(_03693_));
 sky130_fd_sc_hd__nand2_1 _27462_ (.A(_03692_),
    .B(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__inv_2 _27463_ (.A(_03694_),
    .Y(_03695_));
 sky130_fd_sc_hd__nand2_1 _27464_ (.A(_03695_),
    .B(_11671_),
    .Y(_03697_));
 sky130_fd_sc_hd__nand2_1 _27465_ (.A(_03694_),
    .B(_12817_),
    .Y(_03698_));
 sky130_fd_sc_hd__nand2_1 _27466_ (.A(_03697_),
    .B(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__inv_4 _27467_ (.A(_03699_),
    .Y(_03700_));
 sky130_fd_sc_hd__nand3_1 _27468_ (.A(_03659_),
    .B(_03660_),
    .C(_03601_),
    .Y(_03701_));
 sky130_fd_sc_hd__inv_2 _27469_ (.A(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__nand3_1 _27470_ (.A(_03544_),
    .B(_03702_),
    .C(_03583_),
    .Y(_03703_));
 sky130_fd_sc_hd__inv_2 _27471_ (.A(_03599_),
    .Y(_03704_));
 sky130_fd_sc_hd__inv_2 _27472_ (.A(_03660_),
    .Y(_03705_));
 sky130_fd_sc_hd__a21o_1 _27473_ (.A1(_03659_),
    .A2(_03704_),
    .B1(_03705_),
    .X(_03706_));
 sky130_fd_sc_hd__nor2_1 _27474_ (.A(_03588_),
    .B(_03701_),
    .Y(_03708_));
 sky130_fd_sc_hd__nor2_1 _27475_ (.A(_03706_),
    .B(_03708_),
    .Y(_03709_));
 sky130_fd_sc_hd__nand2_1 _27476_ (.A(_03703_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__or2_1 _27477_ (.A(_03700_),
    .B(_03710_),
    .X(_03711_));
 sky130_fd_sc_hd__nand2_1 _27478_ (.A(_03710_),
    .B(_03700_),
    .Y(_03712_));
 sky130_fd_sc_hd__nand3_1 _27479_ (.A(_03711_),
    .B(_03404_),
    .C(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__nand2_1 _27480_ (.A(net239),
    .B(_03695_),
    .Y(_03714_));
 sky130_fd_sc_hd__a21o_1 _27481_ (.A1(_03713_),
    .A2(_03714_),
    .B1(_13304_),
    .X(_03715_));
 sky130_fd_sc_hd__nand3_1 _27482_ (.A(_03713_),
    .B(_13304_),
    .C(_03714_),
    .Y(_03716_));
 sky130_fd_sc_hd__nand2_1 _27483_ (.A(_03715_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__inv_2 _27484_ (.A(_03717_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _27485_ (.A(_03690_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand3_1 _27486_ (.A(_03682_),
    .B(_03717_),
    .C(_03670_),
    .Y(_03721_));
 sky130_fd_sc_hd__nand2_1 _27487_ (.A(_03720_),
    .B(_03721_),
    .Y(_03722_));
 sky130_fd_sc_hd__nand2_1 _27488_ (.A(_03722_),
    .B(_12118_),
    .Y(_03723_));
 sky130_fd_sc_hd__nand3_1 _27489_ (.A(_03720_),
    .B(_12120_),
    .C(_03721_),
    .Y(_03724_));
 sky130_fd_sc_hd__nand2_2 _27490_ (.A(_03723_),
    .B(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__inv_2 _27491_ (.A(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__nand2_1 _27492_ (.A(_03689_),
    .B(_03726_),
    .Y(_03727_));
 sky130_fd_sc_hd__nor2_1 _27493_ (.A(_03717_),
    .B(_03671_),
    .Y(_03728_));
 sky130_fd_sc_hd__nand2_1 _27494_ (.A(_03680_),
    .B(_03728_),
    .Y(_03730_));
 sky130_fd_sc_hd__inv_2 _27495_ (.A(_03716_),
    .Y(_03731_));
 sky130_fd_sc_hd__o21ai_1 _27496_ (.A1(_03670_),
    .A2(_03731_),
    .B1(_03715_),
    .Y(_03732_));
 sky130_fd_sc_hd__inv_2 _27497_ (.A(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand2_1 _27498_ (.A(_03730_),
    .B(_03733_),
    .Y(_03734_));
 sky130_fd_sc_hd__nand2_1 _27499_ (.A(_03712_),
    .B(_03697_),
    .Y(_03735_));
 sky130_fd_sc_hd__nand2_1 _27500_ (.A(_03693_),
    .B(_01912_),
    .Y(_03736_));
 sky130_fd_sc_hd__xor2_1 _27501_ (.A(_01902_),
    .B(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__nand2b_1 _27502_ (.A_N(_03737_),
    .B(_12120_),
    .Y(_03738_));
 sky130_fd_sc_hd__nand2_1 _27503_ (.A(_03737_),
    .B(_12118_),
    .Y(_03739_));
 sky130_fd_sc_hd__nand2_1 _27504_ (.A(_03738_),
    .B(_03739_),
    .Y(_03741_));
 sky130_fd_sc_hd__inv_2 _27505_ (.A(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__nand2_1 _27506_ (.A(_03735_),
    .B(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand3_1 _27507_ (.A(_03712_),
    .B(_03741_),
    .C(_03697_),
    .Y(_03744_));
 sky130_fd_sc_hd__nand2_1 _27508_ (.A(_03743_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__buf_6 _27509_ (.A(_03404_),
    .X(_03746_));
 sky130_fd_sc_hd__nand2_1 _27510_ (.A(_03745_),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand2_1 _27511_ (.A(net239),
    .B(_03737_),
    .Y(_03748_));
 sky130_fd_sc_hd__nand2_1 _27512_ (.A(_03747_),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__nand2_1 _27513_ (.A(_03749_),
    .B(_11715_),
    .Y(_03750_));
 sky130_fd_sc_hd__nand3_2 _27514_ (.A(_03747_),
    .B(_11717_),
    .C(_03748_),
    .Y(_03752_));
 sky130_fd_sc_hd__nand2_1 _27515_ (.A(_03750_),
    .B(_03752_),
    .Y(_03753_));
 sky130_fd_sc_hd__inv_2 _27516_ (.A(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2_2 _27517_ (.A(_03734_),
    .B(_03754_),
    .Y(_03755_));
 sky130_fd_sc_hd__nand2_1 _27518_ (.A(_03755_),
    .B(_03752_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_1 _27519_ (.A(_03742_),
    .B(_03700_),
    .Y(_03757_));
 sky130_fd_sc_hd__inv_2 _27520_ (.A(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2_1 _27521_ (.A(_03710_),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__o21a_1 _27522_ (.A1(_03697_),
    .A2(_03741_),
    .B1(_03738_),
    .X(_03760_));
 sky130_fd_sc_hd__nand2_1 _27523_ (.A(_03759_),
    .B(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__a21o_1 _27524_ (.A1(_01819_),
    .A2(_01915_),
    .B1(_01919_),
    .X(_03763_));
 sky130_fd_sc_hd__xor2_1 _27525_ (.A(_01894_),
    .B(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__inv_2 _27526_ (.A(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__nand2_1 _27527_ (.A(_03765_),
    .B(_12147_),
    .Y(_03766_));
 sky130_fd_sc_hd__nand2_1 _27528_ (.A(_03764_),
    .B(_12149_),
    .Y(_03767_));
 sky130_fd_sc_hd__nand2_1 _27529_ (.A(_03766_),
    .B(_03767_),
    .Y(_03768_));
 sky130_fd_sc_hd__inv_2 _27530_ (.A(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__nand2_1 _27531_ (.A(_03761_),
    .B(_03769_),
    .Y(_03770_));
 sky130_fd_sc_hd__nand3_1 _27532_ (.A(_03759_),
    .B(_03768_),
    .C(_03760_),
    .Y(_03771_));
 sky130_fd_sc_hd__nand3_1 _27533_ (.A(_03770_),
    .B(_03746_),
    .C(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__nand2_1 _27534_ (.A(net239),
    .B(_03765_),
    .Y(_03774_));
 sky130_fd_sc_hd__nand2_1 _27535_ (.A(_03772_),
    .B(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__nand2_1 _27536_ (.A(_03775_),
    .B(_11701_),
    .Y(_03776_));
 sky130_fd_sc_hd__nand3_1 _27537_ (.A(_03772_),
    .B(_11703_),
    .C(_03774_),
    .Y(_03777_));
 sky130_fd_sc_hd__nand2_1 _27538_ (.A(_03776_),
    .B(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__inv_2 _27539_ (.A(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__nand2_1 _27540_ (.A(_03756_),
    .B(_03779_),
    .Y(_03780_));
 sky130_fd_sc_hd__nand3_1 _27541_ (.A(_03755_),
    .B(_03778_),
    .C(_03752_),
    .Y(_03781_));
 sky130_fd_sc_hd__nand2_1 _27542_ (.A(_03780_),
    .B(_03781_),
    .Y(_03782_));
 sky130_fd_sc_hd__nand2_1 _27543_ (.A(_03782_),
    .B(_12894_),
    .Y(_03783_));
 sky130_fd_sc_hd__nand3_1 _27544_ (.A(_03730_),
    .B(_03753_),
    .C(_03733_),
    .Y(_03785_));
 sky130_fd_sc_hd__nand2_1 _27545_ (.A(_03755_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__nand2_1 _27546_ (.A(_03786_),
    .B(_12149_),
    .Y(_03787_));
 sky130_fd_sc_hd__nand3_2 _27547_ (.A(_03755_),
    .B(_12147_),
    .C(_03785_),
    .Y(_03788_));
 sky130_fd_sc_hd__nand2_1 _27548_ (.A(_03787_),
    .B(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__inv_2 _27549_ (.A(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__nand3_2 _27550_ (.A(_03780_),
    .B(_11754_),
    .C(_03781_),
    .Y(_03791_));
 sky130_fd_sc_hd__nand3_1 _27551_ (.A(_03783_),
    .B(_03790_),
    .C(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__nor2_1 _27552_ (.A(_03727_),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__nand2_1 _27553_ (.A(_03651_),
    .B(_03793_),
    .Y(_03794_));
 sky130_fd_sc_hd__clkinvlp_2 _27554_ (.A(_03788_),
    .Y(_03796_));
 sky130_fd_sc_hd__nand3_1 _27555_ (.A(_03783_),
    .B(_03796_),
    .C(_03791_),
    .Y(_03797_));
 sky130_fd_sc_hd__nand2_1 _27556_ (.A(_03797_),
    .B(_03791_),
    .Y(_03798_));
 sky130_fd_sc_hd__a21boi_2 _27557_ (.A1(_03723_),
    .A2(_03684_),
    .B1_N(_03724_),
    .Y(_03799_));
 sky130_fd_sc_hd__nor2_1 _27558_ (.A(_03799_),
    .B(_03792_),
    .Y(_03800_));
 sky130_fd_sc_hd__nor2_2 _27559_ (.A(_03798_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__nand2_2 _27560_ (.A(_03794_),
    .B(_03801_),
    .Y(_03802_));
 sky130_fd_sc_hd__nand2_1 _27561_ (.A(_03770_),
    .B(_03766_),
    .Y(_03803_));
 sky130_fd_sc_hd__a21bo_1 _27562_ (.A1(_03763_),
    .A2(_01891_),
    .B1_N(_01893_),
    .X(_03804_));
 sky130_fd_sc_hd__xor2_1 _27563_ (.A(_01882_),
    .B(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__or2_1 _27564_ (.A(_12894_),
    .B(_03805_),
    .X(_03807_));
 sky130_fd_sc_hd__nand2_1 _27565_ (.A(_03805_),
    .B(_12894_),
    .Y(_03808_));
 sky130_fd_sc_hd__nand2_1 _27566_ (.A(_03807_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__inv_2 _27567_ (.A(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__nand2_1 _27568_ (.A(_03803_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2_1 _27569_ (.A(_03811_),
    .B(_03807_),
    .Y(_03812_));
 sky130_fd_sc_hd__nand2_1 _27570_ (.A(_02011_),
    .B(_02012_),
    .Y(_03813_));
 sky130_fd_sc_hd__xor2_1 _27571_ (.A(_03813_),
    .B(_01922_),
    .X(_03814_));
 sky130_fd_sc_hd__or2_1 _27572_ (.A(_13461_),
    .B(_03814_),
    .X(_03815_));
 sky130_fd_sc_hd__nand2_1 _27573_ (.A(_03814_),
    .B(_13461_),
    .Y(_03816_));
 sky130_fd_sc_hd__nand2_1 _27574_ (.A(_03815_),
    .B(_03816_),
    .Y(_03818_));
 sky130_fd_sc_hd__inv_2 _27575_ (.A(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__nand2_2 _27576_ (.A(_03812_),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__nand3_1 _27577_ (.A(_03811_),
    .B(_03818_),
    .C(_03807_),
    .Y(_03821_));
 sky130_fd_sc_hd__nand2_1 _27578_ (.A(_03820_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__nand2_1 _27579_ (.A(_03822_),
    .B(_03746_),
    .Y(_03823_));
 sky130_fd_sc_hd__nand2_1 _27580_ (.A(\div1i.quot[0] ),
    .B(_03814_),
    .Y(_03824_));
 sky130_fd_sc_hd__nand2_1 _27581_ (.A(_03823_),
    .B(_03824_),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2_1 _27582_ (.A(_03825_),
    .B(_06754_),
    .Y(_03826_));
 sky130_fd_sc_hd__nand3_1 _27583_ (.A(_03823_),
    .B(_13502_),
    .C(_03824_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_1 _27584_ (.A(_03826_),
    .B(_03827_),
    .Y(_03829_));
 sky130_fd_sc_hd__clkinvlp_2 _27585_ (.A(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__nor2_1 _27586_ (.A(_03778_),
    .B(_03753_),
    .Y(_03831_));
 sky130_fd_sc_hd__nand3_1 _27587_ (.A(_03680_),
    .B(_03831_),
    .C(_03728_),
    .Y(_03832_));
 sky130_fd_sc_hd__inv_2 _27588_ (.A(_03777_),
    .Y(_03833_));
 sky130_fd_sc_hd__o21ai_1 _27589_ (.A1(_03752_),
    .A2(_03833_),
    .B1(_03776_),
    .Y(_03834_));
 sky130_fd_sc_hd__a21oi_1 _27590_ (.A1(_03831_),
    .A2(_03732_),
    .B1(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hd__nand2_2 _27591_ (.A(_03832_),
    .B(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__xor2_1 _27592_ (.A(_03809_),
    .B(_03803_),
    .X(_03837_));
 sky130_fd_sc_hd__nand2_1 _27593_ (.A(_03837_),
    .B(_03404_),
    .Y(_03838_));
 sky130_fd_sc_hd__nand2_1 _27594_ (.A(_03805_),
    .B(net239),
    .Y(_03840_));
 sky130_fd_sc_hd__nand2_1 _27595_ (.A(_03838_),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__inv_2 _27596_ (.A(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__nand2_1 _27597_ (.A(_03842_),
    .B(_11840_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _27598_ (.A(_03841_),
    .B(_11838_),
    .Y(_03844_));
 sky130_fd_sc_hd__nand2_1 _27599_ (.A(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__inv_4 _27600_ (.A(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__nand2_1 _27601_ (.A(_03836_),
    .B(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__nand2_1 _27602_ (.A(_03847_),
    .B(_03843_),
    .Y(_03848_));
 sky130_fd_sc_hd__or2_1 _27603_ (.A(_03830_),
    .B(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_1 _27604_ (.A(_03848_),
    .B(_03830_),
    .Y(_03851_));
 sky130_fd_sc_hd__nand2_1 _27605_ (.A(_03849_),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__nand2_1 _27606_ (.A(_03852_),
    .B(_12914_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand3_1 _27607_ (.A(_03849_),
    .B(_11774_),
    .C(_03851_),
    .Y(_03854_));
 sky130_fd_sc_hd__nand2_1 _27608_ (.A(_03853_),
    .B(_03854_),
    .Y(_03855_));
 sky130_fd_sc_hd__inv_2 _27609_ (.A(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__or2_1 _27610_ (.A(_03846_),
    .B(_03836_),
    .X(_03857_));
 sky130_fd_sc_hd__nand2_1 _27611_ (.A(_03857_),
    .B(_03847_),
    .Y(_03858_));
 sky130_fd_sc_hd__nor2_1 _27612_ (.A(_13461_),
    .B(_03858_),
    .Y(_03859_));
 sky130_fd_sc_hd__inv_2 _27613_ (.A(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__nand2_1 _27614_ (.A(_03858_),
    .B(_13461_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _27615_ (.A(_03860_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__clkinvlp_2 _27616_ (.A(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__nand3_2 _27617_ (.A(_03802_),
    .B(_03856_),
    .C(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__a21bo_1 _27618_ (.A1(_01922_),
    .A2(_02011_),
    .B1_N(_02012_),
    .X(_03866_));
 sky130_fd_sc_hd__xor2_1 _27619_ (.A(_02004_),
    .B(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__or2_1 _27620_ (.A(_12914_),
    .B(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__nand2_1 _27621_ (.A(_03867_),
    .B(_12914_),
    .Y(_03869_));
 sky130_fd_sc_hd__nand2_1 _27622_ (.A(_03868_),
    .B(_03869_),
    .Y(_03870_));
 sky130_fd_sc_hd__a21o_1 _27623_ (.A1(_03820_),
    .A2(_03815_),
    .B1(_03870_),
    .X(_03871_));
 sky130_fd_sc_hd__nand3_1 _27624_ (.A(_03820_),
    .B(_03815_),
    .C(_03870_),
    .Y(_03873_));
 sky130_fd_sc_hd__nand2_1 _27625_ (.A(_03871_),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nand2_1 _27626_ (.A(_03874_),
    .B(_03746_),
    .Y(_03875_));
 sky130_fd_sc_hd__nand2_1 _27627_ (.A(\div1i.quot[0] ),
    .B(_03867_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _27628_ (.A(_03875_),
    .B(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _27629_ (.A(_03877_),
    .B(_13537_),
    .Y(_03878_));
 sky130_fd_sc_hd__nand3_2 _27630_ (.A(_03875_),
    .B(_07400_),
    .C(_03876_),
    .Y(_03879_));
 sky130_fd_sc_hd__nand2_1 _27631_ (.A(_03878_),
    .B(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hd__inv_2 _27632_ (.A(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__nand3_2 _27633_ (.A(_03836_),
    .B(_03830_),
    .C(_03846_),
    .Y(_03882_));
 sky130_fd_sc_hd__inv_2 _27634_ (.A(_03843_),
    .Y(_03884_));
 sky130_fd_sc_hd__a21boi_1 _27635_ (.A1(_03884_),
    .A2(_03826_),
    .B1_N(_03827_),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _27636_ (.A(_03882_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand2_2 _27637_ (.A(_03881_),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__nand3_1 _27638_ (.A(_03880_),
    .B(_03882_),
    .C(_03885_),
    .Y(_03888_));
 sky130_fd_sc_hd__nand2_1 _27639_ (.A(_03887_),
    .B(_03888_),
    .Y(_03889_));
 sky130_fd_sc_hd__nand2_1 _27640_ (.A(_03889_),
    .B(_12939_),
    .Y(_03890_));
 sky130_fd_sc_hd__nand3_1 _27641_ (.A(_03887_),
    .B(_03888_),
    .C(_11797_),
    .Y(_03891_));
 sky130_fd_sc_hd__nand2_1 _27642_ (.A(_03890_),
    .B(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__inv_2 _27643_ (.A(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__a21boi_2 _27644_ (.A1(_03853_),
    .A2(_03859_),
    .B1_N(_03854_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand3_1 _27645_ (.A(_03865_),
    .B(_03893_),
    .C(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__nand2_1 _27646_ (.A(_03802_),
    .B(_03864_),
    .Y(_03897_));
 sky130_fd_sc_hd__nand2_1 _27647_ (.A(_03897_),
    .B(_03860_),
    .Y(_03898_));
 sky130_fd_sc_hd__nand2_1 _27648_ (.A(_03898_),
    .B(_03855_),
    .Y(_03899_));
 sky130_fd_sc_hd__nand2_1 _27649_ (.A(_03896_),
    .B(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__nand2_1 _27650_ (.A(_03887_),
    .B(_03879_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _27651_ (.A(_03868_),
    .B(_03815_),
    .Y(_03902_));
 sky130_fd_sc_hd__inv_2 _27652_ (.A(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__nand2_2 _27653_ (.A(_03820_),
    .B(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__nand2_1 _27654_ (.A(_03904_),
    .B(_03869_),
    .Y(_03906_));
 sky130_fd_sc_hd__a21o_1 _27655_ (.A1(_01922_),
    .A2(_02015_),
    .B1(_02017_),
    .X(_03907_));
 sky130_fd_sc_hd__xor2_1 _27656_ (.A(_01995_),
    .B(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__or2_1 _27657_ (.A(_12939_),
    .B(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__nand2_1 _27658_ (.A(_03908_),
    .B(_12939_),
    .Y(_03910_));
 sky130_fd_sc_hd__nand2_1 _27659_ (.A(_03909_),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__nand2_1 _27660_ (.A(_03906_),
    .B(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__inv_2 _27661_ (.A(_03911_),
    .Y(_03913_));
 sky130_fd_sc_hd__nand3_2 _27662_ (.A(_03904_),
    .B(_03913_),
    .C(_03869_),
    .Y(_03914_));
 sky130_fd_sc_hd__nand2_1 _27663_ (.A(_03912_),
    .B(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__nand2_1 _27664_ (.A(_03915_),
    .B(_03746_),
    .Y(_03917_));
 sky130_fd_sc_hd__nand2_1 _27665_ (.A(\div1i.quot[0] ),
    .B(_03908_),
    .Y(_03918_));
 sky130_fd_sc_hd__nand2_1 _27666_ (.A(_03917_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__nand2_1 _27667_ (.A(_03919_),
    .B(_11811_),
    .Y(_03920_));
 sky130_fd_sc_hd__nand3_1 _27668_ (.A(_03917_),
    .B(_11808_),
    .C(_03918_),
    .Y(_03921_));
 sky130_fd_sc_hd__nand2_1 _27669_ (.A(_03920_),
    .B(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__inv_2 _27670_ (.A(_03922_),
    .Y(_03923_));
 sky130_fd_sc_hd__nand2_1 _27671_ (.A(_03901_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__nand3_1 _27672_ (.A(_03887_),
    .B(_03922_),
    .C(_03879_),
    .Y(_03925_));
 sky130_fd_sc_hd__nand2_1 _27673_ (.A(_03924_),
    .B(_03925_),
    .Y(_03926_));
 sky130_fd_sc_hd__nand2_2 _27674_ (.A(_03926_),
    .B(_12992_),
    .Y(_03928_));
 sky130_fd_sc_hd__nand3_2 _27675_ (.A(_03924_),
    .B(_11858_),
    .C(_03925_),
    .Y(_03929_));
 sky130_fd_sc_hd__nand2_1 _27676_ (.A(_03928_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__and2_1 _27677_ (.A(_03930_),
    .B(_03890_),
    .X(_03931_));
 sky130_fd_sc_hd__and2_1 _27678_ (.A(_03725_),
    .B(_03687_),
    .X(_03932_));
 sky130_fd_sc_hd__or2_1 _27679_ (.A(_03488_),
    .B(_03479_),
    .X(_03933_));
 sky130_fd_sc_hd__nand2_1 _27680_ (.A(_03933_),
    .B(_03489_),
    .Y(_03934_));
 sky130_fd_sc_hd__nand2_1 _27681_ (.A(_03467_),
    .B(_03477_),
    .Y(_03935_));
 sky130_fd_sc_hd__xor2_1 _27682_ (.A(_03475_),
    .B(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__nand2_1 _27683_ (.A(_03471_),
    .B(_03473_),
    .Y(_03937_));
 sky130_fd_sc_hd__xor2_1 _27684_ (.A(_03472_),
    .B(_03937_),
    .X(_03939_));
 sky130_fd_sc_hd__and3_1 _27685_ (.A(_03934_),
    .B(_03936_),
    .C(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__nand2_1 _27686_ (.A(_03500_),
    .B(_03461_),
    .Y(_03941_));
 sky130_fd_sc_hd__nand3_1 _27687_ (.A(_03497_),
    .B(_03499_),
    .C(_03460_),
    .Y(_03942_));
 sky130_fd_sc_hd__nand2_1 _27688_ (.A(_03941_),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__nand2_1 _27689_ (.A(_03496_),
    .B(_03499_),
    .Y(_03944_));
 sky130_fd_sc_hd__xor2_1 _27690_ (.A(_03490_),
    .B(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__nand3_1 _27691_ (.A(_03940_),
    .B(_03943_),
    .C(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__nor2_1 _27692_ (.A(_03932_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _27693_ (.A(_03453_),
    .B(_03455_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _27694_ (.A(_03941_),
    .B(_03459_),
    .Y(_03950_));
 sky130_fd_sc_hd__xor2_1 _27695_ (.A(_03948_),
    .B(_03950_),
    .X(_03951_));
 sky130_fd_sc_hd__nand2_1 _27696_ (.A(_03504_),
    .B(_03563_),
    .Y(_03952_));
 sky130_fd_sc_hd__nand3_1 _27697_ (.A(_03501_),
    .B(_03503_),
    .C(_03562_),
    .Y(_03953_));
 sky130_fd_sc_hd__nand2_1 _27698_ (.A(_03952_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hd__nand3_1 _27699_ (.A(_03947_),
    .B(_03951_),
    .C(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__nand2_1 _27700_ (.A(_03571_),
    .B(_03645_),
    .Y(_03956_));
 sky130_fd_sc_hd__nand3_1 _27701_ (.A(_03568_),
    .B(_03570_),
    .C(_03644_),
    .Y(_03957_));
 sky130_fd_sc_hd__nand2_1 _27702_ (.A(_03956_),
    .B(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__inv_2 _27703_ (.A(_03958_),
    .Y(_03959_));
 sky130_fd_sc_hd__nor2_2 _27704_ (.A(_03955_),
    .B(_03959_),
    .Y(_03961_));
 sky130_fd_sc_hd__nand2_1 _27705_ (.A(_03783_),
    .B(_03791_),
    .Y(_03962_));
 sky130_fd_sc_hd__a21o_1 _27706_ (.A1(_03727_),
    .A2(_03799_),
    .B1(_03962_),
    .X(_03963_));
 sky130_fd_sc_hd__nand2_1 _27707_ (.A(_03963_),
    .B(_03790_),
    .Y(_03964_));
 sky130_fd_sc_hd__nand2_1 _27708_ (.A(_03557_),
    .B(_03565_),
    .Y(_03965_));
 sky130_fd_sc_hd__nand2_1 _27709_ (.A(_03952_),
    .B(_03561_),
    .Y(_03966_));
 sky130_fd_sc_hd__xor2_1 _27710_ (.A(_03965_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__nand3_2 _27711_ (.A(_03961_),
    .B(_03964_),
    .C(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hd__nor2_1 _27712_ (.A(_03931_),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__o21ai_1 _27713_ (.A1(_03859_),
    .A2(_03855_),
    .B1(_03863_),
    .Y(_03970_));
 sky130_fd_sc_hd__o21ai_1 _27714_ (.A1(_03970_),
    .A2(_03802_),
    .B1(_03897_),
    .Y(_03972_));
 sky130_fd_sc_hd__nand2_1 _27715_ (.A(_03726_),
    .B(_03686_),
    .Y(_03973_));
 sky130_fd_sc_hd__nand3_1 _27716_ (.A(_03648_),
    .B(_03650_),
    .C(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__nand2_1 _27717_ (.A(_03974_),
    .B(_03688_),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_1 _27718_ (.A(_03962_),
    .B(_03788_),
    .Y(_03976_));
 sky130_fd_sc_hd__nand2_1 _27719_ (.A(_03976_),
    .B(_03797_),
    .Y(_03977_));
 sky130_fd_sc_hd__nand2_1 _27720_ (.A(_03977_),
    .B(_03799_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2_1 _27721_ (.A(_03978_),
    .B(_03789_),
    .Y(_03979_));
 sky130_fd_sc_hd__nand2_1 _27722_ (.A(_03975_),
    .B(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hd__or2_1 _27723_ (.A(_03790_),
    .B(_03727_),
    .X(_03981_));
 sky130_fd_sc_hd__nand2_1 _27724_ (.A(_03651_),
    .B(_03981_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2_1 _27725_ (.A(_03983_),
    .B(_03689_),
    .Y(_03984_));
 sky130_fd_sc_hd__nand2_1 _27726_ (.A(_03956_),
    .B(_03643_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _27727_ (.A(_03634_),
    .B(_03638_),
    .Y(_03986_));
 sky130_fd_sc_hd__inv_2 _27728_ (.A(_03986_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand2_1 _27729_ (.A(_03985_),
    .B(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__nand3_1 _27730_ (.A(_03956_),
    .B(_03986_),
    .C(_03643_),
    .Y(_03989_));
 sky130_fd_sc_hd__nand2_1 _27731_ (.A(_03988_),
    .B(_03989_),
    .Y(_03990_));
 sky130_fd_sc_hd__nand2_1 _27732_ (.A(_03984_),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hd__nor2_2 _27733_ (.A(_03980_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__nand3_1 _27734_ (.A(_03969_),
    .B(_03972_),
    .C(_03992_),
    .Y(_03994_));
 sky130_fd_sc_hd__nor2_1 _27735_ (.A(_03900_),
    .B(_03994_),
    .Y(_03995_));
 sky130_fd_sc_hd__inv_2 _27736_ (.A(_03891_),
    .Y(_03996_));
 sky130_fd_sc_hd__o21ai_1 _27737_ (.A1(_03996_),
    .A2(_03930_),
    .B1(_03895_),
    .Y(_03997_));
 sky130_fd_sc_hd__inv_2 _27738_ (.A(_03865_),
    .Y(_03998_));
 sky130_fd_sc_hd__o21ai_1 _27739_ (.A1(_03997_),
    .A2(_03998_),
    .B1(_03892_),
    .Y(_03999_));
 sky130_fd_sc_hd__nand2_2 _27740_ (.A(_03995_),
    .B(_03999_),
    .Y(_04000_));
 sky130_fd_sc_hd__nand3_1 _27741_ (.A(_03923_),
    .B(_03881_),
    .C(_03886_),
    .Y(_04001_));
 sky130_fd_sc_hd__clkinvlp_2 _27742_ (.A(_03879_),
    .Y(_04002_));
 sky130_fd_sc_hd__a21boi_1 _27743_ (.A1(_04002_),
    .A2(_03920_),
    .B1_N(_03921_),
    .Y(_04003_));
 sky130_fd_sc_hd__nand2_2 _27744_ (.A(_04001_),
    .B(_04003_),
    .Y(_04005_));
 sky130_fd_sc_hd__a21bo_1 _27745_ (.A1(_03907_),
    .A2(_01993_),
    .B1_N(_01994_),
    .X(_04006_));
 sky130_fd_sc_hd__xor2_1 _27746_ (.A(_01984_),
    .B(_04006_),
    .X(_04007_));
 sky130_fd_sc_hd__or2_1 _27747_ (.A(_12992_),
    .B(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__nand2_1 _27748_ (.A(_04007_),
    .B(_12992_),
    .Y(_04009_));
 sky130_fd_sc_hd__nand2_1 _27749_ (.A(_04008_),
    .B(_04009_),
    .Y(_04010_));
 sky130_fd_sc_hd__nand2_1 _27750_ (.A(_03914_),
    .B(_03909_),
    .Y(_04011_));
 sky130_fd_sc_hd__xor2_1 _27751_ (.A(_04010_),
    .B(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__nand2_1 _27752_ (.A(_04012_),
    .B(_03746_),
    .Y(_04013_));
 sky130_fd_sc_hd__nand2_1 _27753_ (.A(_04007_),
    .B(\div1i.quot[0] ),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_1 _27754_ (.A(_04013_),
    .B(_04014_),
    .Y(_04016_));
 sky130_fd_sc_hd__nand2_1 _27755_ (.A(_04016_),
    .B(_11896_),
    .Y(_04017_));
 sky130_fd_sc_hd__nand3_2 _27756_ (.A(_04013_),
    .B(_11899_),
    .C(_04014_),
    .Y(_04018_));
 sky130_fd_sc_hd__nand2_1 _27757_ (.A(_04017_),
    .B(_04018_),
    .Y(_04019_));
 sky130_fd_sc_hd__inv_2 _27758_ (.A(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__nand2_1 _27759_ (.A(_04008_),
    .B(_03909_),
    .Y(_04021_));
 sky130_fd_sc_hd__inv_2 _27760_ (.A(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__nand2_2 _27761_ (.A(_03914_),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hd__nand2_1 _27762_ (.A(_04023_),
    .B(_04009_),
    .Y(_04024_));
 sky130_fd_sc_hd__nand2_1 _27763_ (.A(_02065_),
    .B(_02066_),
    .Y(_04025_));
 sky130_fd_sc_hd__xor2_1 _27764_ (.A(_04025_),
    .B(_02020_),
    .X(_04027_));
 sky130_fd_sc_hd__or2_1 _27765_ (.A(_14113_),
    .B(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__nand2_1 _27766_ (.A(_04027_),
    .B(_14113_),
    .Y(_04029_));
 sky130_fd_sc_hd__nand2_1 _27767_ (.A(_04028_),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_1 _27768_ (.A(_04024_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__inv_2 _27769_ (.A(_04030_),
    .Y(_04032_));
 sky130_fd_sc_hd__nand3_2 _27770_ (.A(_04023_),
    .B(_04032_),
    .C(_04009_),
    .Y(_04033_));
 sky130_fd_sc_hd__nand2_1 _27771_ (.A(_04031_),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__nand2_1 _27772_ (.A(_04034_),
    .B(_03746_),
    .Y(_04035_));
 sky130_fd_sc_hd__nand2_1 _27773_ (.A(\div1i.quot[0] ),
    .B(_04027_),
    .Y(_04036_));
 sky130_fd_sc_hd__nand2_1 _27774_ (.A(_04035_),
    .B(_04036_),
    .Y(_04038_));
 sky130_fd_sc_hd__nand2_1 _27775_ (.A(_04038_),
    .B(_08020_),
    .Y(_04039_));
 sky130_fd_sc_hd__nand3_1 _27776_ (.A(_04035_),
    .B(_13022_),
    .C(_04036_),
    .Y(_04040_));
 sky130_fd_sc_hd__nand2_1 _27777_ (.A(_04039_),
    .B(_04040_),
    .Y(_04041_));
 sky130_fd_sc_hd__inv_2 _27778_ (.A(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__nand3_1 _27779_ (.A(_04005_),
    .B(_04020_),
    .C(_04042_),
    .Y(_04043_));
 sky130_fd_sc_hd__clkinvlp_2 _27780_ (.A(_04018_),
    .Y(_04044_));
 sky130_fd_sc_hd__a21boi_1 _27781_ (.A1(_04044_),
    .A2(_04039_),
    .B1_N(_04040_),
    .Y(_04045_));
 sky130_fd_sc_hd__nand2_1 _27782_ (.A(_04043_),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_1 _27783_ (.A(_04033_),
    .B(_04028_),
    .Y(_04047_));
 sky130_fd_sc_hd__a21bo_1 _27784_ (.A1(_02020_),
    .A2(_02065_),
    .B1_N(_02066_),
    .X(_04049_));
 sky130_fd_sc_hd__xor2_1 _27785_ (.A(_02056_),
    .B(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__or2_1 _27786_ (.A(_13042_),
    .B(_04050_),
    .X(_04051_));
 sky130_fd_sc_hd__nand2_1 _27787_ (.A(_04050_),
    .B(_13042_),
    .Y(_04052_));
 sky130_fd_sc_hd__nand2_1 _27788_ (.A(_04051_),
    .B(_04052_),
    .Y(_04053_));
 sky130_fd_sc_hd__nand2_1 _27789_ (.A(_04047_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__nand3b_1 _27790_ (.A_N(_04053_),
    .B(_04033_),
    .C(_04028_),
    .Y(_04055_));
 sky130_fd_sc_hd__nand3_1 _27791_ (.A(_04054_),
    .B(_04055_),
    .C(_03746_),
    .Y(_04056_));
 sky130_fd_sc_hd__nand2_1 _27792_ (.A(_04050_),
    .B(\div1i.quot[0] ),
    .Y(_04057_));
 sky130_fd_sc_hd__nand2_1 _27793_ (.A(_04056_),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__or2_1 _27794_ (.A(_12506_),
    .B(_04058_),
    .X(_04060_));
 sky130_fd_sc_hd__nand2_1 _27795_ (.A(_04058_),
    .B(_12506_),
    .Y(_04061_));
 sky130_fd_sc_hd__nand2_1 _27796_ (.A(_04060_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hd__inv_2 _27797_ (.A(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2_1 _27798_ (.A(_04046_),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__nand2_1 _27799_ (.A(_04064_),
    .B(_04060_),
    .Y(_04065_));
 sky130_fd_sc_hd__nand2_1 _27800_ (.A(_04047_),
    .B(_04052_),
    .Y(_04066_));
 sky130_fd_sc_hd__a21oi_1 _27801_ (.A1(_02016_),
    .A2(_02019_),
    .B1(_02067_),
    .Y(_04067_));
 sky130_fd_sc_hd__or2_1 _27802_ (.A(_02120_),
    .B(_04067_),
    .X(_04068_));
 sky130_fd_sc_hd__or2_1 _27803_ (.A(_02088_),
    .B(_04068_),
    .X(_04069_));
 sky130_fd_sc_hd__nand2_1 _27804_ (.A(_04068_),
    .B(_02088_),
    .Y(_04071_));
 sky130_fd_sc_hd__nand2_1 _27805_ (.A(_04069_),
    .B(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__or2_1 _27806_ (.A(_13633_),
    .B(_04072_),
    .X(_04073_));
 sky130_fd_sc_hd__nand2_1 _27807_ (.A(_04072_),
    .B(_13633_),
    .Y(_04074_));
 sky130_fd_sc_hd__nand2_1 _27808_ (.A(_04073_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__a21o_1 _27809_ (.A1(_04066_),
    .A2(_04051_),
    .B1(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__nand3_1 _27810_ (.A(_04066_),
    .B(_04051_),
    .C(_04075_),
    .Y(_04077_));
 sky130_fd_sc_hd__nand2_1 _27811_ (.A(_04076_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__nand2_1 _27812_ (.A(_04078_),
    .B(_03746_),
    .Y(_04079_));
 sky130_fd_sc_hd__nand2_1 _27813_ (.A(_04072_),
    .B(\div1i.quot[0] ),
    .Y(_04080_));
 sky130_fd_sc_hd__nand2_1 _27814_ (.A(_04079_),
    .B(_04080_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand2_1 _27815_ (.A(_04082_),
    .B(_11948_),
    .Y(_04083_));
 sky130_fd_sc_hd__nand3_1 _27816_ (.A(_04079_),
    .B(_11946_),
    .C(_04080_),
    .Y(_04084_));
 sky130_fd_sc_hd__nand2_1 _27817_ (.A(_04083_),
    .B(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__inv_2 _27818_ (.A(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__nand2_1 _27819_ (.A(_04065_),
    .B(_04086_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand2_1 _27820_ (.A(_04087_),
    .B(_04084_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand2_1 _27821_ (.A(_04071_),
    .B(_02086_),
    .Y(_04089_));
 sky130_fd_sc_hd__xor2_1 _27822_ (.A(_02114_),
    .B(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__nand3_1 _27823_ (.A(_04076_),
    .B(_03746_),
    .C(_04073_),
    .Y(_04091_));
 sky130_fd_sc_hd__xor2_1 _27824_ (.A(_04090_),
    .B(_04091_),
    .X(_04093_));
 sky130_fd_sc_hd__inv_2 _27825_ (.A(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__nand2b_2 _27826_ (.A_N(_04088_),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__nand2_2 _27827_ (.A(_04088_),
    .B(_04093_),
    .Y(_04096_));
 sky130_fd_sc_hd__nand2_2 _27828_ (.A(_04095_),
    .B(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__nand2b_1 _27829_ (.A_N(_04005_),
    .B(_04019_),
    .Y(_04098_));
 sky130_fd_sc_hd__nand2_2 _27830_ (.A(_04005_),
    .B(_04020_),
    .Y(_04099_));
 sky130_fd_sc_hd__nand2_1 _27831_ (.A(_04098_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__inv_2 _27832_ (.A(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hd__inv_2 _27833_ (.A(_03852_),
    .Y(_04102_));
 sky130_fd_sc_hd__nand3_1 _27834_ (.A(_03683_),
    .B(_03556_),
    .C(_03639_),
    .Y(_04104_));
 sky130_fd_sc_hd__and4_1 _27835_ (.A(_03483_),
    .B(_03466_),
    .C(_05167_),
    .D(_03470_),
    .X(_04105_));
 sky130_fd_sc_hd__and3_1 _27836_ (.A(_04105_),
    .B(_03495_),
    .C(_03457_),
    .X(_04106_));
 sky130_fd_sc_hd__nand3_1 _27837_ (.A(_04106_),
    .B(_03452_),
    .C(_03558_),
    .Y(_04107_));
 sky130_fd_sc_hd__nor2_1 _27838_ (.A(_04104_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__nand2_1 _27839_ (.A(_04108_),
    .B(_03858_),
    .Y(_04109_));
 sky130_fd_sc_hd__inv_2 _27840_ (.A(_04109_),
    .Y(_04110_));
 sky130_fd_sc_hd__and3_1 _27841_ (.A(_03633_),
    .B(_03786_),
    .C(_03722_),
    .X(_04111_));
 sky130_fd_sc_hd__nand3_1 _27842_ (.A(_04110_),
    .B(_04111_),
    .C(_03782_),
    .Y(_04112_));
 sky130_fd_sc_hd__nor2_1 _27843_ (.A(_04102_),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__nand3_1 _27844_ (.A(_04113_),
    .B(_03889_),
    .C(_03926_),
    .Y(_04115_));
 sky130_fd_sc_hd__nor2_1 _27845_ (.A(_04101_),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__nand3_1 _27846_ (.A(_04062_),
    .B(_04043_),
    .C(_04045_),
    .Y(_04117_));
 sky130_fd_sc_hd__nand2_1 _27847_ (.A(_04064_),
    .B(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__nand2_1 _27848_ (.A(_04099_),
    .B(_04018_),
    .Y(_04119_));
 sky130_fd_sc_hd__nand2_1 _27849_ (.A(_04119_),
    .B(_04042_),
    .Y(_04120_));
 sky130_fd_sc_hd__nand3_1 _27850_ (.A(_04099_),
    .B(_04041_),
    .C(_04018_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_1 _27851_ (.A(_04120_),
    .B(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__nand3_1 _27852_ (.A(_04116_),
    .B(_04118_),
    .C(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand3_1 _27853_ (.A(_04095_),
    .B(_04096_),
    .C(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__nand2_2 _27854_ (.A(\div1i.quot[0] ),
    .B(_12221_),
    .Y(_04126_));
 sky130_fd_sc_hd__nand2_1 _27855_ (.A(_04124_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__a21oi_4 _27856_ (.A1(_04000_),
    .A2(_04097_),
    .B1(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__or2_1 _27857_ (.A(_13633_),
    .B(_04118_),
    .X(_04129_));
 sky130_fd_sc_hd__a21boi_1 _27858_ (.A1(_04095_),
    .A2(_04096_),
    .B1_N(_04129_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand3_2 _27859_ (.A(_03928_),
    .B(_03893_),
    .C(_03929_),
    .Y(_04131_));
 sky130_fd_sc_hd__inv_2 _27860_ (.A(_03929_),
    .Y(_04132_));
 sky130_fd_sc_hd__a21o_1 _27861_ (.A1(_03928_),
    .A2(_03996_),
    .B1(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__nor2_1 _27862_ (.A(_03895_),
    .B(_04131_),
    .Y(_04134_));
 sky130_fd_sc_hd__nor2_2 _27863_ (.A(_04133_),
    .B(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hd__o21ai_1 _27864_ (.A1(_04131_),
    .A2(_03865_),
    .B1(_04135_),
    .Y(_04137_));
 sky130_fd_sc_hd__nand2_1 _27865_ (.A(_04100_),
    .B(_14113_),
    .Y(_04138_));
 sky130_fd_sc_hd__nand3_1 _27866_ (.A(_04098_),
    .B(_08554_),
    .C(_04099_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _27867_ (.A(_04138_),
    .B(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__inv_2 _27868_ (.A(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_1 _27869_ (.A(_04122_),
    .B(_13042_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand3_2 _27870_ (.A(_04120_),
    .B(_12495_),
    .C(_04121_),
    .Y(_04143_));
 sky130_fd_sc_hd__nand3_1 _27871_ (.A(_04141_),
    .B(_04142_),
    .C(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__inv_2 _27872_ (.A(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2_1 _27873_ (.A(_04137_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__nand2_1 _27874_ (.A(_04142_),
    .B(_04143_),
    .Y(_04148_));
 sky130_fd_sc_hd__o21a_1 _27875_ (.A1(_04139_),
    .A2(_04148_),
    .B1(_04143_),
    .X(_04149_));
 sky130_fd_sc_hd__nand2_1 _27876_ (.A(_04146_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__nand2_1 _27877_ (.A(_04118_),
    .B(_13633_),
    .Y(_04151_));
 sky130_fd_sc_hd__nand2_1 _27878_ (.A(_04150_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__nand2_1 _27879_ (.A(_04130_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__nand3_1 _27880_ (.A(_04064_),
    .B(_04085_),
    .C(_04060_),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _27881_ (.A(_04087_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__inv_2 _27882_ (.A(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__nand2_2 _27883_ (.A(_04153_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__nand2_4 _27884_ (.A(_04128_),
    .B(_04157_),
    .Y(_04159_));
 sky130_fd_sc_hd__inv_2 _27885_ (.A(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__nand2_1 _27886_ (.A(_02304_),
    .B(net167),
    .Y(_04161_));
 sky130_fd_sc_hd__nand2_1 _27887_ (.A(_04129_),
    .B(_04151_),
    .Y(_04162_));
 sky130_fd_sc_hd__inv_2 _27888_ (.A(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__nand2_1 _27889_ (.A(_04150_),
    .B(_04163_),
    .Y(_04164_));
 sky130_fd_sc_hd__o21ai_1 _27890_ (.A1(_04151_),
    .A2(_04155_),
    .B1(_04129_),
    .Y(_04165_));
 sky130_fd_sc_hd__nand3_1 _27891_ (.A(_04146_),
    .B(_04165_),
    .C(_04149_),
    .Y(_04166_));
 sky130_fd_sc_hd__nand2_2 _27892_ (.A(_04164_),
    .B(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__inv_2 _27893_ (.A(_04131_),
    .Y(_04168_));
 sky130_fd_sc_hd__nand2_1 _27894_ (.A(_03998_),
    .B(_04168_),
    .Y(_04170_));
 sky130_fd_sc_hd__nand3_1 _27895_ (.A(_04170_),
    .B(_04135_),
    .C(_04141_),
    .Y(_04171_));
 sky130_fd_sc_hd__nand2_1 _27896_ (.A(_04148_),
    .B(_04138_),
    .Y(_04172_));
 sky130_fd_sc_hd__nand2_1 _27897_ (.A(_04171_),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__nand3_1 _27898_ (.A(_04142_),
    .B(_04143_),
    .C(_04139_),
    .Y(_04174_));
 sky130_fd_sc_hd__nand3_1 _27899_ (.A(_04170_),
    .B(_04135_),
    .C(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nand2_1 _27900_ (.A(_04175_),
    .B(_04140_),
    .Y(_04176_));
 sky130_fd_sc_hd__inv_2 _27901_ (.A(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__nor2_2 _27902_ (.A(_04173_),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hd__nand2_1 _27903_ (.A(_04167_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__nand2_2 _27904_ (.A(_04179_),
    .B(_04097_),
    .Y(_04181_));
 sky130_fd_sc_hd__nand3_2 _27905_ (.A(_04160_),
    .B(net168),
    .C(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__buf_6 _27906_ (.A(_04182_),
    .X(_04183_));
 sky130_fd_sc_hd__inv_2 _27907_ (.A(net67),
    .Y(_04184_));
 sky130_fd_sc_hd__and3_1 _27908_ (.A(_04184_),
    .B(net66),
    .C(net65),
    .X(_04185_));
 sky130_fd_sc_hd__inv_2 _27909_ (.A(net65),
    .Y(_04186_));
 sky130_fd_sc_hd__and3_1 _27910_ (.A(_04184_),
    .B(_04186_),
    .C(net66),
    .X(_04187_));
 sky130_fd_sc_hd__mux2_4 _27911_ (.A0(_04185_),
    .A1(_04187_),
    .S(net107),
    .X(_04188_));
 sky130_fd_sc_hd__clkinvlp_2 _27912_ (.A(_04188_),
    .Y(_04189_));
 sky130_fd_sc_hd__or3_1 _27913_ (.A(net66),
    .B(net65),
    .C(_04184_),
    .X(_04190_));
 sky130_fd_sc_hd__nor2_4 _27914_ (.A(net168),
    .B(_04190_),
    .Y(_04192_));
 sky130_fd_sc_hd__inv_2 _27915_ (.A(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__buf_6 _27916_ (.A(_04193_),
    .X(_04194_));
 sky130_fd_sc_hd__nand2_1 _27917_ (.A(_04189_),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _27918_ (.A(_04183_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__clkinvlp_2 _27919_ (.A(net189),
    .Y(_04197_));
 sky130_fd_sc_hd__nor2_1 _27920_ (.A(_02203_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__and2_1 _27921_ (.A(_04196_),
    .B(net190),
    .X(_04199_));
 sky130_fd_sc_hd__inv_2 _27922_ (.A(net66),
    .Y(_04200_));
 sky130_fd_sc_hd__and3_1 _27923_ (.A(_04184_),
    .B(_04200_),
    .C(net65),
    .X(_04201_));
 sky130_fd_sc_hd__buf_6 _27924_ (.A(_04201_),
    .X(_04203_));
 sky130_fd_sc_hd__inv_4 _27925_ (.A(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__buf_6 _27926_ (.A(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__o21ai_1 _27927_ (.A1(net190),
    .A2(_04196_),
    .B1(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__nand3_4 _27928_ (.A(_04181_),
    .B(_04157_),
    .C(_04128_),
    .Y(_04207_));
 sky130_fd_sc_hd__inv_2 _27929_ (.A(net190),
    .Y(_04208_));
 sky130_fd_sc_hd__inv_2 _27930_ (.A(net168),
    .Y(_04209_));
 sky130_fd_sc_hd__buf_6 _27931_ (.A(_04209_),
    .X(_04210_));
 sky130_fd_sc_hd__buf_6 _27932_ (.A(_04210_),
    .X(_04211_));
 sky130_fd_sc_hd__buf_6 _27933_ (.A(_04204_),
    .X(_04212_));
 sky130_fd_sc_hd__a31o_1 _27934_ (.A1(_02519_),
    .A2(_02162_),
    .A3(net168),
    .B1(_04212_),
    .X(_04214_));
 sky130_fd_sc_hd__a31o_1 _27935_ (.A1(_04207_),
    .A2(_04208_),
    .A3(_04211_),
    .B1(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__o21ai_1 _27936_ (.A1(_04199_),
    .A2(_04206_),
    .B1(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__and3_1 _27937_ (.A(_04184_),
    .B(_04200_),
    .C(_04186_),
    .X(_04217_));
 sky130_fd_sc_hd__and2b_1 _27938_ (.A_N(net107),
    .B(_04187_),
    .X(_04218_));
 sky130_fd_sc_hd__nand2_1 _27939_ (.A(_04185_),
    .B(net107),
    .Y(_04219_));
 sky130_fd_sc_hd__or3b_1 _27940_ (.A(_04217_),
    .B(_04218_),
    .C_N(_04219_),
    .X(_04220_));
 sky130_fd_sc_hd__buf_6 _27941_ (.A(_04220_),
    .X(_04221_));
 sky130_fd_sc_hd__buf_6 _27942_ (.A(_04221_),
    .X(_04222_));
 sky130_fd_sc_hd__mux2_1 _27943_ (.A0(_04216_),
    .A1(_04208_),
    .S(_04222_),
    .X(_04223_));
 sky130_fd_sc_hd__or2_1 _27944_ (.A(_02652_),
    .B(_04223_),
    .X(_04225_));
 sky130_fd_sc_hd__inv_2 _27945_ (.A(_04225_),
    .Y(_00003_));
 sky130_fd_sc_hd__inv_2 _27946_ (.A(net173),
    .Y(_04226_));
 sky130_fd_sc_hd__nor2_1 _27947_ (.A(_02152_),
    .B(net174),
    .Y(_04227_));
 sky130_fd_sc_hd__clkinvlp_2 _27948_ (.A(net175),
    .Y(_04228_));
 sky130_fd_sc_hd__nand2_1 _27949_ (.A(_04228_),
    .B(_04208_),
    .Y(_04229_));
 sky130_fd_sc_hd__nand2_1 _27950_ (.A(net175),
    .B(net190),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_1 _27951_ (.A(_04229_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__clkinvlp_2 _27952_ (.A(_04231_),
    .Y(_04232_));
 sky130_fd_sc_hd__nand2_1 _27953_ (.A(_04183_),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__a21boi_4 _27954_ (.A1(_04167_),
    .A2(_04178_),
    .B1_N(_04097_),
    .Y(_04235_));
 sky130_fd_sc_hd__nor2_8 _27955_ (.A(_04159_),
    .B(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hd__buf_6 _27956_ (.A(_04236_),
    .X(_04237_));
 sky130_fd_sc_hd__buf_6 _27957_ (.A(net168),
    .X(_04238_));
 sky130_fd_sc_hd__nand3_1 _27958_ (.A(net131),
    .B(_04238_),
    .C(net175),
    .Y(_04239_));
 sky130_fd_sc_hd__buf_6 _27959_ (.A(_04188_),
    .X(_04240_));
 sky130_fd_sc_hd__nand3_1 _27960_ (.A(_04233_),
    .B(_04239_),
    .C(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__buf_6 _27961_ (.A(_04193_),
    .X(_04242_));
 sky130_fd_sc_hd__nor2_1 _27962_ (.A(_04242_),
    .B(_04231_),
    .Y(_04243_));
 sky130_fd_sc_hd__a211o_1 _27963_ (.A1(_04242_),
    .A2(net175),
    .B1(_04240_),
    .C1(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__nand2_1 _27964_ (.A(_04241_),
    .B(_04244_),
    .Y(_04246_));
 sky130_fd_sc_hd__mux2_1 _27965_ (.A0(_04232_),
    .A1(net175),
    .S(net168),
    .X(_04247_));
 sky130_fd_sc_hd__nor2_1 _27966_ (.A(_04205_),
    .B(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21oi_1 _27967_ (.A1(_04246_),
    .A2(_04205_),
    .B1(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__nor2_1 _27968_ (.A(_04222_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__a211o_1 _27969_ (.A1(_04222_),
    .A2(net176),
    .B1(net160),
    .C1(_04250_),
    .X(_04251_));
 sky130_fd_sc_hd__inv_2 _27970_ (.A(_04251_),
    .Y(_00014_));
 sky130_fd_sc_hd__nor2_4 _27971_ (.A(_02155_),
    .B(_02522_),
    .Y(_04252_));
 sky130_fd_sc_hd__inv_2 _27972_ (.A(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__or2_1 _27973_ (.A(_04230_),
    .B(_04253_),
    .X(_04254_));
 sky130_fd_sc_hd__nand2_1 _27974_ (.A(_04253_),
    .B(_04230_),
    .Y(_04256_));
 sky130_fd_sc_hd__nand2_1 _27975_ (.A(_04254_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_8 _27976_ (.A(_04209_),
    .B(_04207_),
    .Y(_04258_));
 sky130_fd_sc_hd__buf_6 _27977_ (.A(_04240_),
    .X(_04259_));
 sky130_fd_sc_hd__nand2_1 _27978_ (.A(_04258_),
    .B(_04252_),
    .Y(_04260_));
 sky130_fd_sc_hd__o211ai_1 _27979_ (.A1(_04257_),
    .A2(_04258_),
    .B1(_04259_),
    .C1(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__buf_6 _27980_ (.A(_04240_),
    .X(_04262_));
 sky130_fd_sc_hd__nor2_1 _27981_ (.A(_04194_),
    .B(_04257_),
    .Y(_04263_));
 sky130_fd_sc_hd__a211o_1 _27982_ (.A1(_04194_),
    .A2(_04252_),
    .B1(_04262_),
    .C1(_04263_),
    .X(_04264_));
 sky130_fd_sc_hd__nand2_1 _27983_ (.A(_04261_),
    .B(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__nand2_1 _27984_ (.A(_04265_),
    .B(_04205_),
    .Y(_04267_));
 sky130_fd_sc_hd__clkbuf_1 _27985_ (.A(net168),
    .X(_04268_));
 sky130_fd_sc_hd__mux2_1 _27986_ (.A0(_04257_),
    .A1(_04253_),
    .S(net169),
    .X(_04269_));
 sky130_fd_sc_hd__buf_6 _27987_ (.A(_04203_),
    .X(_04270_));
 sky130_fd_sc_hd__nand2_1 _27988_ (.A(net170),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand2_1 _27989_ (.A(_04267_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__inv_2 _27990_ (.A(_04221_),
    .Y(_04273_));
 sky130_fd_sc_hd__buf_6 _27991_ (.A(_04273_),
    .X(_04274_));
 sky130_fd_sc_hd__buf_6 _27992_ (.A(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__buf_6 _27993_ (.A(_04275_),
    .X(_04276_));
 sky130_fd_sc_hd__nor2_1 _27994_ (.A(_04276_),
    .B(_04252_),
    .Y(_04278_));
 sky130_fd_sc_hd__a211o_1 _27995_ (.A1(_04272_),
    .A2(_04276_),
    .B1(net160),
    .C1(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__inv_2 _27996_ (.A(_04279_),
    .Y(_00025_));
 sky130_fd_sc_hd__nor2_1 _27997_ (.A(_02170_),
    .B(_02524_),
    .Y(_04280_));
 sky130_fd_sc_hd__inv_4 _27998_ (.A(net184),
    .Y(_04281_));
 sky130_fd_sc_hd__buf_6 _27999_ (.A(_04182_),
    .X(_04282_));
 sky130_fd_sc_hd__or2_1 _28000_ (.A(_04254_),
    .B(_04281_),
    .X(_04283_));
 sky130_fd_sc_hd__nand2_1 _28001_ (.A(_04281_),
    .B(_04254_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_1 _28002_ (.A(_04283_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__inv_2 _28003_ (.A(_04285_),
    .Y(_04286_));
 sky130_fd_sc_hd__nand2_1 _28004_ (.A(_04282_),
    .B(_04286_),
    .Y(_04288_));
 sky130_fd_sc_hd__buf_8 _28005_ (.A(_04237_),
    .X(_04289_));
 sky130_fd_sc_hd__nand3_1 _28006_ (.A(_04289_),
    .B(net169),
    .C(net184),
    .Y(_04290_));
 sky130_fd_sc_hd__nand3_1 _28007_ (.A(_04288_),
    .B(_04290_),
    .C(_04259_),
    .Y(_04291_));
 sky130_fd_sc_hd__buf_6 _28008_ (.A(_04192_),
    .X(_04292_));
 sky130_fd_sc_hd__nor2_1 _28009_ (.A(_04292_),
    .B(_04281_),
    .Y(_04293_));
 sky130_fd_sc_hd__a211o_1 _28010_ (.A1(_04286_),
    .A2(_04292_),
    .B1(_04240_),
    .C1(_04293_),
    .X(_04294_));
 sky130_fd_sc_hd__nand2_1 _28011_ (.A(_04291_),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_1 _28012_ (.A(_04295_),
    .B(_04205_),
    .Y(_04296_));
 sky130_fd_sc_hd__mux2_1 _28013_ (.A0(_04285_),
    .A1(_04281_),
    .S(net168),
    .X(_04297_));
 sky130_fd_sc_hd__nand2_1 _28014_ (.A(_04297_),
    .B(_04270_),
    .Y(_04299_));
 sky130_fd_sc_hd__nand2_1 _28015_ (.A(_04296_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__and2_1 _28016_ (.A(_04300_),
    .B(_04276_),
    .X(_04301_));
 sky130_fd_sc_hd__a211o_1 _28017_ (.A1(_04222_),
    .A2(_04281_),
    .B1(net160),
    .C1(_04301_),
    .X(_04302_));
 sky130_fd_sc_hd__inv_2 _28018_ (.A(_04302_),
    .Y(_00028_));
 sky130_fd_sc_hd__nor2_4 _28019_ (.A(_02193_),
    .B(net196),
    .Y(_04303_));
 sky130_fd_sc_hd__inv_2 _28020_ (.A(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__or2_1 _28021_ (.A(_04283_),
    .B(_04304_),
    .X(_04305_));
 sky130_fd_sc_hd__nand2_1 _28022_ (.A(_04304_),
    .B(_04283_),
    .Y(_04306_));
 sky130_fd_sc_hd__nand2_1 _28023_ (.A(_04305_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__nand3_1 _28024_ (.A(net131),
    .B(_04210_),
    .C(_04307_),
    .Y(_04309_));
 sky130_fd_sc_hd__buf_6 _28025_ (.A(_04209_),
    .X(_04310_));
 sky130_fd_sc_hd__nand3_1 _28026_ (.A(_04207_),
    .B(_04310_),
    .C(_04307_),
    .Y(_04311_));
 sky130_fd_sc_hd__o21a_1 _28027_ (.A1(_04310_),
    .A2(_04303_),
    .B1(_04203_),
    .X(_04312_));
 sky130_fd_sc_hd__nand3_1 _28028_ (.A(_04309_),
    .B(_04311_),
    .C(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__nand2_1 _28029_ (.A(_04313_),
    .B(_04274_),
    .Y(_04314_));
 sky130_fd_sc_hd__inv_2 _28030_ (.A(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__inv_2 _28031_ (.A(_04307_),
    .Y(_04316_));
 sky130_fd_sc_hd__nand2_1 _28032_ (.A(_04282_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__buf_6 _28033_ (.A(_04236_),
    .X(_04318_));
 sky130_fd_sc_hd__nand3_1 _28034_ (.A(_04318_),
    .B(_04238_),
    .C(_04303_),
    .Y(_04320_));
 sky130_fd_sc_hd__nand3_1 _28035_ (.A(_04317_),
    .B(_04320_),
    .C(_04259_),
    .Y(_04321_));
 sky130_fd_sc_hd__mux2_1 _28036_ (.A0(_04307_),
    .A1(_04304_),
    .S(_04193_),
    .X(_04322_));
 sky130_fd_sc_hd__buf_6 _28037_ (.A(_04189_),
    .X(_04323_));
 sky130_fd_sc_hd__a21oi_1 _28038_ (.A1(_04322_),
    .A2(_04323_),
    .B1(_04270_),
    .Y(_04324_));
 sky130_fd_sc_hd__nand2_1 _28039_ (.A(_04321_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__nand2_1 _28040_ (.A(_04315_),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__buf_6 _28041_ (.A(_04221_),
    .X(_04327_));
 sky130_fd_sc_hd__nand2_1 _28042_ (.A(_04304_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__nand2_1 _28043_ (.A(_04326_),
    .B(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__or2_1 _28044_ (.A(_02652_),
    .B(_04329_),
    .X(_04331_));
 sky130_fd_sc_hd__inv_2 _28045_ (.A(_04331_),
    .Y(_00029_));
 sky130_fd_sc_hd__nor2_1 _28046_ (.A(_02195_),
    .B(net198),
    .Y(_04332_));
 sky130_fd_sc_hd__inv_1 _28047_ (.A(net199),
    .Y(_04333_));
 sky130_fd_sc_hd__or2_1 _28048_ (.A(_04305_),
    .B(_04333_),
    .X(_04334_));
 sky130_fd_sc_hd__nand2_1 _28049_ (.A(_04333_),
    .B(_04305_),
    .Y(_04335_));
 sky130_fd_sc_hd__nand2_1 _28050_ (.A(_04334_),
    .B(_04335_),
    .Y(_04336_));
 sky130_fd_sc_hd__inv_2 _28051_ (.A(_04336_),
    .Y(_04337_));
 sky130_fd_sc_hd__nand2_1 _28052_ (.A(_04282_),
    .B(_04337_),
    .Y(_04338_));
 sky130_fd_sc_hd__nand3_1 _28053_ (.A(_04318_),
    .B(net169),
    .C(net199),
    .Y(_04339_));
 sky130_fd_sc_hd__nand3_1 _28054_ (.A(_04338_),
    .B(_04339_),
    .C(_04259_),
    .Y(_04341_));
 sky130_fd_sc_hd__mux2_1 _28055_ (.A0(_04336_),
    .A1(_04333_),
    .S(_04242_),
    .X(_04342_));
 sky130_fd_sc_hd__a21oi_1 _28056_ (.A1(_04342_),
    .A2(_04323_),
    .B1(_04270_),
    .Y(_04343_));
 sky130_fd_sc_hd__nand2_1 _28057_ (.A(_04341_),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hd__buf_6 _28058_ (.A(_04274_),
    .X(_04345_));
 sky130_fd_sc_hd__nor2_2 _28059_ (.A(net168),
    .B(_04236_),
    .Y(_04346_));
 sky130_fd_sc_hd__buf_6 _28060_ (.A(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__nand2_1 _28061_ (.A(_04347_),
    .B(_04336_),
    .Y(_04348_));
 sky130_fd_sc_hd__nand3_1 _28062_ (.A(_04289_),
    .B(_04211_),
    .C(_04336_),
    .Y(_04349_));
 sky130_fd_sc_hd__buf_6 _28063_ (.A(_04310_),
    .X(_04350_));
 sky130_fd_sc_hd__buf_6 _28064_ (.A(_04203_),
    .X(_04352_));
 sky130_fd_sc_hd__o21a_1 _28065_ (.A1(_04350_),
    .A2(net199),
    .B1(_04352_),
    .X(_04353_));
 sky130_fd_sc_hd__nand3_1 _28066_ (.A(_04348_),
    .B(_04349_),
    .C(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__nand3_1 _28067_ (.A(_04344_),
    .B(_04345_),
    .C(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__nand2_1 _28068_ (.A(_04333_),
    .B(_04222_),
    .Y(_04356_));
 sky130_fd_sc_hd__nand2_1 _28069_ (.A(_04355_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__or2_1 _28070_ (.A(_02652_),
    .B(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__inv_2 _28071_ (.A(_04358_),
    .Y(_00030_));
 sky130_fd_sc_hd__nor2_4 _28072_ (.A(_02199_),
    .B(_02531_),
    .Y(_04359_));
 sky130_fd_sc_hd__inv_2 _28073_ (.A(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__or2_1 _28074_ (.A(_04334_),
    .B(_04360_),
    .X(_04362_));
 sky130_fd_sc_hd__nand2_1 _28075_ (.A(_04360_),
    .B(_04334_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _28076_ (.A(_04362_),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__inv_2 _28077_ (.A(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__nand2_1 _28078_ (.A(_04183_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__nand3_1 _28079_ (.A(net131),
    .B(_04238_),
    .C(_04359_),
    .Y(_04367_));
 sky130_fd_sc_hd__nand3_1 _28080_ (.A(_04366_),
    .B(_04367_),
    .C(_04262_),
    .Y(_04368_));
 sky130_fd_sc_hd__mux2_1 _28081_ (.A0(_04364_),
    .A1(_04360_),
    .S(_04193_),
    .X(_04369_));
 sky130_fd_sc_hd__a21oi_1 _28082_ (.A1(_04369_),
    .A2(_04323_),
    .B1(_04352_),
    .Y(_04370_));
 sky130_fd_sc_hd__nand2_1 _28083_ (.A(_04368_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__nand2_1 _28084_ (.A(_04347_),
    .B(_04364_),
    .Y(_04373_));
 sky130_fd_sc_hd__nand3_1 _28085_ (.A(_04318_),
    .B(_04211_),
    .C(_04364_),
    .Y(_04374_));
 sky130_fd_sc_hd__o21a_1 _28086_ (.A1(_04350_),
    .A2(_04359_),
    .B1(_04352_),
    .X(_04375_));
 sky130_fd_sc_hd__nand3_1 _28087_ (.A(_04373_),
    .B(_04374_),
    .C(_04375_),
    .Y(_04376_));
 sky130_fd_sc_hd__nand3_1 _28088_ (.A(_04371_),
    .B(_04345_),
    .C(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__nand2_1 _28089_ (.A(_04360_),
    .B(_04327_),
    .Y(_04378_));
 sky130_fd_sc_hd__nand2_1 _28090_ (.A(_04377_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__or2_1 _28091_ (.A(_02652_),
    .B(_04379_),
    .X(_04380_));
 sky130_fd_sc_hd__inv_2 _28092_ (.A(_04380_),
    .Y(_00031_));
 sky130_fd_sc_hd__nor2_4 _28093_ (.A(_02234_),
    .B(net213),
    .Y(_04381_));
 sky130_fd_sc_hd__clkinvlp_2 _28094_ (.A(_04381_),
    .Y(_04383_));
 sky130_fd_sc_hd__or2_1 _28095_ (.A(_04362_),
    .B(_04383_),
    .X(_04384_));
 sky130_fd_sc_hd__nand2_1 _28096_ (.A(_04383_),
    .B(_04362_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _28097_ (.A(_04384_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hd__nand3_1 _28098_ (.A(_04236_),
    .B(_04210_),
    .C(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__nand3_1 _28099_ (.A(_04207_),
    .B(_04310_),
    .C(_04386_),
    .Y(_04388_));
 sky130_fd_sc_hd__o21a_1 _28100_ (.A1(_04310_),
    .A2(_04381_),
    .B1(_04203_),
    .X(_04389_));
 sky130_fd_sc_hd__nand3_1 _28101_ (.A(_04387_),
    .B(_04388_),
    .C(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hd__nand2_1 _28102_ (.A(_04390_),
    .B(_04273_),
    .Y(_04391_));
 sky130_fd_sc_hd__inv_2 _28103_ (.A(_04391_),
    .Y(_04392_));
 sky130_fd_sc_hd__inv_2 _28104_ (.A(_04386_),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _28105_ (.A(_04282_),
    .B(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand3_1 _28106_ (.A(_04318_),
    .B(_04238_),
    .C(_04381_),
    .Y(_04396_));
 sky130_fd_sc_hd__nand3_1 _28107_ (.A(_04395_),
    .B(_04396_),
    .C(_04262_),
    .Y(_04397_));
 sky130_fd_sc_hd__mux2_1 _28108_ (.A0(_04386_),
    .A1(_04383_),
    .S(_04193_),
    .X(_04398_));
 sky130_fd_sc_hd__a21oi_1 _28109_ (.A1(_04398_),
    .A2(_04323_),
    .B1(_04270_),
    .Y(_04399_));
 sky130_fd_sc_hd__nand2_1 _28110_ (.A(_04397_),
    .B(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__nand2_1 _28111_ (.A(_04392_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _28112_ (.A(_04383_),
    .B(_04221_),
    .Y(_04402_));
 sky130_fd_sc_hd__nand2_1 _28113_ (.A(_04401_),
    .B(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__or2_1 _28114_ (.A(_02652_),
    .B(_04403_),
    .X(_04405_));
 sky130_fd_sc_hd__inv_2 _28115_ (.A(_04405_),
    .Y(_00032_));
 sky130_fd_sc_hd__nor2_4 _28116_ (.A(_02237_),
    .B(_02535_),
    .Y(_04406_));
 sky130_fd_sc_hd__inv_1 _28117_ (.A(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__or2_1 _28118_ (.A(_04384_),
    .B(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__nand2_1 _28119_ (.A(_04407_),
    .B(_04384_),
    .Y(_04409_));
 sky130_fd_sc_hd__nand2_1 _28120_ (.A(_04408_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nand3_1 _28121_ (.A(_04236_),
    .B(_04210_),
    .C(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand3_1 _28122_ (.A(_04207_),
    .B(_04310_),
    .C(_04410_),
    .Y(_04412_));
 sky130_fd_sc_hd__o21a_1 _28123_ (.A1(_04209_),
    .A2(_04406_),
    .B1(_04203_),
    .X(_04413_));
 sky130_fd_sc_hd__nand3_1 _28124_ (.A(_04411_),
    .B(_04412_),
    .C(_04413_),
    .Y(_04415_));
 sky130_fd_sc_hd__nand2_1 _28125_ (.A(_04415_),
    .B(_04273_),
    .Y(_04416_));
 sky130_fd_sc_hd__inv_2 _28126_ (.A(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__inv_2 _28127_ (.A(_04410_),
    .Y(_04418_));
 sky130_fd_sc_hd__nand2_1 _28128_ (.A(_04183_),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__nand3_1 _28129_ (.A(_04237_),
    .B(_04238_),
    .C(_04406_),
    .Y(_04420_));
 sky130_fd_sc_hd__nand3_1 _28130_ (.A(_04419_),
    .B(_04420_),
    .C(_04262_),
    .Y(_04421_));
 sky130_fd_sc_hd__nor2_1 _28131_ (.A(_04192_),
    .B(_04407_),
    .Y(_04422_));
 sky130_fd_sc_hd__nor2_1 _28132_ (.A(_04242_),
    .B(_04410_),
    .Y(_04423_));
 sky130_fd_sc_hd__o31a_1 _28133_ (.A1(_04188_),
    .A2(_04422_),
    .A3(_04423_),
    .B1(_04212_),
    .X(_04424_));
 sky130_fd_sc_hd__nand2_1 _28134_ (.A(_04421_),
    .B(_04424_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand2_1 _28135_ (.A(_04417_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_1 _28136_ (.A(_04407_),
    .B(_04327_),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_1 _28137_ (.A(_04427_),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__or2_1 _28138_ (.A(_02652_),
    .B(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__inv_2 _28139_ (.A(_04430_),
    .Y(_00033_));
 sky130_fd_sc_hd__nor2_4 _28140_ (.A(_02239_),
    .B(_02537_),
    .Y(_04431_));
 sky130_fd_sc_hd__inv_2 _28141_ (.A(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__or2_1 _28142_ (.A(_04408_),
    .B(_04432_),
    .X(_04433_));
 sky130_fd_sc_hd__nand2_1 _28143_ (.A(_04432_),
    .B(_04408_),
    .Y(_04434_));
 sky130_fd_sc_hd__nand2_1 _28144_ (.A(_04433_),
    .B(_04434_),
    .Y(_04436_));
 sky130_fd_sc_hd__nand3_1 _28145_ (.A(_04237_),
    .B(_04210_),
    .C(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__nand3_1 _28146_ (.A(_04207_),
    .B(_04210_),
    .C(_04436_),
    .Y(_04438_));
 sky130_fd_sc_hd__o21a_1 _28147_ (.A1(_04310_),
    .A2(_04431_),
    .B1(_04203_),
    .X(_04439_));
 sky130_fd_sc_hd__nand3_1 _28148_ (.A(_04437_),
    .B(_04438_),
    .C(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__nand2_1 _28149_ (.A(_04440_),
    .B(_04274_),
    .Y(_04441_));
 sky130_fd_sc_hd__inv_2 _28150_ (.A(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__nand2_1 _28151_ (.A(_04258_),
    .B(_04431_),
    .Y(_04443_));
 sky130_fd_sc_hd__clkinvlp_2 _28152_ (.A(_04436_),
    .Y(_04444_));
 sky130_fd_sc_hd__nand2_1 _28153_ (.A(_04183_),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__nand3_1 _28154_ (.A(_04443_),
    .B(_04445_),
    .C(_04259_),
    .Y(_04447_));
 sky130_fd_sc_hd__nand2_1 _28155_ (.A(_04444_),
    .B(_04292_),
    .Y(_04448_));
 sky130_fd_sc_hd__nand2_1 _28156_ (.A(_04431_),
    .B(_04194_),
    .Y(_04449_));
 sky130_fd_sc_hd__a31oi_1 _28157_ (.A1(_04448_),
    .A2(_04323_),
    .A3(_04449_),
    .B1(_04270_),
    .Y(_04450_));
 sky130_fd_sc_hd__nand2_1 _28158_ (.A(_04447_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__nand2_1 _28159_ (.A(_04442_),
    .B(_04451_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_1 _28160_ (.A(_04432_),
    .B(_04327_),
    .Y(_04453_));
 sky130_fd_sc_hd__nand2_1 _28161_ (.A(_04452_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__or2_1 _28162_ (.A(_02652_),
    .B(_04454_),
    .X(_04455_));
 sky130_fd_sc_hd__inv_2 _28163_ (.A(_04455_),
    .Y(_00034_));
 sky130_fd_sc_hd__nor2_4 _28164_ (.A(_02294_),
    .B(_02540_),
    .Y(_04457_));
 sky130_fd_sc_hd__inv_2 _28165_ (.A(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__or2_1 _28166_ (.A(_04433_),
    .B(_04458_),
    .X(_04459_));
 sky130_fd_sc_hd__nand2_1 _28167_ (.A(_04458_),
    .B(_04433_),
    .Y(_04460_));
 sky130_fd_sc_hd__nand2_1 _28168_ (.A(_04459_),
    .B(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand3_1 _28169_ (.A(_04236_),
    .B(_04210_),
    .C(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand3_1 _28170_ (.A(_04207_),
    .B(_04310_),
    .C(_04461_),
    .Y(_04463_));
 sky130_fd_sc_hd__o21a_1 _28171_ (.A1(_04209_),
    .A2(_04457_),
    .B1(_04203_),
    .X(_04464_));
 sky130_fd_sc_hd__nand3_1 _28172_ (.A(_04462_),
    .B(_04463_),
    .C(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__nand2_1 _28173_ (.A(_04465_),
    .B(_04273_),
    .Y(_04466_));
 sky130_fd_sc_hd__inv_2 _28174_ (.A(_04466_),
    .Y(_04468_));
 sky130_fd_sc_hd__inv_2 _28175_ (.A(_04461_),
    .Y(_04469_));
 sky130_fd_sc_hd__nand2_1 _28176_ (.A(_04183_),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__nand3_1 _28177_ (.A(_04318_),
    .B(_04238_),
    .C(_04457_),
    .Y(_04471_));
 sky130_fd_sc_hd__nand3_1 _28178_ (.A(_04470_),
    .B(_04471_),
    .C(_04262_),
    .Y(_04472_));
 sky130_fd_sc_hd__nor2_1 _28179_ (.A(_04192_),
    .B(_04458_),
    .Y(_04473_));
 sky130_fd_sc_hd__nor2_1 _28180_ (.A(_04242_),
    .B(_04461_),
    .Y(_04474_));
 sky130_fd_sc_hd__o31a_1 _28181_ (.A1(_04188_),
    .A2(_04473_),
    .A3(_04474_),
    .B1(_04212_),
    .X(_04475_));
 sky130_fd_sc_hd__nand2_1 _28182_ (.A(_04472_),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__nand2_1 _28183_ (.A(_04468_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand2_1 _28184_ (.A(_04458_),
    .B(_04327_),
    .Y(_04479_));
 sky130_fd_sc_hd__nand2_1 _28185_ (.A(_04477_),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hd__or2_1 _28186_ (.A(_02652_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__inv_2 _28187_ (.A(_04481_),
    .Y(_00004_));
 sky130_fd_sc_hd__clkbuf_2 _28188_ (.A(net160),
    .X(_04482_));
 sky130_fd_sc_hd__nor2_4 _28189_ (.A(_02298_),
    .B(_02542_),
    .Y(_04483_));
 sky130_fd_sc_hd__clkinvlp_2 _28190_ (.A(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__or2_1 _28191_ (.A(_04459_),
    .B(_04484_),
    .X(_04485_));
 sky130_fd_sc_hd__nand2_1 _28192_ (.A(_04484_),
    .B(_04459_),
    .Y(_04486_));
 sky130_fd_sc_hd__nand2_1 _28193_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__inv_2 _28194_ (.A(_04487_),
    .Y(_04489_));
 sky130_fd_sc_hd__nand2_1 _28195_ (.A(_04282_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hd__nand3_1 _28196_ (.A(_04289_),
    .B(net169),
    .C(_04483_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand3_1 _28197_ (.A(_04490_),
    .B(_04491_),
    .C(_04259_),
    .Y(_04492_));
 sky130_fd_sc_hd__nand2_1 _28198_ (.A(_04489_),
    .B(_04292_),
    .Y(_04493_));
 sky130_fd_sc_hd__nand2_1 _28199_ (.A(_04483_),
    .B(_04194_),
    .Y(_04494_));
 sky130_fd_sc_hd__a31oi_1 _28200_ (.A1(_04493_),
    .A2(_04323_),
    .A3(_04494_),
    .B1(_04270_),
    .Y(_04495_));
 sky130_fd_sc_hd__nand2_1 _28201_ (.A(_04492_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__nand2_1 _28202_ (.A(_04347_),
    .B(_04487_),
    .Y(_04497_));
 sky130_fd_sc_hd__nand3_1 _28203_ (.A(_04289_),
    .B(_04211_),
    .C(_04487_),
    .Y(_04498_));
 sky130_fd_sc_hd__o21a_1 _28204_ (.A1(_04350_),
    .A2(_04483_),
    .B1(_04352_),
    .X(_04500_));
 sky130_fd_sc_hd__nand3_1 _28205_ (.A(_04497_),
    .B(_04498_),
    .C(_04500_),
    .Y(_04501_));
 sky130_fd_sc_hd__nand3_1 _28206_ (.A(_04496_),
    .B(_04275_),
    .C(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__nand2_1 _28207_ (.A(_04484_),
    .B(_04222_),
    .Y(_04503_));
 sky130_fd_sc_hd__nand2_1 _28208_ (.A(_04502_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__or2_1 _28209_ (.A(_04482_),
    .B(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__inv_2 _28210_ (.A(_04505_),
    .Y(_00005_));
 sky130_fd_sc_hd__nor2_4 _28211_ (.A(_02301_),
    .B(_02544_),
    .Y(_04506_));
 sky130_fd_sc_hd__inv_2 _28212_ (.A(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__or2_1 _28213_ (.A(_04485_),
    .B(_04507_),
    .X(_04508_));
 sky130_fd_sc_hd__nand2_1 _28214_ (.A(_04507_),
    .B(_04485_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand2_1 _28215_ (.A(_04508_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__inv_2 _28216_ (.A(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hd__nand2_1 _28217_ (.A(_04282_),
    .B(_04512_),
    .Y(_04513_));
 sky130_fd_sc_hd__nand3_1 _28218_ (.A(_04289_),
    .B(net169),
    .C(_04506_),
    .Y(_04514_));
 sky130_fd_sc_hd__nand3_1 _28219_ (.A(_04513_),
    .B(_04514_),
    .C(_04259_),
    .Y(_04515_));
 sky130_fd_sc_hd__nor2_1 _28220_ (.A(_04292_),
    .B(_04507_),
    .Y(_04516_));
 sky130_fd_sc_hd__nor2_1 _28221_ (.A(_04194_),
    .B(_04511_),
    .Y(_04517_));
 sky130_fd_sc_hd__o31a_1 _28222_ (.A1(_04240_),
    .A2(_04516_),
    .A3(_04517_),
    .B1(_04205_),
    .X(_04518_));
 sky130_fd_sc_hd__nand2_1 _28223_ (.A(_04515_),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hd__nand2_1 _28224_ (.A(_04347_),
    .B(_04511_),
    .Y(_04521_));
 sky130_fd_sc_hd__nand3_1 _28225_ (.A(_04289_),
    .B(_04211_),
    .C(_04511_),
    .Y(_04522_));
 sky130_fd_sc_hd__o21a_1 _28226_ (.A1(_04350_),
    .A2(_04506_),
    .B1(_04270_),
    .X(_04523_));
 sky130_fd_sc_hd__nand3_1 _28227_ (.A(_04521_),
    .B(_04522_),
    .C(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__nand3_1 _28228_ (.A(_04519_),
    .B(_04275_),
    .C(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__nand2_1 _28229_ (.A(_04507_),
    .B(_04222_),
    .Y(_04526_));
 sky130_fd_sc_hd__nand2_1 _28230_ (.A(_04525_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__or2_1 _28231_ (.A(_04482_),
    .B(_04527_),
    .X(_04528_));
 sky130_fd_sc_hd__inv_2 _28232_ (.A(_04528_),
    .Y(_00006_));
 sky130_fd_sc_hd__nor2_4 _28233_ (.A(_02349_),
    .B(_02546_),
    .Y(_04529_));
 sky130_fd_sc_hd__inv_2 _28234_ (.A(_04529_),
    .Y(_04531_));
 sky130_fd_sc_hd__or2_1 _28235_ (.A(_04508_),
    .B(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__nand2_1 _28236_ (.A(_04531_),
    .B(_04508_),
    .Y(_04533_));
 sky130_fd_sc_hd__nand2_1 _28237_ (.A(_04532_),
    .B(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand3_1 _28238_ (.A(_04237_),
    .B(_04210_),
    .C(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand3_1 _28239_ (.A(_04207_),
    .B(_04210_),
    .C(_04534_),
    .Y(_04536_));
 sky130_fd_sc_hd__o21a_1 _28240_ (.A1(_04310_),
    .A2(_04529_),
    .B1(_04203_),
    .X(_04537_));
 sky130_fd_sc_hd__nand3_1 _28241_ (.A(_04535_),
    .B(_04536_),
    .C(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_1 _28242_ (.A(_04538_),
    .B(_04274_),
    .Y(_04539_));
 sky130_fd_sc_hd__inv_2 _28243_ (.A(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2_1 _28244_ (.A(_04258_),
    .B(_04529_),
    .Y(_04542_));
 sky130_fd_sc_hd__inv_2 _28245_ (.A(_04534_),
    .Y(_04543_));
 sky130_fd_sc_hd__nand2_1 _28246_ (.A(_04282_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__nand3_1 _28247_ (.A(_04542_),
    .B(_04544_),
    .C(_04259_),
    .Y(_04545_));
 sky130_fd_sc_hd__nand2_1 _28248_ (.A(_04543_),
    .B(_04292_),
    .Y(_04546_));
 sky130_fd_sc_hd__nand2_1 _28249_ (.A(_04529_),
    .B(_04194_),
    .Y(_04547_));
 sky130_fd_sc_hd__a31oi_1 _28250_ (.A1(_04546_),
    .A2(_04323_),
    .A3(_04547_),
    .B1(_04270_),
    .Y(_04548_));
 sky130_fd_sc_hd__nand2_1 _28251_ (.A(_04545_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__nand2_1 _28252_ (.A(_04540_),
    .B(_04549_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand2_1 _28253_ (.A(_04531_),
    .B(_04327_),
    .Y(_04551_));
 sky130_fd_sc_hd__nand2_1 _28254_ (.A(_04550_),
    .B(_04551_),
    .Y(_04553_));
 sky130_fd_sc_hd__or2_1 _28255_ (.A(_04482_),
    .B(_04553_),
    .X(_04554_));
 sky130_fd_sc_hd__inv_2 _28256_ (.A(_04554_),
    .Y(_00007_));
 sky130_fd_sc_hd__nor2_4 _28257_ (.A(_02363_),
    .B(_02548_),
    .Y(_04555_));
 sky130_fd_sc_hd__inv_2 _28258_ (.A(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__or2_1 _28259_ (.A(_04532_),
    .B(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__nand2_1 _28260_ (.A(_04556_),
    .B(_04532_),
    .Y(_04558_));
 sky130_fd_sc_hd__nand2_1 _28261_ (.A(_04557_),
    .B(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__inv_2 _28262_ (.A(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__nand2_1 _28263_ (.A(_04282_),
    .B(_04560_),
    .Y(_04561_));
 sky130_fd_sc_hd__nand3_1 _28264_ (.A(_04318_),
    .B(net169),
    .C(_04555_),
    .Y(_04563_));
 sky130_fd_sc_hd__nand3_1 _28265_ (.A(_04561_),
    .B(_04563_),
    .C(_04259_),
    .Y(_04564_));
 sky130_fd_sc_hd__nor2_1 _28266_ (.A(_04192_),
    .B(_04556_),
    .Y(_04565_));
 sky130_fd_sc_hd__nor2_1 _28267_ (.A(_04242_),
    .B(_04559_),
    .Y(_04566_));
 sky130_fd_sc_hd__o31a_1 _28268_ (.A1(_04240_),
    .A2(_04565_),
    .A3(_04566_),
    .B1(_04212_),
    .X(_04567_));
 sky130_fd_sc_hd__nand2_1 _28269_ (.A(_04564_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__nand2_1 _28270_ (.A(_04347_),
    .B(_04559_),
    .Y(_04569_));
 sky130_fd_sc_hd__nand3_1 _28271_ (.A(_04289_),
    .B(_04211_),
    .C(_04559_),
    .Y(_04570_));
 sky130_fd_sc_hd__o21a_1 _28272_ (.A1(_04350_),
    .A2(_04555_),
    .B1(_04352_),
    .X(_04571_));
 sky130_fd_sc_hd__nand3_1 _28273_ (.A(_04569_),
    .B(_04570_),
    .C(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand3_1 _28274_ (.A(_04568_),
    .B(_04345_),
    .C(_04572_),
    .Y(_04574_));
 sky130_fd_sc_hd__nand2_1 _28275_ (.A(_04556_),
    .B(_04222_),
    .Y(_04575_));
 sky130_fd_sc_hd__nand2_1 _28276_ (.A(_04574_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hd__or2_1 _28277_ (.A(_04482_),
    .B(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__inv_2 _28278_ (.A(_04577_),
    .Y(_00008_));
 sky130_fd_sc_hd__nand2_4 _28279_ (.A(_02551_),
    .B(_02421_),
    .Y(_04578_));
 sky130_fd_sc_hd__or2_1 _28280_ (.A(_04578_),
    .B(_04557_),
    .X(_04579_));
 sky130_fd_sc_hd__nand2_1 _28281_ (.A(_04557_),
    .B(_04578_),
    .Y(_04580_));
 sky130_fd_sc_hd__nand2_1 _28282_ (.A(_04579_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__inv_2 _28283_ (.A(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__nand2_1 _28284_ (.A(_04282_),
    .B(_04582_),
    .Y(_04584_));
 sky130_fd_sc_hd__clkinvlp_2 _28285_ (.A(_04578_),
    .Y(_04585_));
 sky130_fd_sc_hd__nand3_1 _28286_ (.A(_04318_),
    .B(_04238_),
    .C(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__nand3_1 _28287_ (.A(_04584_),
    .B(_04586_),
    .C(_04262_),
    .Y(_04587_));
 sky130_fd_sc_hd__nand2_1 _28288_ (.A(_04582_),
    .B(_04292_),
    .Y(_04588_));
 sky130_fd_sc_hd__nand2_1 _28289_ (.A(_04585_),
    .B(_04194_),
    .Y(_04589_));
 sky130_fd_sc_hd__a31oi_1 _28290_ (.A1(_04588_),
    .A2(_04323_),
    .A3(_04589_),
    .B1(_04352_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _28291_ (.A(_04587_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nand2_1 _28292_ (.A(_04347_),
    .B(_04581_),
    .Y(_04592_));
 sky130_fd_sc_hd__nand3_1 _28293_ (.A(_04289_),
    .B(_04211_),
    .C(_04581_),
    .Y(_04593_));
 sky130_fd_sc_hd__a21oi_1 _28294_ (.A1(_04578_),
    .A2(_04238_),
    .B1(_04212_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand3_1 _28295_ (.A(_04592_),
    .B(_04593_),
    .C(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__nand3_1 _28296_ (.A(_04591_),
    .B(_04345_),
    .C(_04596_),
    .Y(_04597_));
 sky130_fd_sc_hd__nand2_1 _28297_ (.A(_04578_),
    .B(_04327_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_1 _28298_ (.A(_04597_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__or2_1 _28299_ (.A(_04482_),
    .B(_04599_),
    .X(_04600_));
 sky130_fd_sc_hd__inv_2 _28300_ (.A(_04600_),
    .Y(_00009_));
 sky130_fd_sc_hd__nand2_1 _28301_ (.A(_04236_),
    .B(_04310_),
    .Y(_04601_));
 sky130_fd_sc_hd__or4_1 _28302_ (.A(_04485_),
    .B(_04507_),
    .C(_04531_),
    .D(_04556_),
    .X(_04602_));
 sky130_fd_sc_hd__nand2_4 _28303_ (.A(_02552_),
    .B(_02367_),
    .Y(_04603_));
 sky130_fd_sc_hd__or3_1 _28304_ (.A(_04578_),
    .B(_04602_),
    .C(_04603_),
    .X(_04605_));
 sky130_fd_sc_hd__nand2_1 _28305_ (.A(_04603_),
    .B(_04579_),
    .Y(_04606_));
 sky130_fd_sc_hd__nand2_2 _28306_ (.A(_04605_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__nand2b_1 _28307_ (.A_N(_04601_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__nand2_1 _28308_ (.A(_04347_),
    .B(_04607_),
    .Y(_04609_));
 sky130_fd_sc_hd__a21oi_1 _28309_ (.A1(_04603_),
    .A2(net169),
    .B1(_04205_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand3_1 _28310_ (.A(_04608_),
    .B(_04609_),
    .C(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__inv_2 _28311_ (.A(_04603_),
    .Y(_04612_));
 sky130_fd_sc_hd__nand2_1 _28312_ (.A(_04258_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__clkinvlp_2 _28313_ (.A(_04607_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2_1 _28314_ (.A(_04183_),
    .B(_04614_),
    .Y(_04616_));
 sky130_fd_sc_hd__nand3_1 _28315_ (.A(_04613_),
    .B(_04616_),
    .C(_04262_),
    .Y(_04617_));
 sky130_fd_sc_hd__nor2_1 _28316_ (.A(_04192_),
    .B(_04603_),
    .Y(_04618_));
 sky130_fd_sc_hd__nor2_1 _28317_ (.A(_04242_),
    .B(_04607_),
    .Y(_04619_));
 sky130_fd_sc_hd__o31a_1 _28318_ (.A1(_04188_),
    .A2(_04618_),
    .A3(_04619_),
    .B1(_04212_),
    .X(_04620_));
 sky130_fd_sc_hd__nand2_1 _28319_ (.A(_04617_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__nand3_1 _28320_ (.A(_04611_),
    .B(_04621_),
    .C(_04345_),
    .Y(_04622_));
 sky130_fd_sc_hd__nand2_1 _28321_ (.A(_04603_),
    .B(_04327_),
    .Y(_04623_));
 sky130_fd_sc_hd__nand2_1 _28322_ (.A(_04622_),
    .B(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__or2_1 _28323_ (.A(_04482_),
    .B(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__inv_2 _28324_ (.A(_04625_),
    .Y(_00010_));
 sky130_fd_sc_hd__nand2_4 _28325_ (.A(_02553_),
    .B(_02433_),
    .Y(_04627_));
 sky130_fd_sc_hd__clkinvlp_2 _28326_ (.A(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__or2_1 _28327_ (.A(_04627_),
    .B(_04605_),
    .X(_04629_));
 sky130_fd_sc_hd__nand2_1 _28328_ (.A(_04605_),
    .B(_04627_),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _28329_ (.A(_04629_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__inv_2 _28330_ (.A(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand2_1 _28331_ (.A(_04282_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__nand3_1 _28332_ (.A(_04318_),
    .B(net169),
    .C(_04628_),
    .Y(_04634_));
 sky130_fd_sc_hd__nand3_1 _28333_ (.A(_04633_),
    .B(_04634_),
    .C(_04259_),
    .Y(_04635_));
 sky130_fd_sc_hd__nand2_1 _28334_ (.A(_04632_),
    .B(_04292_),
    .Y(_04637_));
 sky130_fd_sc_hd__nand2_1 _28335_ (.A(_04628_),
    .B(_04194_),
    .Y(_04638_));
 sky130_fd_sc_hd__a31oi_1 _28336_ (.A1(_04637_),
    .A2(_04323_),
    .A3(_04638_),
    .B1(_04270_),
    .Y(_04639_));
 sky130_fd_sc_hd__nand2_1 _28337_ (.A(_04635_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2_1 _28338_ (.A(_04347_),
    .B(_04631_),
    .Y(_04641_));
 sky130_fd_sc_hd__nand3_1 _28339_ (.A(_04289_),
    .B(_04211_),
    .C(_04631_),
    .Y(_04642_));
 sky130_fd_sc_hd__a21oi_1 _28340_ (.A1(_04627_),
    .A2(net169),
    .B1(_04205_),
    .Y(_04643_));
 sky130_fd_sc_hd__nand3_1 _28341_ (.A(_04641_),
    .B(_04642_),
    .C(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hd__nand3_1 _28342_ (.A(_04640_),
    .B(_04345_),
    .C(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__o21ai_1 _28343_ (.A1(_04345_),
    .A2(_04628_),
    .B1(_04645_),
    .Y(_04646_));
 sky130_fd_sc_hd__or2_1 _28344_ (.A(_04482_),
    .B(_04646_),
    .X(_04648_));
 sky130_fd_sc_hd__inv_2 _28345_ (.A(_04648_),
    .Y(_00011_));
 sky130_fd_sc_hd__nand2_4 _28346_ (.A(_02554_),
    .B(_02436_),
    .Y(_04649_));
 sky130_fd_sc_hd__inv_2 _28347_ (.A(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__nand2_1 _28348_ (.A(_04258_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__or2_1 _28349_ (.A(_04629_),
    .B(_04649_),
    .X(_04652_));
 sky130_fd_sc_hd__nand2_1 _28350_ (.A(_04649_),
    .B(_04629_),
    .Y(_04653_));
 sky130_fd_sc_hd__nand2_1 _28351_ (.A(_04652_),
    .B(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__clkinvlp_2 _28352_ (.A(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hd__nand2_1 _28353_ (.A(_04183_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__nand3_1 _28354_ (.A(_04651_),
    .B(_04656_),
    .C(_04262_),
    .Y(_04658_));
 sky130_fd_sc_hd__nor2_1 _28355_ (.A(_04192_),
    .B(_04649_),
    .Y(_04659_));
 sky130_fd_sc_hd__nor2_1 _28356_ (.A(_04242_),
    .B(_04654_),
    .Y(_04660_));
 sky130_fd_sc_hd__o31a_1 _28357_ (.A1(_04240_),
    .A2(_04659_),
    .A3(_04660_),
    .B1(_04212_),
    .X(_04661_));
 sky130_fd_sc_hd__nand2_1 _28358_ (.A(_04658_),
    .B(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__nand2_1 _28359_ (.A(_04347_),
    .B(_04654_),
    .Y(_04663_));
 sky130_fd_sc_hd__nand3_1 _28360_ (.A(_04289_),
    .B(_04211_),
    .C(_04654_),
    .Y(_04664_));
 sky130_fd_sc_hd__a21oi_1 _28361_ (.A1(_04649_),
    .A2(net169),
    .B1(_04212_),
    .Y(_04665_));
 sky130_fd_sc_hd__nand3_1 _28362_ (.A(_04663_),
    .B(_04664_),
    .C(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__nand3_1 _28363_ (.A(_04662_),
    .B(_04345_),
    .C(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hd__nand2_1 _28364_ (.A(_04649_),
    .B(_04327_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand2_1 _28365_ (.A(_04667_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__or2_1 _28366_ (.A(_04482_),
    .B(_04670_),
    .X(_04671_));
 sky130_fd_sc_hd__inv_2 _28367_ (.A(_04671_),
    .Y(_00012_));
 sky130_fd_sc_hd__nor2_2 _28368_ (.A(_02511_),
    .B(_02556_),
    .Y(_04672_));
 sky130_fd_sc_hd__inv_2 _28369_ (.A(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__or2_1 _28370_ (.A(_04652_),
    .B(_04673_),
    .X(_04674_));
 sky130_fd_sc_hd__nand2_1 _28371_ (.A(_04673_),
    .B(_04652_),
    .Y(_04675_));
 sky130_fd_sc_hd__nand2_1 _28372_ (.A(_04674_),
    .B(_04675_),
    .Y(_04676_));
 sky130_fd_sc_hd__inv_2 _28373_ (.A(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand2_1 _28374_ (.A(_04183_),
    .B(_04677_),
    .Y(_04679_));
 sky130_fd_sc_hd__nand3_1 _28375_ (.A(_04237_),
    .B(_04238_),
    .C(_04672_),
    .Y(_04680_));
 sky130_fd_sc_hd__nand3_1 _28376_ (.A(_04679_),
    .B(_04680_),
    .C(_04262_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand2_1 _28377_ (.A(_04677_),
    .B(_04292_),
    .Y(_04682_));
 sky130_fd_sc_hd__nand2_1 _28378_ (.A(_04672_),
    .B(_04242_),
    .Y(_04683_));
 sky130_fd_sc_hd__a31oi_1 _28379_ (.A1(_04682_),
    .A2(_04189_),
    .A3(_04683_),
    .B1(_04352_),
    .Y(_04684_));
 sky130_fd_sc_hd__nand2_1 _28380_ (.A(_04681_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__nand2_1 _28381_ (.A(_04346_),
    .B(_04676_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand3_1 _28382_ (.A(_04318_),
    .B(_04350_),
    .C(_04676_),
    .Y(_04687_));
 sky130_fd_sc_hd__o21a_1 _28383_ (.A1(_04350_),
    .A2(_04672_),
    .B1(_04352_),
    .X(_04688_));
 sky130_fd_sc_hd__nand3_1 _28384_ (.A(_04686_),
    .B(_04687_),
    .C(_04688_),
    .Y(_04690_));
 sky130_fd_sc_hd__nand3_1 _28385_ (.A(_04685_),
    .B(_04274_),
    .C(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__nand2_1 _28386_ (.A(_04673_),
    .B(_04221_),
    .Y(_04692_));
 sky130_fd_sc_hd__nand2_1 _28387_ (.A(_04691_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__or2_1 _28388_ (.A(_04482_),
    .B(_04693_),
    .X(_04694_));
 sky130_fd_sc_hd__inv_2 _28389_ (.A(_04694_),
    .Y(_00013_));
 sky130_fd_sc_hd__nand2_2 _28390_ (.A(_02558_),
    .B(_02512_),
    .Y(_04695_));
 sky130_fd_sc_hd__inv_1 _28391_ (.A(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__nand2_1 _28392_ (.A(_04674_),
    .B(_04695_),
    .Y(_04697_));
 sky130_fd_sc_hd__or2_1 _28393_ (.A(_04695_),
    .B(_04674_),
    .X(_04698_));
 sky130_fd_sc_hd__nand3_1 _28394_ (.A(_04182_),
    .B(_04697_),
    .C(_04698_),
    .Y(_04700_));
 sky130_fd_sc_hd__nand2_1 _28395_ (.A(_04258_),
    .B(_04696_),
    .Y(_04701_));
 sky130_fd_sc_hd__nand3_1 _28396_ (.A(_04700_),
    .B(_04701_),
    .C(_04240_),
    .Y(_04702_));
 sky130_fd_sc_hd__nor2_1 _28397_ (.A(_04192_),
    .B(_04695_),
    .Y(_04703_));
 sky130_fd_sc_hd__nand2_1 _28398_ (.A(_04698_),
    .B(_04697_),
    .Y(_04704_));
 sky130_fd_sc_hd__nor2_1 _28399_ (.A(_04193_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__o31a_1 _28400_ (.A1(_04188_),
    .A2(_04703_),
    .A3(_04705_),
    .B1(_04204_),
    .X(_04706_));
 sky130_fd_sc_hd__nand2_1 _28401_ (.A(_04702_),
    .B(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__nand2_1 _28402_ (.A(_04346_),
    .B(_04704_),
    .Y(_04708_));
 sky130_fd_sc_hd__nand3_1 _28403_ (.A(net131),
    .B(_04350_),
    .C(_04704_),
    .Y(_04709_));
 sky130_fd_sc_hd__a21oi_1 _28404_ (.A1(_04695_),
    .A2(net168),
    .B1(_04212_),
    .Y(_04711_));
 sky130_fd_sc_hd__nand3_1 _28405_ (.A(_04708_),
    .B(_04709_),
    .C(_04711_),
    .Y(_04712_));
 sky130_fd_sc_hd__nand3_1 _28406_ (.A(_04707_),
    .B(_04274_),
    .C(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__o21ai_2 _28407_ (.A1(_04274_),
    .A2(_04696_),
    .B1(_04713_),
    .Y(_04714_));
 sky130_fd_sc_hd__or2_1 _28408_ (.A(_04482_),
    .B(_04714_),
    .X(_04715_));
 sky130_fd_sc_hd__inv_2 _28409_ (.A(_04715_),
    .Y(_00015_));
 sky130_fd_sc_hd__nor2_2 _28410_ (.A(_02564_),
    .B(_02562_),
    .Y(_04716_));
 sky130_fd_sc_hd__clkinvlp_2 _28411_ (.A(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__or2_1 _28412_ (.A(_04698_),
    .B(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__nand2_1 _28413_ (.A(_04717_),
    .B(_04698_),
    .Y(_04719_));
 sky130_fd_sc_hd__nand2_1 _28414_ (.A(_04718_),
    .B(_04719_),
    .Y(_04721_));
 sky130_fd_sc_hd__inv_2 _28415_ (.A(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _28416_ (.A(_04183_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__nand3_1 _28417_ (.A(net131),
    .B(_04238_),
    .C(_04716_),
    .Y(_04724_));
 sky130_fd_sc_hd__nand3_1 _28418_ (.A(_04723_),
    .B(_04724_),
    .C(_04262_),
    .Y(_04725_));
 sky130_fd_sc_hd__nand2_1 _28419_ (.A(_04722_),
    .B(_04292_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_1 _28420_ (.A(_04716_),
    .B(_04194_),
    .Y(_04727_));
 sky130_fd_sc_hd__a31oi_1 _28421_ (.A1(_04726_),
    .A2(_04323_),
    .A3(_04727_),
    .B1(_04352_),
    .Y(_04728_));
 sky130_fd_sc_hd__nand2_1 _28422_ (.A(_04725_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__nand2_1 _28423_ (.A(_04347_),
    .B(_04721_),
    .Y(_04730_));
 sky130_fd_sc_hd__nand3_1 _28424_ (.A(_04318_),
    .B(_04350_),
    .C(_04721_),
    .Y(_04732_));
 sky130_fd_sc_hd__o21a_1 _28425_ (.A1(_04350_),
    .A2(_04716_),
    .B1(_04352_),
    .X(_04733_));
 sky130_fd_sc_hd__nand3_1 _28426_ (.A(_04730_),
    .B(_04732_),
    .C(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__nand3_1 _28427_ (.A(_04729_),
    .B(_04345_),
    .C(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hd__nand2_1 _28428_ (.A(_04717_),
    .B(_04327_),
    .Y(_04736_));
 sky130_fd_sc_hd__nand2_1 _28429_ (.A(_04735_),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__or2_1 _28430_ (.A(net160),
    .B(_04737_),
    .X(_04738_));
 sky130_fd_sc_hd__inv_2 _28431_ (.A(_04738_),
    .Y(_00016_));
 sky130_fd_sc_hd__nor2_2 _28432_ (.A(_02567_),
    .B(_02565_),
    .Y(_04739_));
 sky130_fd_sc_hd__inv_2 _28433_ (.A(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__or2_1 _28434_ (.A(_04718_),
    .B(_04740_),
    .X(_04742_));
 sky130_fd_sc_hd__nand2_1 _28435_ (.A(_04740_),
    .B(_04718_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _28436_ (.A(_04742_),
    .B(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__nand2b_1 _28437_ (.A_N(_04744_),
    .B(_04182_),
    .Y(_04745_));
 sky130_fd_sc_hd__nand2_1 _28438_ (.A(_04258_),
    .B(_04739_),
    .Y(_04746_));
 sky130_fd_sc_hd__nand3_1 _28439_ (.A(_04745_),
    .B(_04240_),
    .C(_04746_),
    .Y(_04747_));
 sky130_fd_sc_hd__nor2_1 _28440_ (.A(_04192_),
    .B(_04740_),
    .Y(_04748_));
 sky130_fd_sc_hd__nor2_1 _28441_ (.A(_04242_),
    .B(_04744_),
    .Y(_04749_));
 sky130_fd_sc_hd__o31a_1 _28442_ (.A1(_04188_),
    .A2(_04748_),
    .A3(_04749_),
    .B1(_04212_),
    .X(_04750_));
 sky130_fd_sc_hd__nand2_1 _28443_ (.A(_04747_),
    .B(_04750_),
    .Y(_04751_));
 sky130_fd_sc_hd__nand2b_1 _28444_ (.A_N(_04601_),
    .B(_04744_),
    .Y(_04753_));
 sky130_fd_sc_hd__nand2_1 _28445_ (.A(_04346_),
    .B(_04744_),
    .Y(_04754_));
 sky130_fd_sc_hd__o21a_1 _28446_ (.A1(_04210_),
    .A2(_04739_),
    .B1(_04203_),
    .X(_04755_));
 sky130_fd_sc_hd__nand3_1 _28447_ (.A(_04753_),
    .B(_04754_),
    .C(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__nand3_1 _28448_ (.A(_04751_),
    .B(_04274_),
    .C(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _28449_ (.A(_04740_),
    .B(_04222_),
    .Y(_04758_));
 sky130_fd_sc_hd__nand2_1 _28450_ (.A(_04757_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hd__nand2_1 _28451_ (.A(_02134_),
    .B(net148),
    .Y(_04760_));
 sky130_fd_sc_hd__o21ai_1 _28452_ (.A1(_02652_),
    .A2(_04759_),
    .B1(net149),
    .Y(_00017_));
 sky130_fd_sc_hd__nand2_1 _28453_ (.A(_04379_),
    .B(_04359_),
    .Y(_04761_));
 sky130_fd_sc_hd__nand3_1 _28454_ (.A(_04377_),
    .B(_04275_),
    .C(_04360_),
    .Y(_04763_));
 sky130_fd_sc_hd__nand2_1 _28455_ (.A(_04761_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__nand2_1 _28456_ (.A(_04670_),
    .B(_04650_),
    .Y(_04765_));
 sky130_fd_sc_hd__buf_6 _28457_ (.A(_04274_),
    .X(_04766_));
 sky130_fd_sc_hd__nand3_1 _28458_ (.A(_04667_),
    .B(_04766_),
    .C(_04649_),
    .Y(_04767_));
 sky130_fd_sc_hd__nand2_1 _28459_ (.A(_04765_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__nor2_1 _28460_ (.A(_04764_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__nand3_1 _28461_ (.A(_04645_),
    .B(_04275_),
    .C(_04627_),
    .Y(_04770_));
 sky130_fd_sc_hd__nand3_1 _28462_ (.A(_04735_),
    .B(_04275_),
    .C(_04717_),
    .Y(_04771_));
 sky130_fd_sc_hd__nand2_1 _28463_ (.A(_04770_),
    .B(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__nand3_1 _28464_ (.A(_04713_),
    .B(_04766_),
    .C(_04695_),
    .Y(_04774_));
 sky130_fd_sc_hd__nand2_1 _28465_ (.A(_04737_),
    .B(_04716_),
    .Y(_04775_));
 sky130_fd_sc_hd__nand2_1 _28466_ (.A(_04774_),
    .B(_04775_),
    .Y(_04776_));
 sky130_fd_sc_hd__nor2_1 _28467_ (.A(_04772_),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__nand2_1 _28468_ (.A(_04769_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_1 _28469_ (.A(_04599_),
    .B(_04585_),
    .Y(_04779_));
 sky130_fd_sc_hd__nand3_1 _28470_ (.A(_04691_),
    .B(_04766_),
    .C(_04673_),
    .Y(_04780_));
 sky130_fd_sc_hd__nand2_1 _28471_ (.A(_04779_),
    .B(_04780_),
    .Y(_04781_));
 sky130_fd_sc_hd__nand2_1 _28472_ (.A(_04646_),
    .B(_04628_),
    .Y(_04782_));
 sky130_fd_sc_hd__nand2_1 _28473_ (.A(_04624_),
    .B(_04612_),
    .Y(_04783_));
 sky130_fd_sc_hd__nand2_1 _28474_ (.A(_04782_),
    .B(_04783_),
    .Y(_04785_));
 sky130_fd_sc_hd__nor2_1 _28475_ (.A(_04781_),
    .B(_04785_),
    .Y(_04786_));
 sky130_fd_sc_hd__nand3_1 _28476_ (.A(_04622_),
    .B(_04766_),
    .C(_04603_),
    .Y(_04787_));
 sky130_fd_sc_hd__nand2_1 _28477_ (.A(_04693_),
    .B(_04672_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand2_1 _28478_ (.A(_04787_),
    .B(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__nand3_1 _28479_ (.A(_04355_),
    .B(_04766_),
    .C(_04333_),
    .Y(_04790_));
 sky130_fd_sc_hd__o21ai_1 _28480_ (.A1(_04381_),
    .A2(_04403_),
    .B1(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__nor2_1 _28481_ (.A(_04789_),
    .B(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand2_1 _28482_ (.A(_04786_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__nor2_1 _28483_ (.A(_04778_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand3b_1 _28484_ (.A_N(_04216_),
    .B(_04208_),
    .C(_04276_),
    .Y(_04796_));
 sky130_fd_sc_hd__nand3_1 _28485_ (.A(_04216_),
    .B(net190),
    .C(_04276_),
    .Y(_04797_));
 sky130_fd_sc_hd__nand2_1 _28486_ (.A(_04796_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__nand2_1 _28487_ (.A(_04714_),
    .B(_04696_),
    .Y(_04799_));
 sky130_fd_sc_hd__nand3_1 _28488_ (.A(_04757_),
    .B(_04345_),
    .C(_04740_),
    .Y(_04800_));
 sky130_fd_sc_hd__nand2_1 _28489_ (.A(_04799_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__inv_2 _28490_ (.A(_04801_),
    .Y(_04802_));
 sky130_fd_sc_hd__a21oi_1 _28491_ (.A1(_04759_),
    .A2(_04739_),
    .B1(_04211_),
    .Y(_04803_));
 sky130_fd_sc_hd__nand2_1 _28492_ (.A(_04802_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__nor2_1 _28493_ (.A(_04798_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hd__nand2_1 _28494_ (.A(_04794_),
    .B(_04805_),
    .Y(_04807_));
 sky130_fd_sc_hd__nand2_1 _28495_ (.A(_04480_),
    .B(_04457_),
    .Y(_04808_));
 sky130_fd_sc_hd__nand3_1 _28496_ (.A(_04477_),
    .B(_04275_),
    .C(_04458_),
    .Y(_04809_));
 sky130_fd_sc_hd__nand2_1 _28497_ (.A(_04808_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__nand2_1 _28498_ (.A(_04454_),
    .B(_04431_),
    .Y(_04811_));
 sky130_fd_sc_hd__nand3_1 _28499_ (.A(_04452_),
    .B(_04766_),
    .C(_04432_),
    .Y(_04812_));
 sky130_fd_sc_hd__nand2_1 _28500_ (.A(_04811_),
    .B(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__nor2_1 _28501_ (.A(_04810_),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__nand3_1 _28502_ (.A(_04427_),
    .B(_04275_),
    .C(_04407_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand3_1 _28503_ (.A(_04550_),
    .B(_04275_),
    .C(_04531_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2_1 _28504_ (.A(_04815_),
    .B(_04816_),
    .Y(_04818_));
 sky130_fd_sc_hd__nand2_1 _28505_ (.A(_04403_),
    .B(_04381_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _28506_ (.A(_04429_),
    .B(_04406_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand2_1 _28507_ (.A(_04819_),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__nor2_1 _28508_ (.A(_04818_),
    .B(_04821_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand2_1 _28509_ (.A(_04814_),
    .B(_04822_),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_1 _28510_ (.A(_04553_),
    .B(_04529_),
    .Y(_04824_));
 sky130_fd_sc_hd__nand3_1 _28511_ (.A(_04574_),
    .B(_04766_),
    .C(_04556_),
    .Y(_04825_));
 sky130_fd_sc_hd__nand2_1 _28512_ (.A(_04824_),
    .B(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__nand2_1 _28513_ (.A(_04357_),
    .B(net199),
    .Y(_04827_));
 sky130_fd_sc_hd__nand3_1 _28514_ (.A(_04502_),
    .B(_04766_),
    .C(_04484_),
    .Y(_04829_));
 sky130_fd_sc_hd__nand2_1 _28515_ (.A(_04827_),
    .B(_04829_),
    .Y(_04830_));
 sky130_fd_sc_hd__nor2_1 _28516_ (.A(_04826_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__nand2_1 _28517_ (.A(_04329_),
    .B(_04303_),
    .Y(_04832_));
 sky130_fd_sc_hd__nand3_1 _28518_ (.A(_04326_),
    .B(_04766_),
    .C(_04304_),
    .Y(_04833_));
 sky130_fd_sc_hd__nand2_1 _28519_ (.A(_04832_),
    .B(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__nand2_1 _28520_ (.A(_04576_),
    .B(_04555_),
    .Y(_04835_));
 sky130_fd_sc_hd__nand3_1 _28521_ (.A(_04597_),
    .B(_04766_),
    .C(_04578_),
    .Y(_04836_));
 sky130_fd_sc_hd__nand2_1 _28522_ (.A(_04835_),
    .B(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__nor2_1 _28523_ (.A(_04834_),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__nand2_1 _28524_ (.A(_04831_),
    .B(_04838_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_1 _28525_ (.A(_04823_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__nor3_1 _28526_ (.A(_04222_),
    .B(_04252_),
    .C(_04272_),
    .Y(_04842_));
 sky130_fd_sc_hd__nand3_1 _28527_ (.A(_04272_),
    .B(_04276_),
    .C(_04252_),
    .Y(_04843_));
 sky130_fd_sc_hd__nand3b_1 _28528_ (.A_N(_04300_),
    .B(_04276_),
    .C(_04281_),
    .Y(_04844_));
 sky130_fd_sc_hd__nand2_1 _28529_ (.A(_04843_),
    .B(_04844_),
    .Y(_04845_));
 sky130_fd_sc_hd__nor2_1 _28530_ (.A(_04842_),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2_1 _28531_ (.A(_04246_),
    .B(_04205_),
    .Y(_04847_));
 sky130_fd_sc_hd__o21ai_1 _28532_ (.A1(_04205_),
    .A2(_04247_),
    .B1(_04847_),
    .Y(_04848_));
 sky130_fd_sc_hd__nand3_1 _28533_ (.A(_04848_),
    .B(_04275_),
    .C(net175),
    .Y(_04849_));
 sky130_fd_sc_hd__inv_2 _28534_ (.A(_04849_),
    .Y(_04851_));
 sky130_fd_sc_hd__nand3_1 _28535_ (.A(_04249_),
    .B(_04276_),
    .C(_04228_),
    .Y(_04852_));
 sky130_fd_sc_hd__nand3_1 _28536_ (.A(_04300_),
    .B(_04276_),
    .C(net184),
    .Y(_04853_));
 sky130_fd_sc_hd__nand2_1 _28537_ (.A(_04852_),
    .B(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__nand2_1 _28538_ (.A(_04504_),
    .B(_04483_),
    .Y(_04855_));
 sky130_fd_sc_hd__nand2_1 _28539_ (.A(_04527_),
    .B(_04506_),
    .Y(_04856_));
 sky130_fd_sc_hd__nand3_1 _28540_ (.A(_04525_),
    .B(_04276_),
    .C(_04507_),
    .Y(_04857_));
 sky130_fd_sc_hd__nand3_1 _28541_ (.A(_04855_),
    .B(_04856_),
    .C(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__nor3_2 _28542_ (.A(_04851_),
    .B(_04854_),
    .C(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__nand3_2 _28543_ (.A(_04841_),
    .B(_04846_),
    .C(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__nor2_1 _28544_ (.A(_04807_),
    .B(_04860_),
    .Y(_04862_));
 sky130_fd_sc_hd__nor2_1 _28545_ (.A(_02134_),
    .B(_04862_),
    .Y(_00001_));
 sky130_fd_sc_hd__nand2_1 _28546_ (.A(_02134_),
    .B(net142),
    .Y(_04863_));
 sky130_fd_sc_hd__inv_2 _28547_ (.A(net143),
    .Y(_00000_));
 sky130_fd_sc_hd__nand2_1 _28548_ (.A(_02134_),
    .B(net145),
    .Y(_04864_));
 sky130_fd_sc_hd__inv_2 _28549_ (.A(net146),
    .Y(_00002_));
 sky130_fd_sc_hd__or3b_1 _28550_ (.A(_02651_),
    .B(_02756_),
    .C_N(_02867_),
    .X(_04865_));
 sky130_fd_sc_hd__or3_1 _28551_ (.A(_02966_),
    .B(_04865_),
    .C(_03087_),
    .X(_04866_));
 sky130_fd_sc_hd__inv_2 _28552_ (.A(_03286_),
    .Y(_04867_));
 sky130_fd_sc_hd__and4b_1 _28553_ (.A_N(_04866_),
    .B(_04867_),
    .C(_03325_),
    .D(_03188_),
    .X(_04868_));
 sky130_fd_sc_hd__o21a_1 _28554_ (.A1(_03296_),
    .A2(_04868_),
    .B1(_02653_),
    .X(_00036_));
 sky130_fd_sc_hd__nand2_1 _28555_ (.A(_02756_),
    .B(_02651_),
    .Y(_04870_));
 sky130_fd_sc_hd__or3b_1 _28556_ (.A(_02867_),
    .B(_04870_),
    .C_N(_02966_),
    .X(_04871_));
 sky130_fd_sc_hd__or3b_1 _28557_ (.A(_04871_),
    .B(_03188_),
    .C_N(_03087_),
    .X(_04872_));
 sky130_fd_sc_hd__or3_1 _28558_ (.A(_04872_),
    .B(_03325_),
    .C(_04867_),
    .X(_04873_));
 sky130_fd_sc_hd__or3b_1 _28559_ (.A(_02774_),
    .B(_02885_),
    .C_N(_02673_),
    .X(_04874_));
 sky130_fd_sc_hd__or3_1 _28560_ (.A(_02990_),
    .B(_03106_),
    .C(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__or3_4 _28561_ (.A(_03206_),
    .B(_03294_),
    .C(_04875_),
    .X(_04876_));
 sky130_fd_sc_hd__a21oi_1 _28562_ (.A1(_04873_),
    .A2(_04876_),
    .B1(_02134_),
    .Y(_00035_));
 sky130_fd_sc_hd__inv_2 _28563_ (.A(net57),
    .Y(_04877_));
 sky130_fd_sc_hd__nand2_1 _28564_ (.A(net54),
    .B(net53),
    .Y(_04879_));
 sky130_fd_sc_hd__inv_2 _28565_ (.A(net48),
    .Y(_04880_));
 sky130_fd_sc_hd__nand2_1 _28566_ (.A(net52),
    .B(net51),
    .Y(_04881_));
 sky130_fd_sc_hd__nand2_1 _28567_ (.A(net50),
    .B(net49),
    .Y(_04882_));
 sky130_fd_sc_hd__or2_1 _28568_ (.A(_04881_),
    .B(_04882_),
    .X(_04883_));
 sky130_fd_sc_hd__or4_4 _28569_ (.A(_11935_),
    .B(_08554_),
    .C(_12495_),
    .D(_09943_),
    .X(_04884_));
 sky130_fd_sc_hd__or4_1 _28570_ (.A(_04880_),
    .B(_03287_),
    .C(_04883_),
    .D(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__or4_1 _28571_ (.A(_04877_),
    .B(_05386_),
    .C(_04879_),
    .D(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__or4_2 _28572_ (.A(net57),
    .B(_05386_),
    .C(_04879_),
    .D(_04885_),
    .X(_04887_));
 sky130_fd_sc_hd__nand2_1 _28573_ (.A(_02569_),
    .B(_03288_),
    .Y(_04888_));
 sky130_fd_sc_hd__or4_1 _28574_ (.A(net20),
    .B(net19),
    .C(net18),
    .D(net17),
    .X(_04890_));
 sky130_fd_sc_hd__or4_1 _28575_ (.A(net22),
    .B(net21),
    .C(_04888_),
    .D(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__or4_1 _28576_ (.A(net11),
    .B(net10),
    .C(net9),
    .D(net8),
    .X(_04892_));
 sky130_fd_sc_hd__or4_1 _28577_ (.A(net26),
    .B(net1),
    .C(net12),
    .D(net23),
    .X(_04893_));
 sky130_fd_sc_hd__or4_1 _28578_ (.A(net27),
    .B(net30),
    .C(net29),
    .D(net28),
    .X(_04894_));
 sky130_fd_sc_hd__or4_1 _28579_ (.A(net3),
    .B(net2),
    .C(net32),
    .D(net31),
    .X(_04895_));
 sky130_fd_sc_hd__or4_1 _28580_ (.A(net7),
    .B(net6),
    .C(net5),
    .D(net4),
    .X(_04896_));
 sky130_fd_sc_hd__or4_4 _28581_ (.A(_04893_),
    .B(_04894_),
    .C(_04895_),
    .D(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__nor3_1 _28582_ (.A(net15),
    .B(net14),
    .C(net13),
    .Y(_04898_));
 sky130_fd_sc_hd__or4b_4 _28583_ (.A(_04891_),
    .B(_04892_),
    .C(_04897_),
    .D_N(_04898_),
    .X(_04899_));
 sky130_fd_sc_hd__and3_1 _28584_ (.A(_04886_),
    .B(_04887_),
    .C(_04899_),
    .X(_04901_));
 sky130_fd_sc_hd__or2_1 _28585_ (.A(net54),
    .B(net53),
    .X(_04902_));
 sky130_fd_sc_hd__or4_1 _28586_ (.A(net52),
    .B(net51),
    .C(net50),
    .D(net49),
    .X(_04903_));
 sky130_fd_sc_hd__or4_1 _28587_ (.A(net48),
    .B(net56),
    .C(_04903_),
    .D(_04884_),
    .X(_04904_));
 sky130_fd_sc_hd__or3_1 _28588_ (.A(net57),
    .B(_04902_),
    .C(_04904_),
    .X(_04905_));
 sky130_fd_sc_hd__nor2_1 _28589_ (.A(_05386_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__or4_1 _28590_ (.A(_04877_),
    .B(_05386_),
    .C(_04902_),
    .D(_04904_),
    .X(_04907_));
 sky130_fd_sc_hd__and2b_1 _28591_ (.A_N(_04906_),
    .B(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__nand2_1 _28592_ (.A(_04901_),
    .B(_04908_),
    .Y(_04909_));
 sky130_fd_sc_hd__inv_2 _28593_ (.A(_04909_),
    .Y(_04910_));
 sky130_fd_sc_hd__nand2_1 _28594_ (.A(_04886_),
    .B(_04887_),
    .Y(_04912_));
 sky130_fd_sc_hd__inv_2 _28595_ (.A(_04912_),
    .Y(_04913_));
 sky130_fd_sc_hd__or3b_1 _28596_ (.A(_02569_),
    .B(_04892_),
    .C_N(_04898_),
    .X(_04914_));
 sky130_fd_sc_hd__and4_1 _28597_ (.A(net24),
    .B(net22),
    .C(net18),
    .D(net17),
    .X(_04915_));
 sky130_fd_sc_hd__and3_1 _28598_ (.A(net21),
    .B(net20),
    .C(net19),
    .X(_04916_));
 sky130_fd_sc_hd__nand2_1 _28599_ (.A(_04915_),
    .B(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hd__or4_1 _28600_ (.A(_04897_),
    .B(_04914_),
    .C(_04917_),
    .D(_04913_),
    .X(_04918_));
 sky130_fd_sc_hd__o21a_1 _28601_ (.A1(_04899_),
    .A2(_04913_),
    .B1(_04918_),
    .X(_04919_));
 sky130_fd_sc_hd__o21ai_4 _28602_ (.A1(_04908_),
    .A2(_04899_),
    .B1(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__nor2_8 _28603_ (.A(_04910_),
    .B(_04920_),
    .Y(div_zero_f_c));
 sky130_fd_sc_hd__inv_2 _28604_ (.A(div_zero_f_c),
    .Y(\out_f_c[22] ));
 sky130_fd_sc_hd__or2_1 _28605_ (.A(_04901_),
    .B(_04920_),
    .X(_04922_));
 sky130_fd_sc_hd__buf_4 _28606_ (.A(_04922_),
    .X(\out_f_c[23] ));
 sky130_fd_sc_hd__a21boi_1 _28607_ (.A1(_04907_),
    .A2(_04886_),
    .B1_N(_04887_),
    .Y(_04923_));
 sky130_fd_sc_hd__nand3b_1 _28608_ (.A_N(_04906_),
    .B(_04887_),
    .C(net25),
    .Y(_04924_));
 sky130_fd_sc_hd__o2111a_4 _28609_ (.A1(net25),
    .A2(_04923_),
    .B1(_04899_),
    .C1(_04924_),
    .D1(_04918_),
    .X(\out_f_c[31] ));
 sky130_fd_sc_hd__or4_4 _28610_ (.A(net25),
    .B(_04897_),
    .C(_04917_),
    .D(_04914_),
    .X(_04925_));
 sky130_fd_sc_hd__nand2_8 _28611_ (.A(_04910_),
    .B(_04925_),
    .Y(forward_c));
 sky130_fd_sc_hd__inv_2 _28612_ (.A(div_zero_f_c),
    .Y(inv_f_c));
 sky130_fd_sc_hd__dfrtp_1 _28613_ (.CLK(clknet_3_1_0_clk),
    .D(\div1i.quot[0] ),
    .RESET_B(net115),
    .Q(\M00r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _28614_ (.CLK(clknet_3_0_0_clk),
    .D(\div1i.quot[1] ),
    .RESET_B(net115),
    .Q(\M00r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _28615_ (.CLK(clknet_3_0_0_clk),
    .D(\div1i.quot[2] ),
    .RESET_B(net116),
    .Q(\M00r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _28616_ (.CLK(clknet_3_1_0_clk),
    .D(\div1i.quot[3] ),
    .RESET_B(net116),
    .Q(\M00r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _28617_ (.CLK(clknet_3_1_0_clk),
    .D(\div1i.quot[4] ),
    .RESET_B(net116),
    .Q(\M00r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _28618_ (.CLK(clknet_3_0_0_clk),
    .D(\div1i.quot[5] ),
    .RESET_B(net116),
    .Q(\M00r[5] ));
 sky130_fd_sc_hd__dfrtp_1 _28619_ (.CLK(clknet_3_1_0_clk),
    .D(\div1i.quot[6] ),
    .RESET_B(net116),
    .Q(\M00r[6] ));
 sky130_fd_sc_hd__dfrtp_1 _28620_ (.CLK(clknet_3_0_0_clk),
    .D(\div1i.quot[7] ),
    .RESET_B(net116),
    .Q(\M00r[7] ));
 sky130_fd_sc_hd__dfrtp_1 _28621_ (.CLK(clknet_3_0_0_clk),
    .D(\div1i.quot[8] ),
    .RESET_B(net116),
    .Q(\M00r[8] ));
 sky130_fd_sc_hd__dfrtp_1 _28622_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[9] ),
    .RESET_B(net108),
    .Q(\M00r[9] ));
 sky130_fd_sc_hd__dfrtp_1 _28623_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[10] ),
    .RESET_B(net108),
    .Q(\M00r[10] ));
 sky130_fd_sc_hd__dfrtp_1 _28624_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[11] ),
    .RESET_B(net108),
    .Q(\M00r[11] ));
 sky130_fd_sc_hd__dfrtp_1 _28625_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[12] ),
    .RESET_B(net108),
    .Q(\M00r[12] ));
 sky130_fd_sc_hd__dfrtp_1 _28626_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[13] ),
    .RESET_B(net108),
    .Q(\M00r[13] ));
 sky130_fd_sc_hd__dfrtp_1 _28627_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[14] ),
    .RESET_B(net108),
    .Q(\M00r[14] ));
 sky130_fd_sc_hd__dfrtp_1 _28628_ (.CLK(clknet_3_3_0_clk),
    .D(net222),
    .RESET_B(net108),
    .Q(\M00r[15] ));
 sky130_fd_sc_hd__dfrtp_1 _28629_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[16] ),
    .RESET_B(net108),
    .Q(\M00r[16] ));
 sky130_fd_sc_hd__dfrtp_1 _28630_ (.CLK(clknet_3_3_0_clk),
    .D(\div1i.quot[17] ),
    .RESET_B(net108),
    .Q(\M00r[17] ));
 sky130_fd_sc_hd__dfrtp_2 _28631_ (.CLK(clknet_3_2_0_clk),
    .D(\div1i.quot[18] ),
    .RESET_B(net109),
    .Q(\M00r[18] ));
 sky130_fd_sc_hd__dfrtp_1 _28632_ (.CLK(clknet_3_2_0_clk),
    .D(\div1i.quot[19] ),
    .RESET_B(net109),
    .Q(\M00r[19] ));
 sky130_fd_sc_hd__dfrtp_2 _28633_ (.CLK(clknet_3_2_0_clk),
    .D(\div1i.quot[20] ),
    .RESET_B(net109),
    .Q(\M00r[20] ));
 sky130_fd_sc_hd__dfrtp_4 _28634_ (.CLK(clknet_3_2_0_clk),
    .D(\div1i.quot[21] ),
    .RESET_B(net109),
    .Q(\M00r[21] ));
 sky130_fd_sc_hd__dfrtp_1 _28635_ (.CLK(clknet_3_2_0_clk),
    .D(\div1i.quot[22] ),
    .RESET_B(net109),
    .Q(\M00r[22] ));
 sky130_fd_sc_hd__dfrtp_1 _28636_ (.CLK(clknet_3_2_0_clk),
    .D(\div1i.quot[23] ),
    .RESET_B(net109),
    .Q(\M00r[23] ));
 sky130_fd_sc_hd__dfrtp_1 _28637_ (.CLK(clknet_3_2_0_clk),
    .D(net118),
    .RESET_B(net108),
    .Q(\M00r[24] ));
 sky130_fd_sc_hd__conb_1 _28637__118 (.HI(net118));
 sky130_fd_sc_hd__dfrtp_2 _28638_ (.CLK(clknet_3_5_0_clk),
    .D(_00003_),
    .RESET_B(net110),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_2 _28639_ (.CLK(clknet_3_5_0_clk),
    .D(_00014_),
    .RESET_B(net115),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_2 _28640_ (.CLK(clknet_3_5_0_clk),
    .D(_00025_),
    .RESET_B(net110),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_2 _28641_ (.CLK(clknet_3_4_0_clk),
    .D(_00028_),
    .RESET_B(net111),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _28642_ (.CLK(clknet_3_5_0_clk),
    .D(_00029_),
    .RESET_B(net110),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_2 _28643_ (.CLK(clknet_3_5_0_clk),
    .D(_00030_),
    .RESET_B(net111),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_2 _28644_ (.CLK(clknet_3_4_0_clk),
    .D(_00031_),
    .RESET_B(net111),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_2 _28645_ (.CLK(clknet_3_4_0_clk),
    .D(_00032_),
    .RESET_B(net111),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _28646_ (.CLK(clknet_3_4_0_clk),
    .D(_00033_),
    .RESET_B(net111),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _28647_ (.CLK(clknet_3_5_0_clk),
    .D(_00034_),
    .RESET_B(net110),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _28648_ (.CLK(clknet_3_4_0_clk),
    .D(_00004_),
    .RESET_B(net110),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _28649_ (.CLK(clknet_3_5_0_clk),
    .D(_00005_),
    .RESET_B(net110),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _28650_ (.CLK(clknet_3_4_0_clk),
    .D(_00006_),
    .RESET_B(net110),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _28651_ (.CLK(clknet_3_5_0_clk),
    .D(_00007_),
    .RESET_B(net111),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _28652_ (.CLK(clknet_3_5_0_clk),
    .D(_00008_),
    .RESET_B(net111),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _28653_ (.CLK(clknet_3_4_0_clk),
    .D(_00009_),
    .RESET_B(net111),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _28654_ (.CLK(clknet_3_6_0_clk),
    .D(_00010_),
    .RESET_B(net113),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _28655_ (.CLK(clknet_3_6_0_clk),
    .D(_00011_),
    .RESET_B(net113),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _28656_ (.CLK(clknet_3_6_0_clk),
    .D(_00012_),
    .RESET_B(net113),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _28657_ (.CLK(clknet_3_5_0_clk),
    .D(_00013_),
    .RESET_B(net110),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _28658_ (.CLK(clknet_3_5_0_clk),
    .D(_00015_),
    .RESET_B(net110),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _28659_ (.CLK(clknet_3_5_0_clk),
    .D(_00016_),
    .RESET_B(net110),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _28660_ (.CLK(clknet_3_7_0_clk),
    .D(_00017_),
    .RESET_B(net113),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _28661_ (.CLK(clknet_3_6_0_clk),
    .D(_00018_),
    .RESET_B(net113),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _28662_ (.CLK(clknet_3_4_0_clk),
    .D(_00019_),
    .RESET_B(net111),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _28663_ (.CLK(clknet_3_6_0_clk),
    .D(net162),
    .RESET_B(net113),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _28664_ (.CLK(clknet_3_4_0_clk),
    .D(_00021_),
    .RESET_B(net115),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _28665_ (.CLK(clknet_3_6_0_clk),
    .D(_00022_),
    .RESET_B(net113),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _28666_ (.CLK(clknet_3_7_0_clk),
    .D(net158),
    .RESET_B(net112),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _28667_ (.CLK(clknet_3_7_0_clk),
    .D(net165),
    .RESET_B(net112),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _28668_ (.CLK(clknet_3_7_0_clk),
    .D(net155),
    .RESET_B(net112),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _28669_ (.CLK(clknet_3_6_0_clk),
    .D(net152),
    .RESET_B(net113),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _28670_ (.CLK(clknet_3_7_0_clk),
    .D(_00035_),
    .RESET_B(net112),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_1 _28671_ (.CLK(clknet_3_7_0_clk),
    .D(_00036_),
    .RESET_B(net114),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_1 _28672_ (.CLK(clknet_3_7_0_clk),
    .D(net216),
    .RESET_B(net112),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _28673_ (.CLK(clknet_3_7_0_clk),
    .D(net147),
    .RESET_B(net112),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _28674_ (.CLK(clknet_3_7_0_clk),
    .D(net144),
    .RESET_B(net113),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _28675_ (.CLK(clknet_3_7_0_clk),
    .D(_00001_),
    .RESET_B(net113),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _28676_ (.CLK(clknet_3_6_0_clk),
    .D(net117),
    .RESET_B(net112),
    .Q(done0_reg));
 sky130_fd_sc_hd__conb_1 _28676__117 (.HI(net117));
 sky130_fd_sc_hd__dfrtp_1 _28677_ (.CLK(clknet_3_7_0_clk),
    .D(\out_f_c[22] ),
    .RESET_B(net112),
    .Q(\out_f[22] ));
 sky130_fd_sc_hd__dfrtp_1 _28678_ (.CLK(clknet_3_1_0_clk),
    .D(\out_f_c[23] ),
    .RESET_B(net114),
    .Q(\out_f[23] ));
 sky130_fd_sc_hd__dfrtp_1 _28679_ (.CLK(clknet_3_1_0_clk),
    .D(\out_f_c[31] ),
    .RESET_B(net114),
    .Q(\out_f[31] ));
 sky130_fd_sc_hd__dfrtp_1 _28680_ (.CLK(clknet_3_7_0_clk),
    .D(inv_f_c),
    .RESET_B(net112),
    .Q(inv_f));
 sky130_fd_sc_hd__dfrtp_1 _28681_ (.CLK(clknet_3_6_0_clk),
    .D(div_zero_f_c),
    .RESET_B(net112),
    .Q(div_zero_f));
 sky130_fd_sc_hd__dfrtp_1 _28682_ (.CLK(clknet_3_1_0_clk),
    .D(forward_c),
    .RESET_B(net114),
    .Q(forward));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(net68),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net115),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(net114),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 fanout116 (.A(net68),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_02440_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\out_f[22] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(done0_reg),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net215),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(div_zero_f),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_04863_),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_00000_),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(inv_f),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_04864_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_00002_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net219),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_04760_),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\out_f[31] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_02136_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_00027_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net166),
    .X(net153));
 sky130_fd_sc_hd__buf_1 hold36 (.A(_02654_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_00026_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 hold38 (.A(net164),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_00023_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net163),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_4 hold42 (.A(net156),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_00020_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(forward),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net159),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_00024_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\out_f[23] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\M00r[0] ),
    .X(net167));
 sky130_fd_sc_hd__buf_4 hold50 (.A(net186),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 hold51 (.A(_04268_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_04269_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\M00r[2] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_02441_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_02520_),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_04226_),
    .X(net174));
 sky130_fd_sc_hd__buf_2 hold57 (.A(_04227_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_04228_),
    .X(net176));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold59 (.A(\M00r[22] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_02140_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_02147_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_02148_),
    .X(net180));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold63 (.A(_02150_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_02151_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_02156_),
    .X(net183));
 sky130_fd_sc_hd__buf_2 hold66 (.A(_04280_),
    .X(net184));
 sky130_fd_sc_hd__buf_2 hold67 (.A(\M00r[24] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_04161_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\M00r[1] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_02518_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_02519_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_2 hold72 (.A(_04198_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\M00r[5] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_02368_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_02446_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_02447_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_02448_),
    .X(net195));
 sky130_fd_sc_hd__buf_1 hold78 (.A(_02526_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_02528_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_02529_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 hold81 (.A(_04332_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 hold82 (.A(\M00r[23] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\M00r[19] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_02161_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_02167_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_02172_),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_02174_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\M00r[7] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_02371_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_02372_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_02374_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_02453_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_02454_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_02455_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_02533_),
    .X(net213));
 sky130_fd_sc_hd__buf_1 hold96 (.A(\M00r[21] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net220),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net141),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\M00r[3] ),
    .X(net217));
 sky130_fd_sc_hd__buf_2 input1 (.A(in1[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(in1[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(in1[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in1[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(in1[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(in1[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(in1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in1[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(in1[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(in1[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(in1[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(in1[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in1[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in1[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in1[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(in1[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(in1[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(in1[3]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(in1[4]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(in1[5]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(in1[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(in1[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(in1[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in1[8]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(in1[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_4 input33 (.A(in2[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(in2[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_4 input35 (.A(in2[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_6 input36 (.A(in2[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(in2[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_6 input38 (.A(in2[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(in2[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(in1[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input40 (.A(in2[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_4 input41 (.A(in2[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(in2[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 input43 (.A(in2[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 input44 (.A(in2[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(in2[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(in2[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(in2[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in2[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(in2[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(in1[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(in2[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(in2[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(in2[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(in2[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(in2[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_4 input55 (.A(in2[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(in2[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_2 input57 (.A(in2[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input58 (.A(in2[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 input59 (.A(in2[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(in1[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(in2[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(in2[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(in2[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_4 input63 (.A(in2[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(in2[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_8 input65 (.A(round_m[0]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 input66 (.A(round_m[1]),
    .X(net66));
 sky130_fd_sc_hd__buf_4 input67 (.A(round_m[2]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 input68 (.A(rst),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input7 (.A(in1[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(in1[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(in1[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(out[5]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(out[6]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(out[7]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(out[8]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(out[9]));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(ov));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(un));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(div_zero));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(done));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(inexact));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(inv));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(out[0]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(out[10]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(out[11]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(out[12]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(out[13]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(out[14]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(out[15]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(out[16]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(out[17]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(out[18]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(out[19]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(out[20]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(out[21]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(out[22]));
 sky130_fd_sc_hd__clkbuf_4 output88 (.A(net88),
    .X(out[23]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(out[24]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(out[25]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(out[26]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(out[27]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(out[28]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(out[29]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(out[2]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(out[30]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(out[31]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(out[3]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(out[4]));
 sky130_fd_sc_hd__clkbuf_2 rebuffer10 (.A(_06383_),
    .X(net128));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer11 (.A(_07538_),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 rebuffer12 (.A(_06383_),
    .X(net130));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer13 (.A(_07007_),
    .X(net136));
 sky130_fd_sc_hd__buf_6 rebuffer16 (.A(_06385_),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer17 (.A(_06269_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer18 (.A(_06951_),
    .X(net140));
 sky130_fd_sc_hd__buf_6 rebuffer20 (.A(_06971_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_2 rebuffer31 (.A(_06387_),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 rebuffer37 (.A(_06624_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 rebuffer40 (.A(_06860_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer41 (.A(_10009_),
    .X(net241));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer44 (.A(_05927_),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 rebuffer5 (.A(_06969_),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 rebuffer6 (.A(_06969_),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 rebuffer7 (.A(_06969_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 rebuffer8 (.A(_06969_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 rebuffer9 (.A(_06969_),
    .X(net127));
 sky130_fd_sc_hd__buf_6 split1 (.A(_01588_),
    .X(net119));
 sky130_fd_sc_hd__buf_6 split11 (.A(_01586_),
    .X(net129));
 sky130_fd_sc_hd__buf_4 split13 (.A(_04237_),
    .X(net131));
 sky130_fd_sc_hd__buf_6 split14 (.A(_02112_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 split15 (.A(_08582_),
    .X(net137));
 sky130_fd_sc_hd__buf_6 split19 (.A(_06972_),
    .X(net157));
 sky130_fd_sc_hd__buf_2 split2 (.A(_09724_),
    .X(net120));
 sky130_fd_sc_hd__buf_6 split21 (.A(_08101_),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 split22 (.A(\div1i.quot[15] ),
    .X(net222));
 sky130_fd_sc_hd__buf_6 split23 (.A(_12555_),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 split24 (.A(_09743_),
    .X(net224));
 sky130_fd_sc_hd__buf_6 split25 (.A(_10300_),
    .X(net225));
 sky130_fd_sc_hd__buf_6 split26 (.A(_13664_),
    .X(net226));
 sky130_fd_sc_hd__buf_6 split27 (.A(_11397_),
    .X(net227));
 sky130_fd_sc_hd__buf_6 split28 (.A(_00502_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 split29 (.A(_08644_),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 split3 (.A(_08571_),
    .X(net121));
 sky130_fd_sc_hd__buf_6 split30 (.A(_13104_),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_2 split32 (.A(_14202_),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 split33 (.A(_01590_),
    .X(net233));
 sky130_fd_sc_hd__buf_6 split34 (.A(_05010_),
    .X(net234));
 sky130_fd_sc_hd__buf_6 split35 (.A(_05834_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 split36 (.A(_13102_),
    .X(net236));
 sky130_fd_sc_hd__buf_6 split38 (.A(_09200_),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 split39 (.A(_02132_),
    .X(net239));
 sky130_fd_sc_hd__buf_6 split4 (.A(_02131_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 split42 (.A(_11971_),
    .X(net242));
 sky130_fd_sc_hd__buf_2 split43 (.A(_07055_),
    .X(net243));
 sky130_fd_sc_hd__buf_6 split5 (.A(_12974_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_2 split6 (.A(_07011_),
    .X(net134));
 sky130_fd_sc_hd__buf_4 wire107 (.A(_02135_),
    .X(net107));
endmodule

