// This is the unpowered netlist.
module fp_add (clk,
    done,
    inexact,
    inv,
    ov,
    rst,
    un,
    in1,
    in2,
    out,
    round_m);
 input clk;
 output done;
 output inexact;
 output inv;
 output ov;
 input rst;
 output un;
 input [31:0] in1;
 input [31:0] in2;
 output [31:0] out;
 input [2:0] round_m;

 wire \M000[0] ;
 wire \M000[10] ;
 wire \M000[11] ;
 wire \M000[12] ;
 wire \M000[13] ;
 wire \M000[14] ;
 wire \M000[15] ;
 wire \M000[16] ;
 wire \M000[17] ;
 wire \M000[18] ;
 wire \M000[19] ;
 wire \M000[1] ;
 wire \M000[20] ;
 wire \M000[21] ;
 wire \M000[22] ;
 wire \M000[23] ;
 wire \M000[24] ;
 wire \M000[25] ;
 wire \M000[26] ;
 wire \M000[2] ;
 wire \M000[3] ;
 wire \M000[4] ;
 wire \M000[5] ;
 wire \M000[6] ;
 wire \M000[7] ;
 wire \M000[8] ;
 wire \M000[9] ;
 wire \M00[0] ;
 wire \M00[10] ;
 wire \M00[11] ;
 wire \M00[12] ;
 wire \M00[13] ;
 wire \M00[14] ;
 wire \M00[15] ;
 wire \M00[16] ;
 wire \M00[17] ;
 wire \M00[18] ;
 wire \M00[19] ;
 wire \M00[1] ;
 wire \M00[20] ;
 wire \M00[21] ;
 wire \M00[22] ;
 wire \M00[23] ;
 wire \M00[24] ;
 wire \M00[25] ;
 wire \M00[26] ;
 wire \M00[2] ;
 wire \M00[3] ;
 wire \M00[4] ;
 wire \M00[5] ;
 wire \M00[6] ;
 wire \M00[7] ;
 wire \M00[8] ;
 wire \M00[9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire done0_r;
 wire forward;
 wire forward_c;
 wire inv_f;
 wire inv_f_c;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \out_f[31] ;
 wire \out_f_c[31] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__S (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__C (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__B (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__B (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A0 (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__B1 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__S (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A (.DIODE(_2739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__B_N (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__S (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A2 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__S (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__S (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__S (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__S (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A1 (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A1 (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__B1 (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A2 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A1 (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A1 (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A1 (.DIODE(_1630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3735__S (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__C1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A2 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__C (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__S (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__S (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3852__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3854__S (.DIODE(_1124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A2 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B (.DIODE(_2329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3865__A1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3898__C (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__S (.DIODE(_2809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A1 (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__S (.DIODE(_1729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4173__A (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__A (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A (.DIODE(_0074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__A (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A2 (.DIODE(_2717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A3 (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__B1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__C (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__C (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__B (.DIODE(_0089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__C (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__A (.DIODE(_0089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__B (.DIODE(_0095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__A (.DIODE(_0089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4217__A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__A1 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A (.DIODE(_0095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__B (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__B (.DIODE(_0089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__A (.DIODE(_0089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__C (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__S (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__B (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__B_N (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__S (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__C (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__S (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__C (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__C (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B_N (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__S (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__C (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__C (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__S (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__S (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__C (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__C (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__C (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__S (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__C (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__C (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__C (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__B (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__C (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A1 (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__B (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__S (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A2 (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__B (.DIODE(_0960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__B (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__C (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__B (.DIODE(_0491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__B (.DIODE(_1767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__B (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__B1 (.DIODE(_1041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__B1 (.DIODE(_1199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__S (.DIODE(_1674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__B (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__B (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__B (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A1 (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A2 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__B1 (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A (.DIODE(_1968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__C (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A2 (.DIODE(_2072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(_1823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__B (.DIODE(_0095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A (.DIODE(_0089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A2 (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A3 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__S (.DIODE(_0074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A1 (.DIODE(_2740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A (.DIODE(_1767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__B1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A1 (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A3 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A1 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A2 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__C1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__B1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A1 (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A2 (.DIODE(_2034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__B (.DIODE(_0078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__B1 (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__C1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__S (.DIODE(_0074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__S (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__B1 (.DIODE(_0067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A3 (.DIODE(_1696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A2 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A2 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A3 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__A2 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__A2 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A2 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__S (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A1_N (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A2_N (.DIODE(_2308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__B (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A2_N (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__B2 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__S (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__A (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A2 (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A2 (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A2 (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A2_N (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__B (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A1 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__B1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__B (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__B (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A2 (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__B (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A2 (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A2 (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A1 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__B (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A2 (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A1_N (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__B1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__B (.DIODE(_2305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A1 (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__A1 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__B1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__B (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A1_N (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__B (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__B (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__B (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__B1 (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__B (.DIODE(_0058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__B (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__B (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A1 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__B1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__B (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A1 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__B1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__B (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__B (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__B1 (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A2 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B1 (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A1_N (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__B (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__B1 (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A2 (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A2 (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B1 (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__B (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A2 (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B (.DIODE(_2306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A2 (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A2 (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__B (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A1 (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A (.DIODE(_2331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A (.DIODE(_2325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__B1 (.DIODE(_2328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A2 (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__B2 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A1 (.DIODE(_2345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A (.DIODE(_2337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__D (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__RESET_B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold10_A (.DIODE(_0026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold64_A (.DIODE(_1770_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold66_A (.DIODE(_1760_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__buf_6 _3313_ (.A(net157),
    .X(_0684_));
 sky130_fd_sc_hd__buf_4 _3314_ (.A(_0684_),
    .X(_0695_));
 sky130_fd_sc_hd__clkbuf_4 _3315_ (.A(_0695_),
    .X(_0706_));
 sky130_fd_sc_hd__mux2_1 _3316_ (.A0(\M000[1] ),
    .A1(net135),
    .S(_0706_),
    .X(_0717_));
 sky130_fd_sc_hd__inv_2 _3317_ (.A(\M000[1] ),
    .Y(_0728_));
 sky130_fd_sc_hd__nand2_1 _3318_ (.A(_0728_),
    .B(_0706_),
    .Y(_0739_));
 sky130_fd_sc_hd__o21a_1 _3319_ (.A1(_0706_),
    .A2(net128),
    .B1(_0739_),
    .X(_0750_));
 sky130_fd_sc_hd__nor2_4 _3320_ (.A(_0684_),
    .B(net179),
    .Y(_0761_));
 sky130_fd_sc_hd__buf_2 _3321_ (.A(_0761_),
    .X(_0772_));
 sky130_fd_sc_hd__clkbuf_4 _3322_ (.A(_0772_),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _3323_ (.A0(net136),
    .A1(net129),
    .S(_0783_),
    .X(_0794_));
 sky130_fd_sc_hd__inv_2 _3324_ (.A(net157),
    .Y(_0805_));
 sky130_fd_sc_hd__inv_2 _3325_ (.A(\M000[25] ),
    .Y(_0816_));
 sky130_fd_sc_hd__inv_2 _3326_ (.A(net144),
    .Y(_0827_));
 sky130_fd_sc_hd__and3_1 _3327_ (.A(_0805_),
    .B(_0816_),
    .C(_0827_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_2 _3328_ (.A(net158),
    .X(_0849_));
 sky130_fd_sc_hd__inv_2 _3329_ (.A(_0849_),
    .Y(_0860_));
 sky130_fd_sc_hd__clkbuf_4 _3330_ (.A(_0860_),
    .X(_0871_));
 sky130_fd_sc_hd__nand2_1 _3331_ (.A(net137),
    .B(_0871_),
    .Y(_0882_));
 sky130_fd_sc_hd__inv_2 _3332_ (.A(net138),
    .Y(_0893_));
 sky130_fd_sc_hd__inv_2 _3333_ (.A(net19),
    .Y(_0904_));
 sky130_fd_sc_hd__nand2_1 _3334_ (.A(_0904_),
    .B(net51),
    .Y(_0915_));
 sky130_fd_sc_hd__inv_2 _3335_ (.A(net51),
    .Y(_0926_));
 sky130_fd_sc_hd__nand2_1 _3336_ (.A(_0926_),
    .B(net19),
    .Y(_0937_));
 sky130_fd_sc_hd__nand2_1 _3337_ (.A(_0915_),
    .B(_0937_),
    .Y(_0948_));
 sky130_fd_sc_hd__inv_2 _3338_ (.A(_0948_),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_2 _3339_ (.A(net49),
    .Y(_0970_));
 sky130_fd_sc_hd__nand2_1 _3340_ (.A(_0970_),
    .B(net17),
    .Y(_0981_));
 sky130_fd_sc_hd__inv_2 _3341_ (.A(net17),
    .Y(_0992_));
 sky130_fd_sc_hd__nand2_1 _3342_ (.A(_0992_),
    .B(net49),
    .Y(_1003_));
 sky130_fd_sc_hd__inv_2 _3343_ (.A(net48),
    .Y(_1014_));
 sky130_fd_sc_hd__nand2_1 _3344_ (.A(_1014_),
    .B(net16),
    .Y(_1025_));
 sky130_fd_sc_hd__nand3_1 _3345_ (.A(_0981_),
    .B(_1003_),
    .C(_1025_),
    .Y(_1036_));
 sky130_fd_sc_hd__nand2_2 _3346_ (.A(_1036_),
    .B(_1003_),
    .Y(_1047_));
 sky130_fd_sc_hd__inv_2 _3347_ (.A(net50),
    .Y(_1058_));
 sky130_fd_sc_hd__nand2_1 _3348_ (.A(_1058_),
    .B(net18),
    .Y(_1069_));
 sky130_fd_sc_hd__inv_2 _3349_ (.A(net18),
    .Y(_1080_));
 sky130_fd_sc_hd__nand2_1 _3350_ (.A(_1080_),
    .B(net50),
    .Y(_1091_));
 sky130_fd_sc_hd__inv_2 _3351_ (.A(_1091_),
    .Y(_1102_));
 sky130_fd_sc_hd__a21o_1 _3352_ (.A1(_1047_),
    .A2(_1069_),
    .B1(_1102_),
    .X(_1113_));
 sky130_fd_sc_hd__xor2_4 _3353_ (.A(_0959_),
    .B(_1113_),
    .X(_1124_));
 sky130_fd_sc_hd__clkbuf_4 _3354_ (.A(_1124_),
    .X(_1135_));
 sky130_fd_sc_hd__and2_1 _3355_ (.A(_0981_),
    .B(_1003_),
    .X(_1146_));
 sky130_fd_sc_hd__inv_2 _3356_ (.A(net16),
    .Y(_1157_));
 sky130_fd_sc_hd__nand2_1 _3357_ (.A(_1157_),
    .B(net48),
    .Y(_1168_));
 sky130_fd_sc_hd__nand2_1 _3358_ (.A(_1146_),
    .B(_1168_),
    .Y(_1179_));
 sky130_fd_sc_hd__nand2_1 _3359_ (.A(_1179_),
    .B(_0981_),
    .Y(_1190_));
 sky130_fd_sc_hd__nand2_1 _3360_ (.A(_1069_),
    .B(_1091_),
    .Y(_1201_));
 sky130_fd_sc_hd__inv_2 _3361_ (.A(_1201_),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _3362_ (.A(_1190_),
    .B(_1212_),
    .Y(_1223_));
 sky130_fd_sc_hd__nand2_2 _3363_ (.A(_1223_),
    .B(_1069_),
    .Y(_1234_));
 sky130_fd_sc_hd__xor2_4 _3364_ (.A(_0959_),
    .B(_1234_),
    .X(_1245_));
 sky130_fd_sc_hd__nor2_1 _3365_ (.A(_0948_),
    .B(_1201_),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _3366_ (.A(_1047_),
    .B(_1256_),
    .Y(_1267_));
 sky130_fd_sc_hd__a21boi_1 _3367_ (.A1(_1102_),
    .A2(_0937_),
    .B1_N(_0915_),
    .Y(_1278_));
 sky130_fd_sc_hd__nand2_2 _3368_ (.A(_1267_),
    .B(_1278_),
    .Y(_1289_));
 sky130_fd_sc_hd__inv_2 _3369_ (.A(net53),
    .Y(_1300_));
 sky130_fd_sc_hd__nand2_1 _3370_ (.A(_1300_),
    .B(net21),
    .Y(_1311_));
 sky130_fd_sc_hd__inv_2 _3371_ (.A(net21),
    .Y(_1322_));
 sky130_fd_sc_hd__nand2_1 _3372_ (.A(_1322_),
    .B(net53),
    .Y(_1333_));
 sky130_fd_sc_hd__nand2_2 _3373_ (.A(_1311_),
    .B(_1333_),
    .Y(_1344_));
 sky130_fd_sc_hd__inv_2 _3374_ (.A(net52),
    .Y(_1355_));
 sky130_fd_sc_hd__nand2_1 _3375_ (.A(_1355_),
    .B(net20),
    .Y(_1366_));
 sky130_fd_sc_hd__inv_2 _3376_ (.A(net20),
    .Y(_1377_));
 sky130_fd_sc_hd__nand2_1 _3377_ (.A(_1377_),
    .B(net52),
    .Y(_1388_));
 sky130_fd_sc_hd__nand2_1 _3378_ (.A(_1366_),
    .B(_1388_),
    .Y(_1399_));
 sky130_fd_sc_hd__nor2_1 _3379_ (.A(_1344_),
    .B(_1399_),
    .Y(_1410_));
 sky130_fd_sc_hd__inv_2 _3380_ (.A(net24),
    .Y(_1421_));
 sky130_fd_sc_hd__nand2_1 _3381_ (.A(_1421_),
    .B(net56),
    .Y(_1432_));
 sky130_fd_sc_hd__inv_2 _3382_ (.A(net56),
    .Y(_1443_));
 sky130_fd_sc_hd__nand2_1 _3383_ (.A(_1443_),
    .B(net24),
    .Y(_1454_));
 sky130_fd_sc_hd__nand2_1 _3384_ (.A(_1432_),
    .B(_1454_),
    .Y(_1465_));
 sky130_fd_sc_hd__inv_2 _3385_ (.A(net54),
    .Y(_1476_));
 sky130_fd_sc_hd__nand2_1 _3386_ (.A(_1476_),
    .B(net22),
    .Y(_1487_));
 sky130_fd_sc_hd__inv_2 _3387_ (.A(net22),
    .Y(_1498_));
 sky130_fd_sc_hd__nand2_1 _3388_ (.A(_1498_),
    .B(net54),
    .Y(_1509_));
 sky130_fd_sc_hd__nand2_1 _3389_ (.A(_1487_),
    .B(_1509_),
    .Y(_1520_));
 sky130_fd_sc_hd__nor2_1 _3390_ (.A(_1465_),
    .B(_1520_),
    .Y(_1531_));
 sky130_fd_sc_hd__and2_1 _3391_ (.A(_1410_),
    .B(_1531_),
    .X(_1542_));
 sky130_fd_sc_hd__nand2_1 _3392_ (.A(_1289_),
    .B(_1542_),
    .Y(_1553_));
 sky130_fd_sc_hd__inv_2 _3393_ (.A(_1311_),
    .Y(_1564_));
 sky130_fd_sc_hd__o21ai_1 _3394_ (.A1(_1388_),
    .A2(_1564_),
    .B1(_1333_),
    .Y(_1575_));
 sky130_fd_sc_hd__o21ai_1 _3395_ (.A1(_1509_),
    .A2(_1465_),
    .B1(_1432_),
    .Y(_1586_));
 sky130_fd_sc_hd__a21oi_1 _3396_ (.A1(_1575_),
    .A2(_1531_),
    .B1(_1586_),
    .Y(_1597_));
 sky130_fd_sc_hd__nand2_4 _3397_ (.A(_1553_),
    .B(_1597_),
    .Y(_1608_));
 sky130_fd_sc_hd__and2_1 _3398_ (.A(_1168_),
    .B(_1025_),
    .X(_1619_));
 sky130_fd_sc_hd__buf_4 _3399_ (.A(_1619_),
    .X(_1630_));
 sky130_fd_sc_hd__and3_1 _3400_ (.A(_1256_),
    .B(_1146_),
    .C(_1630_),
    .X(_1641_));
 sky130_fd_sc_hd__nand2_4 _3401_ (.A(_1641_),
    .B(_1542_),
    .Y(_1652_));
 sky130_fd_sc_hd__nand2_4 _3402_ (.A(_1608_),
    .B(_1652_),
    .Y(_1663_));
 sky130_fd_sc_hd__buf_4 _3403_ (.A(_1663_),
    .X(_1674_));
 sky130_fd_sc_hd__inv_2 _3404_ (.A(_1674_),
    .Y(_1685_));
 sky130_fd_sc_hd__inv_2 _3405_ (.A(net126),
    .Y(_1696_));
 sky130_fd_sc_hd__nand2_2 _3406_ (.A(_1685_),
    .B(_1696_),
    .Y(_1707_));
 sky130_fd_sc_hd__mux2_2 _3407_ (.A0(_1135_),
    .A1(_1245_),
    .S(_1707_),
    .X(_1718_));
 sky130_fd_sc_hd__xor2_4 _3408_ (.A(_1212_),
    .B(_1047_),
    .X(_1729_));
 sky130_fd_sc_hd__or2_1 _3409_ (.A(_1212_),
    .B(_1190_),
    .X(_1740_));
 sky130_fd_sc_hd__and2_1 _3410_ (.A(_1740_),
    .B(_1223_),
    .X(_1751_));
 sky130_fd_sc_hd__clkbuf_4 _3411_ (.A(_1751_),
    .X(_1762_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(_1729_),
    .A1(_1762_),
    .S(_1707_),
    .X(_1773_));
 sky130_fd_sc_hd__and3_1 _3413_ (.A(_1432_),
    .B(_1454_),
    .C(_1487_),
    .X(_1784_));
 sky130_fd_sc_hd__a21bo_1 _3414_ (.A1(_1234_),
    .A2(_0915_),
    .B1_N(_0937_),
    .X(_1795_));
 sky130_fd_sc_hd__inv_2 _3415_ (.A(_1399_),
    .Y(_1806_));
 sky130_fd_sc_hd__nand2_1 _3416_ (.A(_1795_),
    .B(_1806_),
    .Y(_1817_));
 sky130_fd_sc_hd__nand2_1 _3417_ (.A(_1817_),
    .B(_1366_),
    .Y(_1828_));
 sky130_fd_sc_hd__inv_2 _3418_ (.A(_1344_),
    .Y(_1839_));
 sky130_fd_sc_hd__nand2_1 _3419_ (.A(_1828_),
    .B(_1839_),
    .Y(_1850_));
 sky130_fd_sc_hd__nand2_1 _3420_ (.A(_1850_),
    .B(_1311_),
    .Y(_1861_));
 sky130_fd_sc_hd__o21ai_1 _3421_ (.A1(_1465_),
    .A2(_1861_),
    .B1(_1509_),
    .Y(_1872_));
 sky130_fd_sc_hd__or2_1 _3422_ (.A(_1784_),
    .B(_1872_),
    .X(_1883_));
 sky130_fd_sc_hd__o21ai_1 _3423_ (.A1(_1861_),
    .A2(_1784_),
    .B1(_1872_),
    .Y(_1894_));
 sky130_fd_sc_hd__nand2_2 _3424_ (.A(_1883_),
    .B(_1894_),
    .Y(_1905_));
 sky130_fd_sc_hd__inv_2 _3425_ (.A(_1905_),
    .Y(_1916_));
 sky130_fd_sc_hd__buf_2 _3426_ (.A(_1916_),
    .X(_1927_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(_1465_),
    .Y(_1938_));
 sky130_fd_sc_hd__nand2_1 _3428_ (.A(_1938_),
    .B(_1509_),
    .Y(_1949_));
 sky130_fd_sc_hd__a21oi_1 _3429_ (.A1(_1289_),
    .A2(_1410_),
    .B1(_1575_),
    .Y(_1960_));
 sky130_fd_sc_hd__a21bo_1 _3430_ (.A1(_1960_),
    .A2(_1938_),
    .B1_N(_1487_),
    .X(_1971_));
 sky130_fd_sc_hd__inv_2 _3431_ (.A(_1971_),
    .Y(_1982_));
 sky130_fd_sc_hd__a21o_1 _3432_ (.A1(_1949_),
    .A2(_1960_),
    .B1(_1982_),
    .X(_1993_));
 sky130_fd_sc_hd__nand2_1 _3433_ (.A(_1982_),
    .B(_1949_),
    .Y(_2004_));
 sky130_fd_sc_hd__nand2_2 _3434_ (.A(_1993_),
    .B(_2004_),
    .Y(_2015_));
 sky130_fd_sc_hd__inv_2 _3435_ (.A(_2015_),
    .Y(_2026_));
 sky130_fd_sc_hd__buf_2 _3436_ (.A(_2026_),
    .X(_2037_));
 sky130_fd_sc_hd__inv_2 _3437_ (.A(_1707_),
    .Y(_2048_));
 sky130_fd_sc_hd__mux2_2 _3438_ (.A0(_1927_),
    .A1(_2037_),
    .S(_2048_),
    .X(_2059_));
 sky130_fd_sc_hd__or2_1 _3439_ (.A(_1025_),
    .B(_1146_),
    .X(_2070_));
 sky130_fd_sc_hd__nand2_2 _3440_ (.A(_2070_),
    .B(_1036_),
    .Y(_2080_));
 sky130_fd_sc_hd__clkbuf_4 _3441_ (.A(_2080_),
    .X(_2090_));
 sky130_fd_sc_hd__or2_1 _3442_ (.A(_1168_),
    .B(_1146_),
    .X(_2101_));
 sky130_fd_sc_hd__nand2_1 _3443_ (.A(_2101_),
    .B(_1179_),
    .Y(_2111_));
 sky130_fd_sc_hd__clkbuf_4 _3444_ (.A(_2111_),
    .X(_2120_));
 sky130_fd_sc_hd__mux2_1 _3445_ (.A0(_2090_),
    .A1(_2120_),
    .S(_1707_),
    .X(_2129_));
 sky130_fd_sc_hd__nand2_1 _3446_ (.A(_2059_),
    .B(_2129_),
    .Y(_2138_));
 sky130_fd_sc_hd__or2_1 _3447_ (.A(_1773_),
    .B(_2138_),
    .X(_2148_));
 sky130_fd_sc_hd__or2_1 _3448_ (.A(_1806_),
    .B(_1795_),
    .X(_2158_));
 sky130_fd_sc_hd__and2_1 _3449_ (.A(_2158_),
    .B(_1817_),
    .X(_2168_));
 sky130_fd_sc_hd__clkbuf_4 _3450_ (.A(_2168_),
    .X(_2177_));
 sky130_fd_sc_hd__xor2_2 _3451_ (.A(_1806_),
    .B(_1289_),
    .X(_2187_));
 sky130_fd_sc_hd__mux2_4 _3452_ (.A0(_2177_),
    .A1(_2187_),
    .S(_2048_),
    .X(_2197_));
 sky130_fd_sc_hd__o21ai_1 _3453_ (.A1(_1718_),
    .A2(_2148_),
    .B1(_2197_),
    .Y(_2206_));
 sky130_fd_sc_hd__or2_1 _3454_ (.A(_1839_),
    .B(_1828_),
    .X(_2216_));
 sky130_fd_sc_hd__nand2_1 _3455_ (.A(_2216_),
    .B(_1850_),
    .Y(_2226_));
 sky130_fd_sc_hd__a21bo_1 _3456_ (.A1(_1289_),
    .A2(_1366_),
    .B1_N(_1388_),
    .X(_2235_));
 sky130_fd_sc_hd__xor2_2 _3457_ (.A(_1344_),
    .B(_2235_),
    .X(_2245_));
 sky130_fd_sc_hd__mux2_1 _3458_ (.A0(_2226_),
    .A1(_2245_),
    .S(_2048_),
    .X(_2255_));
 sky130_fd_sc_hd__inv_2 _3459_ (.A(_2255_),
    .Y(_2259_));
 sky130_fd_sc_hd__nor2_1 _3460_ (.A(_2197_),
    .B(_2059_),
    .Y(_2267_));
 sky130_fd_sc_hd__or2_2 _3461_ (.A(_2259_),
    .B(_2267_),
    .X(_2278_));
 sky130_fd_sc_hd__inv_2 _3462_ (.A(_2278_),
    .Y(_2289_));
 sky130_fd_sc_hd__nand2_1 _3463_ (.A(_2206_),
    .B(_2289_),
    .Y(_2300_));
 sky130_fd_sc_hd__inv_2 _3464_ (.A(_1630_),
    .Y(_2311_));
 sky130_fd_sc_hd__clkbuf_4 _3465_ (.A(_2311_),
    .X(_2320_));
 sky130_fd_sc_hd__clkbuf_4 _3466_ (.A(_2320_),
    .X(_2329_));
 sky130_fd_sc_hd__clkbuf_4 _3467_ (.A(_2329_),
    .X(_2339_));
 sky130_fd_sc_hd__inv_2 _3468_ (.A(_2059_),
    .Y(_2349_));
 sky130_fd_sc_hd__or3b_1 _3469_ (.A(_2339_),
    .B(_2349_),
    .C_N(_2129_),
    .X(_2360_));
 sky130_fd_sc_hd__nor2_1 _3470_ (.A(_1773_),
    .B(_2360_),
    .Y(_2370_));
 sky130_fd_sc_hd__inv_2 _3471_ (.A(_1718_),
    .Y(_2380_));
 sky130_fd_sc_hd__inv_2 _3472_ (.A(_2197_),
    .Y(_2390_));
 sky130_fd_sc_hd__a21o_1 _3473_ (.A1(_2370_),
    .A2(_2380_),
    .B1(_2390_),
    .X(_2400_));
 sky130_fd_sc_hd__nand2_1 _3474_ (.A(_2400_),
    .B(_2289_),
    .Y(_2411_));
 sky130_fd_sc_hd__or3_1 _3475_ (.A(_2197_),
    .B(_2259_),
    .C(_2349_),
    .X(_2421_));
 sky130_fd_sc_hd__inv_2 _3476_ (.A(_1773_),
    .Y(_2431_));
 sky130_fd_sc_hd__clkbuf_4 _3477_ (.A(_1630_),
    .X(_2441_));
 sky130_fd_sc_hd__o21ai_1 _3478_ (.A1(_2441_),
    .A2(_2129_),
    .B1(_2059_),
    .Y(_2451_));
 sky130_fd_sc_hd__nand2_1 _3479_ (.A(_2059_),
    .B(_2431_),
    .Y(_2462_));
 sky130_fd_sc_hd__o21ai_1 _3480_ (.A1(_2431_),
    .A2(_2451_),
    .B1(_2462_),
    .Y(_2472_));
 sky130_fd_sc_hd__nand2_1 _3481_ (.A(_2349_),
    .B(_2380_),
    .Y(_2482_));
 sky130_fd_sc_hd__nand2_2 _3482_ (.A(_2255_),
    .B(_2390_),
    .Y(_2493_));
 sky130_fd_sc_hd__inv_2 _3483_ (.A(_2493_),
    .Y(_2503_));
 sky130_fd_sc_hd__nand2_1 _3484_ (.A(_2482_),
    .B(_2503_),
    .Y(_2513_));
 sky130_fd_sc_hd__inv_2 _3485_ (.A(_2513_),
    .Y(_2523_));
 sky130_fd_sc_hd__o21ai_1 _3486_ (.A1(_2380_),
    .A2(_2472_),
    .B1(_2523_),
    .Y(_2534_));
 sky130_fd_sc_hd__a22o_1 _3487_ (.A1(net37),
    .A2(_2421_),
    .B1(_2534_),
    .B2(net36),
    .X(_2544_));
 sky130_fd_sc_hd__a221o_1 _3488_ (.A1(net39),
    .A2(_2300_),
    .B1(net38),
    .B2(_2411_),
    .C1(_2544_),
    .X(_2554_));
 sky130_fd_sc_hd__and2_1 _3489_ (.A(_2462_),
    .B(_2138_),
    .X(_2564_));
 sky130_fd_sc_hd__a21o_1 _3490_ (.A1(_2564_),
    .A2(_1718_),
    .B1(_2513_),
    .X(_2575_));
 sky130_fd_sc_hd__nand2_1 _3491_ (.A(_2360_),
    .B(_2462_),
    .Y(_2585_));
 sky130_fd_sc_hd__o21ai_1 _3492_ (.A1(_2380_),
    .A2(_2585_),
    .B1(_2523_),
    .Y(_2596_));
 sky130_fd_sc_hd__nor2_1 _3493_ (.A(_1773_),
    .B(_2451_),
    .Y(_2606_));
 sky130_fd_sc_hd__o21ai_1 _3494_ (.A1(_2380_),
    .A2(_2606_),
    .B1(_2523_),
    .Y(_2616_));
 sky130_fd_sc_hd__nor2_1 _3495_ (.A(_1718_),
    .B(_2349_),
    .Y(_2627_));
 sky130_fd_sc_hd__inv_2 _3496_ (.A(_2627_),
    .Y(_2637_));
 sky130_fd_sc_hd__and2_1 _3497_ (.A(_2637_),
    .B(_2462_),
    .X(_2648_));
 sky130_fd_sc_hd__o21ai_1 _3498_ (.A1(_2493_),
    .A2(_2648_),
    .B1(net64),
    .Y(_2658_));
 sky130_fd_sc_hd__a21bo_1 _3499_ (.A1(net63),
    .A2(_2616_),
    .B1_N(_2658_),
    .X(_2662_));
 sky130_fd_sc_hd__a221o_1 _3500_ (.A1(net35),
    .A2(_2575_),
    .B1(net34),
    .B2(_2596_),
    .C1(_2662_),
    .X(_2663_));
 sky130_fd_sc_hd__or2_1 _3501_ (.A(_1718_),
    .B(_2421_),
    .X(_2664_));
 sky130_fd_sc_hd__nand2_1 _3502_ (.A(_2472_),
    .B(_2380_),
    .Y(_2665_));
 sky130_fd_sc_hd__or2_1 _3503_ (.A(_2493_),
    .B(_2665_),
    .X(_2666_));
 sky130_fd_sc_hd__and2_1 _3504_ (.A(_2666_),
    .B(net59),
    .X(_2667_));
 sky130_fd_sc_hd__nand2_1 _3505_ (.A(_2148_),
    .B(_2637_),
    .Y(_2668_));
 sky130_fd_sc_hd__nand2_1 _3506_ (.A(_2668_),
    .B(_2503_),
    .Y(_2669_));
 sky130_fd_sc_hd__o21ai_1 _3507_ (.A1(_2380_),
    .A2(_2370_),
    .B1(_2482_),
    .Y(_2670_));
 sky130_fd_sc_hd__or2_1 _3508_ (.A(_2493_),
    .B(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__a22o_1 _3509_ (.A1(net62),
    .A2(_2669_),
    .B1(_2671_),
    .B2(net61),
    .X(_2672_));
 sky130_fd_sc_hd__nor2_1 _3510_ (.A(_1718_),
    .B(_2564_),
    .Y(_2673_));
 sky130_fd_sc_hd__nand2_1 _3511_ (.A(_2673_),
    .B(_2503_),
    .Y(_2674_));
 sky130_fd_sc_hd__nand2_1 _3512_ (.A(_2585_),
    .B(_2380_),
    .Y(_2675_));
 sky130_fd_sc_hd__or2_1 _3513_ (.A(_2493_),
    .B(_2675_),
    .X(_2676_));
 sky130_fd_sc_hd__or2_1 _3514_ (.A(_1718_),
    .B(_2462_),
    .X(_2677_));
 sky130_fd_sc_hd__or2_1 _3515_ (.A(_2493_),
    .B(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__nand2_1 _3516_ (.A(_2606_),
    .B(_2380_),
    .Y(_2679_));
 sky130_fd_sc_hd__or2_1 _3517_ (.A(_2493_),
    .B(_2679_),
    .X(_2680_));
 sky130_fd_sc_hd__a22o_1 _3518_ (.A1(_2678_),
    .A2(net44),
    .B1(_2680_),
    .B2(net33),
    .X(_2681_));
 sky130_fd_sc_hd__a221o_1 _3519_ (.A1(net58),
    .A2(_2674_),
    .B1(_2676_),
    .B2(net55),
    .C1(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__a2111o_1 _3520_ (.A1(net60),
    .A2(_2664_),
    .B1(_2667_),
    .C1(_2672_),
    .D1(_2682_),
    .X(_2683_));
 sky130_fd_sc_hd__a21o_1 _3521_ (.A1(_2670_),
    .A2(_2197_),
    .B1(_2278_),
    .X(_2684_));
 sky130_fd_sc_hd__o21ai_1 _3522_ (.A1(_2390_),
    .A2(_2668_),
    .B1(_2289_),
    .Y(_2685_));
 sky130_fd_sc_hd__inv_2 _3523_ (.A(net46),
    .Y(_2686_));
 sky130_fd_sc_hd__o211a_1 _3524_ (.A1(_2390_),
    .A2(_2380_),
    .B1(_2255_),
    .C1(_2059_),
    .X(_2687_));
 sky130_fd_sc_hd__a21o_1 _3525_ (.A1(_2665_),
    .A2(_2197_),
    .B1(_2278_),
    .X(_2688_));
 sky130_fd_sc_hd__a2bb2o_1 _3526_ (.A1_N(_2686_),
    .A2_N(_2687_),
    .B1(net45),
    .B2(_2688_),
    .X(_2689_));
 sky130_fd_sc_hd__o21ai_1 _3527_ (.A1(_2390_),
    .A2(_2673_),
    .B1(_2289_),
    .Y(_2690_));
 sky130_fd_sc_hd__a21o_1 _3528_ (.A1(_2675_),
    .A2(_2197_),
    .B1(_2278_),
    .X(_2691_));
 sky130_fd_sc_hd__a21o_1 _3529_ (.A1(_2679_),
    .A2(_2197_),
    .B1(_2278_),
    .X(_2692_));
 sky130_fd_sc_hd__a211o_1 _3530_ (.A1(_2677_),
    .A2(_2197_),
    .B1(_2259_),
    .C1(_2267_),
    .X(_2693_));
 sky130_fd_sc_hd__a22o_1 _3531_ (.A1(net40),
    .A2(_2692_),
    .B1(_2693_),
    .B2(net41),
    .X(_2694_));
 sky130_fd_sc_hd__a221o_1 _3532_ (.A1(net43),
    .A2(_2690_),
    .B1(net42),
    .B2(_2691_),
    .C1(_2694_),
    .X(_2695_));
 sky130_fd_sc_hd__a2111o_1 _3533_ (.A1(net47),
    .A2(_2684_),
    .B1(_2685_),
    .C1(_2689_),
    .D1(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__inv_2 _3534_ (.A(_1608_),
    .Y(_2697_));
 sky130_fd_sc_hd__o41a_1 _3535_ (.A1(_2554_),
    .A2(_2663_),
    .A3(_2683_),
    .A4(_2696_),
    .B1(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__and2_1 _3536_ (.A(_2534_),
    .B(net4),
    .X(_2699_));
 sky130_fd_sc_hd__a22o_1 _3537_ (.A1(net7),
    .A2(_2300_),
    .B1(_2411_),
    .B2(net6),
    .X(_2700_));
 sky130_fd_sc_hd__o21a_1 _3538_ (.A1(_2493_),
    .A2(_2648_),
    .B1(net32),
    .X(_2701_));
 sky130_fd_sc_hd__a22o_1 _3539_ (.A1(_2575_),
    .A2(net3),
    .B1(_2596_),
    .B2(net2),
    .X(_2702_));
 sky130_fd_sc_hd__a211o_1 _3540_ (.A1(net31),
    .A2(_2616_),
    .B1(_2701_),
    .C1(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__a2111o_1 _3541_ (.A1(net5),
    .A2(_2421_),
    .B1(_2699_),
    .C1(_2700_),
    .D1(_2703_),
    .X(_2704_));
 sky130_fd_sc_hd__inv_2 _3542_ (.A(net14),
    .Y(_2705_));
 sky130_fd_sc_hd__a2bb2o_1 _3543_ (.A1_N(_2705_),
    .A2_N(_2687_),
    .B1(net13),
    .B2(_2688_),
    .X(_2706_));
 sky130_fd_sc_hd__and2_1 _3544_ (.A(_2691_),
    .B(net10),
    .X(_2707_));
 sky130_fd_sc_hd__a22o_1 _3545_ (.A1(net8),
    .A2(_2692_),
    .B1(_2693_),
    .B2(net9),
    .X(_2708_));
 sky130_fd_sc_hd__a211o_1 _3546_ (.A1(net11),
    .A2(_2690_),
    .B1(_2707_),
    .C1(_2708_),
    .X(_2709_));
 sky130_fd_sc_hd__a2111o_1 _3547_ (.A1(net15),
    .A2(_2684_),
    .B1(_2685_),
    .C1(_2706_),
    .D1(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__and2_1 _3548_ (.A(_2674_),
    .B(net26),
    .X(_2711_));
 sky130_fd_sc_hd__a22o_1 _3549_ (.A1(_2678_),
    .A2(net12),
    .B1(_2680_),
    .B2(net1),
    .X(_2712_));
 sky130_fd_sc_hd__a22o_1 _3550_ (.A1(net30),
    .A2(_2669_),
    .B1(_2671_),
    .B2(net29),
    .X(_2713_));
 sky130_fd_sc_hd__a221o_1 _3551_ (.A1(net28),
    .A2(_2664_),
    .B1(net27),
    .B2(_2666_),
    .C1(_2713_),
    .X(_2714_));
 sky130_fd_sc_hd__a2111o_1 _3552_ (.A1(net23),
    .A2(_2676_),
    .B1(_2711_),
    .C1(_2712_),
    .D1(_2714_),
    .X(_2715_));
 sky130_fd_sc_hd__o31a_1 _3553_ (.A1(_2704_),
    .A2(_2710_),
    .A3(_2715_),
    .B1(_1685_),
    .X(_2716_));
 sky130_fd_sc_hd__or2_4 _3554_ (.A(_2698_),
    .B(_2716_),
    .X(_2717_));
 sky130_fd_sc_hd__inv_2 _3555_ (.A(_0761_),
    .Y(_2718_));
 sky130_fd_sc_hd__buf_6 _3556_ (.A(_2718_),
    .X(_2719_));
 sky130_fd_sc_hd__a21oi_1 _3557_ (.A1(_2719_),
    .A2(net129),
    .B1(_2717_),
    .Y(_2720_));
 sky130_fd_sc_hd__inv_2 _3558_ (.A(net130),
    .Y(_2721_));
 sky130_fd_sc_hd__nor2_1 _3559_ (.A(net138),
    .B(net131),
    .Y(_2722_));
 sky130_fd_sc_hd__mux2_1 _3560_ (.A0(net135),
    .A1(net139),
    .S(_0706_),
    .X(_2723_));
 sky130_fd_sc_hd__mux2_1 _3561_ (.A0(net140),
    .A1(net136),
    .S(_0783_),
    .X(_2724_));
 sky130_fd_sc_hd__clkbuf_4 _3562_ (.A(_0849_),
    .X(_2725_));
 sky130_fd_sc_hd__clkbuf_4 _3563_ (.A(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__mux2_1 _3564_ (.A0(net141),
    .A1(net137),
    .S(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__mux2_1 _3565_ (.A0(net171),
    .A1(net144),
    .S(_0684_),
    .X(_2728_));
 sky130_fd_sc_hd__o21a_1 _3566_ (.A1(_0684_),
    .A2(net144),
    .B1(\M000[25] ),
    .X(_2729_));
 sky130_fd_sc_hd__a21oi_1 _3567_ (.A1(_2728_),
    .A2(_0761_),
    .B1(net145),
    .Y(_2730_));
 sky130_fd_sc_hd__nand2_1 _3568_ (.A(net146),
    .B(_0849_),
    .Y(_2731_));
 sky130_fd_sc_hd__buf_2 _3569_ (.A(net147),
    .X(_2732_));
 sky130_fd_sc_hd__clkbuf_4 _3570_ (.A(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__nand2_1 _3571_ (.A(net142),
    .B(_2733_),
    .Y(_2734_));
 sky130_fd_sc_hd__nand2_1 _3572_ (.A(_2722_),
    .B(net143),
    .Y(_2735_));
 sky130_fd_sc_hd__nand2_2 _3573_ (.A(_2735_),
    .B(_0893_),
    .Y(_2736_));
 sky130_fd_sc_hd__inv_2 _3574_ (.A(net67),
    .Y(_2737_));
 sky130_fd_sc_hd__inv_2 _3575_ (.A(net66),
    .Y(_2738_));
 sky130_fd_sc_hd__and3_2 _3576_ (.A(_2737_),
    .B(_2738_),
    .C(net65),
    .X(_2739_));
 sky130_fd_sc_hd__buf_2 _3577_ (.A(_2739_),
    .X(_2740_));
 sky130_fd_sc_hd__or2b_1 _3578_ (.A(_2736_),
    .B_N(_2740_),
    .X(_2741_));
 sky130_fd_sc_hd__buf_2 _3579_ (.A(_2026_),
    .X(_2742_));
 sky130_fd_sc_hd__nand2_1 _3580_ (.A(_2742_),
    .B(net31),
    .Y(_2743_));
 sky130_fd_sc_hd__nand2_1 _3581_ (.A(_2026_),
    .B(net32),
    .Y(_2744_));
 sky130_fd_sc_hd__mux2_1 _3582_ (.A0(_2743_),
    .A1(_2744_),
    .S(_2320_),
    .X(_2745_));
 sky130_fd_sc_hd__nand2_1 _3583_ (.A(_2742_),
    .B(net2),
    .Y(_2746_));
 sky130_fd_sc_hd__nand2_1 _3584_ (.A(_2026_),
    .B(net3),
    .Y(_2747_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(_2746_),
    .A1(_2747_),
    .S(_2320_),
    .X(_2748_));
 sky130_fd_sc_hd__inv_2 _3586_ (.A(_2080_),
    .Y(_2749_));
 sky130_fd_sc_hd__mux2_1 _3587_ (.A0(_2745_),
    .A1(_2748_),
    .S(_2749_),
    .X(_2750_));
 sky130_fd_sc_hd__nand2_1 _3588_ (.A(_2742_),
    .B(net27),
    .Y(_2751_));
 sky130_fd_sc_hd__nand2_1 _3589_ (.A(_2742_),
    .B(net28),
    .Y(_2752_));
 sky130_fd_sc_hd__clkbuf_4 _3590_ (.A(_2311_),
    .X(_2753_));
 sky130_fd_sc_hd__mux2_1 _3591_ (.A0(_2751_),
    .A1(_2752_),
    .S(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__nand2_1 _3592_ (.A(_2742_),
    .B(net29),
    .Y(_2755_));
 sky130_fd_sc_hd__nand2_1 _3593_ (.A(_2742_),
    .B(net30),
    .Y(_2756_));
 sky130_fd_sc_hd__mux2_1 _3594_ (.A0(_2755_),
    .A1(_2756_),
    .S(_2753_),
    .X(_2757_));
 sky130_fd_sc_hd__clkbuf_4 _3595_ (.A(_2749_),
    .X(_2758_));
 sky130_fd_sc_hd__mux2_1 _3596_ (.A0(_2754_),
    .A1(_2757_),
    .S(_2758_),
    .X(_2759_));
 sky130_fd_sc_hd__inv_2 _3597_ (.A(_1729_),
    .Y(_2760_));
 sky130_fd_sc_hd__mux2_1 _3598_ (.A0(_2750_),
    .A1(_2759_),
    .S(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__nand2_1 _3599_ (.A(_2742_),
    .B(net8),
    .Y(_2762_));
 sky130_fd_sc_hd__nand2_1 _3600_ (.A(_2026_),
    .B(net9),
    .Y(_2763_));
 sky130_fd_sc_hd__mux2_1 _3601_ (.A0(_2762_),
    .A1(_2763_),
    .S(_2753_),
    .X(_2764_));
 sky130_fd_sc_hd__nand2_1 _3602_ (.A(_2026_),
    .B(net10),
    .Y(_2765_));
 sky130_fd_sc_hd__nand2_1 _3603_ (.A(_2037_),
    .B(net11),
    .Y(_2766_));
 sky130_fd_sc_hd__mux2_1 _3604_ (.A0(_2765_),
    .A1(_2766_),
    .S(_2753_),
    .X(_2767_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(_2764_),
    .A1(_2767_),
    .S(_2758_),
    .X(_2768_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(_2742_),
    .B(net4),
    .Y(_2769_));
 sky130_fd_sc_hd__nand2_1 _3607_ (.A(_2026_),
    .B(net5),
    .Y(_2770_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(_2769_),
    .A1(_2770_),
    .S(_2320_),
    .X(_2771_));
 sky130_fd_sc_hd__nand2_1 _3609_ (.A(_2026_),
    .B(net6),
    .Y(_2772_));
 sky130_fd_sc_hd__nand2_1 _3610_ (.A(_2742_),
    .B(net7),
    .Y(_2773_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(_2772_),
    .A1(_2773_),
    .S(_2320_),
    .X(_2774_));
 sky130_fd_sc_hd__mux2_1 _3612_ (.A0(_2771_),
    .A1(_2774_),
    .S(_2749_),
    .X(_2775_));
 sky130_fd_sc_hd__mux2_1 _3613_ (.A0(_2768_),
    .A1(_2775_),
    .S(_2760_),
    .X(_2776_));
 sky130_fd_sc_hd__mux2_1 _3614_ (.A0(_2761_),
    .A1(_2776_),
    .S(_1124_),
    .X(_2777_));
 sky130_fd_sc_hd__clkbuf_4 _3615_ (.A(_2187_),
    .X(_2778_));
 sky130_fd_sc_hd__inv_2 _3616_ (.A(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__clkbuf_4 _3617_ (.A(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__nand2_1 _3618_ (.A(_2777_),
    .B(_2780_),
    .Y(_2781_));
 sky130_fd_sc_hd__clkbuf_4 _3619_ (.A(_2758_),
    .X(_2782_));
 sky130_fd_sc_hd__nand2_1 _3620_ (.A(_2037_),
    .B(net13),
    .Y(_2783_));
 sky130_fd_sc_hd__nand2_1 _3621_ (.A(_2037_),
    .B(net14),
    .Y(_2784_));
 sky130_fd_sc_hd__mux2_1 _3622_ (.A0(_2783_),
    .A1(_2784_),
    .S(_2339_),
    .X(_2785_));
 sky130_fd_sc_hd__o21ai_1 _3623_ (.A1(net15),
    .A2(_2339_),
    .B1(_2037_),
    .Y(_2786_));
 sky130_fd_sc_hd__or2_1 _3624_ (.A(_2090_),
    .B(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__o21ai_1 _3625_ (.A1(_2782_),
    .A2(_2785_),
    .B1(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__clkbuf_4 _3626_ (.A(_2760_),
    .X(_2789_));
 sky130_fd_sc_hd__nand2_1 _3627_ (.A(_2788_),
    .B(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__or2_1 _3628_ (.A(_1135_),
    .B(_2790_),
    .X(_2791_));
 sky130_fd_sc_hd__inv_2 _3629_ (.A(_2245_),
    .Y(_2792_));
 sky130_fd_sc_hd__nor2_2 _3630_ (.A(_1674_),
    .B(_2792_),
    .Y(_2793_));
 sky130_fd_sc_hd__inv_2 _3631_ (.A(_2793_),
    .Y(_2794_));
 sky130_fd_sc_hd__a21oi_1 _3632_ (.A1(_2791_),
    .A2(_2778_),
    .B1(_2794_),
    .Y(_2795_));
 sky130_fd_sc_hd__a22o_1 _3633_ (.A1(net27),
    .A2(_1674_),
    .B1(_2781_),
    .B2(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__inv_2 _3634_ (.A(_2796_),
    .Y(_2797_));
 sky130_fd_sc_hd__buf_2 _3635_ (.A(_1916_),
    .X(_2798_));
 sky130_fd_sc_hd__nand2_1 _3636_ (.A(_2798_),
    .B(net63),
    .Y(_2799_));
 sky130_fd_sc_hd__nand2_1 _3637_ (.A(_2798_),
    .B(net64),
    .Y(_2800_));
 sky130_fd_sc_hd__mux2_1 _3638_ (.A0(_2799_),
    .A1(_2800_),
    .S(_2329_),
    .X(_2801_));
 sky130_fd_sc_hd__nand2_1 _3639_ (.A(_2798_),
    .B(net34),
    .Y(_2802_));
 sky130_fd_sc_hd__nand2_1 _3640_ (.A(_2798_),
    .B(net35),
    .Y(_2803_));
 sky130_fd_sc_hd__mux2_1 _3641_ (.A0(_2802_),
    .A1(_2803_),
    .S(_2329_),
    .X(_2804_));
 sky130_fd_sc_hd__inv_2 _3642_ (.A(_2111_),
    .Y(_2805_));
 sky130_fd_sc_hd__mux2_1 _3643_ (.A0(_2801_),
    .A1(_2804_),
    .S(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__nand2_1 _3644_ (.A(_1927_),
    .B(net59),
    .Y(_2807_));
 sky130_fd_sc_hd__nand2_1 _3645_ (.A(_2798_),
    .B(net60),
    .Y(_2808_));
 sky130_fd_sc_hd__buf_4 _3646_ (.A(_2753_),
    .X(_2809_));
 sky130_fd_sc_hd__mux2_1 _3647_ (.A0(_2807_),
    .A1(_2808_),
    .S(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__nand2_1 _3648_ (.A(_2798_),
    .B(net61),
    .Y(_2811_));
 sky130_fd_sc_hd__nand2_1 _3649_ (.A(_1927_),
    .B(net62),
    .Y(_2812_));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(_2811_),
    .A1(_2812_),
    .S(_2809_),
    .X(_2813_));
 sky130_fd_sc_hd__clkbuf_4 _3651_ (.A(_2805_),
    .X(_2814_));
 sky130_fd_sc_hd__mux2_1 _3652_ (.A0(_2810_),
    .A1(_2813_),
    .S(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__inv_2 _3653_ (.A(_1762_),
    .Y(_2816_));
 sky130_fd_sc_hd__mux2_1 _3654_ (.A0(_2806_),
    .A1(_2815_),
    .S(_2816_),
    .X(_2817_));
 sky130_fd_sc_hd__nand2_1 _3655_ (.A(_2798_),
    .B(net40),
    .Y(_2818_));
 sky130_fd_sc_hd__nand2_1 _3656_ (.A(_1916_),
    .B(net41),
    .Y(_2819_));
 sky130_fd_sc_hd__mux2_1 _3657_ (.A0(_2818_),
    .A1(_2819_),
    .S(_2809_),
    .X(_2820_));
 sky130_fd_sc_hd__nand2_1 _3658_ (.A(_2798_),
    .B(net42),
    .Y(_2821_));
 sky130_fd_sc_hd__nand2_1 _3659_ (.A(_1916_),
    .B(net43),
    .Y(_2822_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(_2821_),
    .A1(_2822_),
    .S(_2809_),
    .X(_2823_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(_2820_),
    .A1(_2823_),
    .S(_2814_),
    .X(_2824_));
 sky130_fd_sc_hd__nand2_1 _3662_ (.A(_2798_),
    .B(net36),
    .Y(_2825_));
 sky130_fd_sc_hd__nand2_1 _3663_ (.A(_1916_),
    .B(net37),
    .Y(_2826_));
 sky130_fd_sc_hd__mux2_1 _3664_ (.A0(_2825_),
    .A1(_2826_),
    .S(_2809_),
    .X(_2827_));
 sky130_fd_sc_hd__nand2_1 _3665_ (.A(_1916_),
    .B(net38),
    .Y(_2828_));
 sky130_fd_sc_hd__nand2_1 _3666_ (.A(_1916_),
    .B(net39),
    .Y(_2829_));
 sky130_fd_sc_hd__mux2_1 _3667_ (.A0(_2828_),
    .A1(_2829_),
    .S(_2329_),
    .X(_2830_));
 sky130_fd_sc_hd__mux2_1 _3668_ (.A0(_2827_),
    .A1(_2830_),
    .S(_2805_),
    .X(_2831_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(_2824_),
    .A1(_2831_),
    .S(_2816_),
    .X(_2832_));
 sky130_fd_sc_hd__mux2_1 _3670_ (.A0(_2817_),
    .A1(_2832_),
    .S(_1245_),
    .X(_2833_));
 sky130_fd_sc_hd__inv_2 _3671_ (.A(_2177_),
    .Y(_2834_));
 sky130_fd_sc_hd__nand2_1 _3672_ (.A(_2833_),
    .B(_2834_),
    .Y(_2835_));
 sky130_fd_sc_hd__inv_2 _3673_ (.A(_2226_),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_1 _3674_ (.A(_1608_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__clkbuf_4 _3675_ (.A(_2837_),
    .X(_2838_));
 sky130_fd_sc_hd__clkbuf_4 _3676_ (.A(_1245_),
    .X(_2839_));
 sky130_fd_sc_hd__buf_2 _3677_ (.A(_2814_),
    .X(_2840_));
 sky130_fd_sc_hd__nand2_1 _3678_ (.A(_2798_),
    .B(net45),
    .Y(_2841_));
 sky130_fd_sc_hd__nand2_1 _3679_ (.A(_1927_),
    .B(net46),
    .Y(_2842_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(_2841_),
    .A1(_2842_),
    .S(_2339_),
    .X(_2843_));
 sky130_fd_sc_hd__o21ai_1 _3681_ (.A1(net47),
    .A2(_2339_),
    .B1(_1927_),
    .Y(_2844_));
 sky130_fd_sc_hd__or2_1 _3682_ (.A(_2120_),
    .B(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__o21ai_1 _3683_ (.A1(_2840_),
    .A2(_2843_),
    .B1(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__clkbuf_4 _3684_ (.A(_2816_),
    .X(_2847_));
 sky130_fd_sc_hd__nand2_1 _3685_ (.A(_2846_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__or2_1 _3686_ (.A(_2839_),
    .B(_2848_),
    .X(_2849_));
 sky130_fd_sc_hd__nand2_1 _3687_ (.A(_2849_),
    .B(_2177_),
    .Y(_2850_));
 sky130_fd_sc_hd__buf_2 _3688_ (.A(_1608_),
    .X(_2851_));
 sky130_fd_sc_hd__a32o_1 _3689_ (.A1(_2835_),
    .A2(_2838_),
    .A3(_2850_),
    .B1(net59),
    .B2(_2851_),
    .X(_2852_));
 sky130_fd_sc_hd__or2_1 _3690_ (.A(_2797_),
    .B(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__nand2_1 _3691_ (.A(_2852_),
    .B(_2797_),
    .Y(_2854_));
 sky130_fd_sc_hd__nand2_1 _3692_ (.A(_2853_),
    .B(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(_2766_),
    .A1(_2783_),
    .S(_2329_),
    .X(_2856_));
 sky130_fd_sc_hd__or2_1 _3694_ (.A(_2311_),
    .B(_2763_),
    .X(_2857_));
 sky130_fd_sc_hd__o21a_1 _3695_ (.A1(_1630_),
    .A2(_2765_),
    .B1(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__or2_1 _3696_ (.A(_2749_),
    .B(_2858_),
    .X(_2859_));
 sky130_fd_sc_hd__o21a_1 _3697_ (.A1(_2080_),
    .A2(_2856_),
    .B1(_2859_),
    .X(_2860_));
 sky130_fd_sc_hd__or2_1 _3698_ (.A(_2320_),
    .B(_2770_),
    .X(_2861_));
 sky130_fd_sc_hd__o21a_1 _3699_ (.A1(_1630_),
    .A2(_2772_),
    .B1(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__mux2_1 _3700_ (.A0(_2773_),
    .A1(_2762_),
    .S(_2320_),
    .X(_2863_));
 sky130_fd_sc_hd__mux2_1 _3701_ (.A0(_2862_),
    .A1(_2863_),
    .S(_2758_),
    .X(_2864_));
 sky130_fd_sc_hd__mux2_1 _3702_ (.A0(_2860_),
    .A1(_2864_),
    .S(_2760_),
    .X(_2865_));
 sky130_fd_sc_hd__mux2_1 _3703_ (.A0(_2752_),
    .A1(_2755_),
    .S(_2753_),
    .X(_2866_));
 sky130_fd_sc_hd__mux2_1 _3704_ (.A0(_2756_),
    .A1(_2743_),
    .S(_2753_),
    .X(_2867_));
 sky130_fd_sc_hd__mux2_1 _3705_ (.A0(_2866_),
    .A1(_2867_),
    .S(_2758_),
    .X(_2868_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(_2744_),
    .A1(_2746_),
    .S(_2753_),
    .X(_2869_));
 sky130_fd_sc_hd__mux2_1 _3707_ (.A0(_2747_),
    .A1(_2769_),
    .S(_2753_),
    .X(_2870_));
 sky130_fd_sc_hd__mux2_1 _3708_ (.A0(_2869_),
    .A1(_2870_),
    .S(_2758_),
    .X(_2871_));
 sky130_fd_sc_hd__mux2_1 _3709_ (.A0(_2868_),
    .A1(_2871_),
    .S(_1729_),
    .X(_2872_));
 sky130_fd_sc_hd__inv_2 _3710_ (.A(_1124_),
    .Y(_2873_));
 sky130_fd_sc_hd__mux2_1 _3711_ (.A0(_2865_),
    .A1(_2872_),
    .S(_2873_),
    .X(_2874_));
 sky130_fd_sc_hd__nand2_1 _3712_ (.A(_2874_),
    .B(_2780_),
    .Y(_2875_));
 sky130_fd_sc_hd__nand2_1 _3713_ (.A(_2329_),
    .B(net15),
    .Y(_2876_));
 sky130_fd_sc_hd__o22a_1 _3714_ (.A1(_2015_),
    .A2(_2876_),
    .B1(_2809_),
    .B2(_2784_),
    .X(_2877_));
 sky130_fd_sc_hd__nor2_1 _3715_ (.A(_2758_),
    .B(_2877_),
    .Y(_2878_));
 sky130_fd_sc_hd__a31o_1 _3716_ (.A1(_2441_),
    .A2(_2758_),
    .A3(_2037_),
    .B1(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__nand2_1 _3717_ (.A(_2879_),
    .B(_2789_),
    .Y(_2880_));
 sky130_fd_sc_hd__or2_1 _3718_ (.A(_1124_),
    .B(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__a21oi_1 _3719_ (.A1(_2881_),
    .A2(_2778_),
    .B1(_2794_),
    .Y(_2882_));
 sky130_fd_sc_hd__a22o_1 _3720_ (.A1(net28),
    .A2(_1674_),
    .B1(_2875_),
    .B2(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__inv_2 _3721_ (.A(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__or2_1 _3722_ (.A(_2753_),
    .B(_2819_),
    .X(_2885_));
 sky130_fd_sc_hd__o21ai_1 _3723_ (.A1(_1630_),
    .A2(_2821_),
    .B1(_2885_),
    .Y(_2886_));
 sky130_fd_sc_hd__or2_1 _3724_ (.A(_2320_),
    .B(_2822_),
    .X(_2887_));
 sky130_fd_sc_hd__o21ai_1 _3725_ (.A1(_1630_),
    .A2(_2841_),
    .B1(_2887_),
    .Y(_2888_));
 sky130_fd_sc_hd__mux2_1 _3726_ (.A0(_2886_),
    .A1(_2888_),
    .S(_2805_),
    .X(_2889_));
 sky130_fd_sc_hd__or2_1 _3727_ (.A(_2320_),
    .B(_2829_),
    .X(_2890_));
 sky130_fd_sc_hd__o21ai_1 _3728_ (.A1(_1630_),
    .A2(_2818_),
    .B1(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__mux2_1 _3729_ (.A0(_2826_),
    .A1(_2828_),
    .S(_2320_),
    .X(_2892_));
 sky130_fd_sc_hd__nand2_1 _3730_ (.A(_2892_),
    .B(_2111_),
    .Y(_2893_));
 sky130_fd_sc_hd__o21ai_1 _3731_ (.A1(_2120_),
    .A2(_2891_),
    .B1(_2893_),
    .Y(_2894_));
 sky130_fd_sc_hd__inv_2 _3732_ (.A(_2894_),
    .Y(_2895_));
 sky130_fd_sc_hd__mux2_1 _3733_ (.A0(_2889_),
    .A1(_2895_),
    .S(_2816_),
    .X(_2896_));
 sky130_fd_sc_hd__inv_2 _3734_ (.A(_2896_),
    .Y(_2897_));
 sky130_fd_sc_hd__mux2_1 _3735_ (.A0(_2808_),
    .A1(_2811_),
    .S(_2329_),
    .X(_2898_));
 sky130_fd_sc_hd__mux2_1 _3736_ (.A0(_2812_),
    .A1(_2799_),
    .S(_2809_),
    .X(_2899_));
 sky130_fd_sc_hd__mux2_1 _3737_ (.A0(_2898_),
    .A1(_2899_),
    .S(_2814_),
    .X(_2900_));
 sky130_fd_sc_hd__mux2_1 _3738_ (.A0(_2800_),
    .A1(_2802_),
    .S(_2809_),
    .X(_2901_));
 sky130_fd_sc_hd__o2111ai_1 _3739_ (.A1(_1784_),
    .A2(_1872_),
    .B1(net35),
    .C1(_2441_),
    .D1(_1894_),
    .Y(_2902_));
 sky130_fd_sc_hd__o21a_1 _3740_ (.A1(_2441_),
    .A2(_2825_),
    .B1(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(_2901_),
    .A1(_2903_),
    .S(_2805_),
    .X(_2904_));
 sky130_fd_sc_hd__mux2_1 _3742_ (.A0(_2900_),
    .A1(_2904_),
    .S(_1762_),
    .X(_2905_));
 sky130_fd_sc_hd__inv_2 _3743_ (.A(_1245_),
    .Y(_2906_));
 sky130_fd_sc_hd__mux2_1 _3744_ (.A0(_2897_),
    .A1(_2905_),
    .S(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__nand2_1 _3745_ (.A(_2907_),
    .B(_2834_),
    .Y(_2908_));
 sky130_fd_sc_hd__nand2_1 _3746_ (.A(_2339_),
    .B(net47),
    .Y(_2909_));
 sky130_fd_sc_hd__o22a_1 _3747_ (.A1(_1905_),
    .A2(_2909_),
    .B1(_2339_),
    .B2(_2842_),
    .X(_2910_));
 sky130_fd_sc_hd__nor2_1 _3748_ (.A(_2814_),
    .B(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__a31o_1 _3749_ (.A1(_2840_),
    .A2(_2441_),
    .A3(_1927_),
    .B1(_2911_),
    .X(_2912_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(_2912_),
    .B(_2816_),
    .Y(_2913_));
 sky130_fd_sc_hd__or2_1 _3751_ (.A(_2839_),
    .B(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__nand2_1 _3752_ (.A(_2914_),
    .B(_2177_),
    .Y(_2915_));
 sky130_fd_sc_hd__a32o_1 _3753_ (.A1(_2908_),
    .A2(_2838_),
    .A3(_2915_),
    .B1(net60),
    .B2(_1608_),
    .X(_2916_));
 sky130_fd_sc_hd__or2_1 _3754_ (.A(_2884_),
    .B(_2916_),
    .X(_2917_));
 sky130_fd_sc_hd__nand2_1 _3755_ (.A(_2916_),
    .B(_2884_),
    .Y(_2918_));
 sky130_fd_sc_hd__nand2_2 _3756_ (.A(_2917_),
    .B(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__or2_1 _3757_ (.A(_2855_),
    .B(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__clkbuf_4 _3758_ (.A(_1762_),
    .X(_2921_));
 sky130_fd_sc_hd__nand2_1 _3759_ (.A(_1927_),
    .B(net58),
    .Y(_2922_));
 sky130_fd_sc_hd__mux2_1 _3760_ (.A0(_2922_),
    .A1(_2807_),
    .S(_2339_),
    .X(_2923_));
 sky130_fd_sc_hd__or2_1 _3761_ (.A(_2840_),
    .B(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__o21ai_1 _3762_ (.A1(_2120_),
    .A2(_2898_),
    .B1(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__mux2_1 _3763_ (.A0(_2899_),
    .A1(_2901_),
    .S(_2840_),
    .X(_2926_));
 sky130_fd_sc_hd__nand2_1 _3764_ (.A(_2926_),
    .B(_2921_),
    .Y(_2927_));
 sky130_fd_sc_hd__o21ai_1 _3765_ (.A1(_2921_),
    .A2(_2925_),
    .B1(_2927_),
    .Y(_2928_));
 sky130_fd_sc_hd__mux2_1 _3766_ (.A0(_2891_),
    .A1(_2886_),
    .S(_2840_),
    .X(_2929_));
 sky130_fd_sc_hd__mux2_1 _3767_ (.A0(_2892_),
    .A1(_2903_),
    .S(_2120_),
    .X(_2930_));
 sky130_fd_sc_hd__nand2_1 _3768_ (.A(_2930_),
    .B(_2847_),
    .Y(_2931_));
 sky130_fd_sc_hd__o21ai_1 _3769_ (.A1(_2847_),
    .A2(_2929_),
    .B1(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__mux2_1 _3770_ (.A0(_2928_),
    .A1(_2932_),
    .S(_2839_),
    .X(_2933_));
 sky130_fd_sc_hd__clkbuf_4 _3771_ (.A(_2834_),
    .X(_2934_));
 sky130_fd_sc_hd__nand2_1 _3772_ (.A(_2933_),
    .B(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__nand2_1 _3773_ (.A(_2910_),
    .B(_2814_),
    .Y(_2936_));
 sky130_fd_sc_hd__o21ai_1 _3774_ (.A1(_2840_),
    .A2(_2888_),
    .B1(_2936_),
    .Y(_2937_));
 sky130_fd_sc_hd__inv_2 _3775_ (.A(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__and3_1 _3776_ (.A(_1927_),
    .B(_2120_),
    .C(_2441_),
    .X(_2939_));
 sky130_fd_sc_hd__mux2_1 _3777_ (.A0(_2938_),
    .A1(_2939_),
    .S(_1762_),
    .X(_2940_));
 sky130_fd_sc_hd__buf_2 _3778_ (.A(_2906_),
    .X(_2941_));
 sky130_fd_sc_hd__a21o_1 _3779_ (.A1(_2940_),
    .A2(_2941_),
    .B1(_2934_),
    .X(_2942_));
 sky130_fd_sc_hd__a32o_1 _3780_ (.A1(_2935_),
    .A2(_2838_),
    .A3(_2942_),
    .B1(net58),
    .B2(_2851_),
    .X(_2943_));
 sky130_fd_sc_hd__mux2_1 _3781_ (.A0(_2858_),
    .A1(_2863_),
    .S(_2090_),
    .X(_2944_));
 sky130_fd_sc_hd__mux2_1 _3782_ (.A0(_2862_),
    .A1(_2870_),
    .S(_2090_),
    .X(_2945_));
 sky130_fd_sc_hd__mux2_1 _3783_ (.A0(_2944_),
    .A1(_2945_),
    .S(_2789_),
    .X(_2946_));
 sky130_fd_sc_hd__nand2_1 _3784_ (.A(_2037_),
    .B(net26),
    .Y(_2947_));
 sky130_fd_sc_hd__mux2_1 _3785_ (.A0(_2947_),
    .A1(_2751_),
    .S(_2809_),
    .X(_2948_));
 sky130_fd_sc_hd__mux2_1 _3786_ (.A0(_2948_),
    .A1(_2866_),
    .S(_2782_),
    .X(_2949_));
 sky130_fd_sc_hd__mux2_1 _3787_ (.A0(_2867_),
    .A1(_2869_),
    .S(_2782_),
    .X(_2950_));
 sky130_fd_sc_hd__buf_2 _3788_ (.A(_1729_),
    .X(_2951_));
 sky130_fd_sc_hd__mux2_1 _3789_ (.A0(_2949_),
    .A1(_2950_),
    .S(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__buf_2 _3790_ (.A(_2873_),
    .X(_2953_));
 sky130_fd_sc_hd__mux2_1 _3791_ (.A0(_2946_),
    .A1(_2952_),
    .S(_2953_),
    .X(_2954_));
 sky130_fd_sc_hd__nand2_1 _3792_ (.A(_2954_),
    .B(_2780_),
    .Y(_2955_));
 sky130_fd_sc_hd__or2_1 _3793_ (.A(_2090_),
    .B(_2877_),
    .X(_2956_));
 sky130_fd_sc_hd__o21a_1 _3794_ (.A1(_2782_),
    .A2(_2856_),
    .B1(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__and3_1 _3795_ (.A(_2037_),
    .B(_2441_),
    .C(_2090_),
    .X(_2958_));
 sky130_fd_sc_hd__nand2_1 _3796_ (.A(_2958_),
    .B(_2951_),
    .Y(_2959_));
 sky130_fd_sc_hd__o21ai_1 _3797_ (.A1(_2951_),
    .A2(_2957_),
    .B1(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__buf_2 _3798_ (.A(_2953_),
    .X(_2961_));
 sky130_fd_sc_hd__nand2_1 _3799_ (.A(_2960_),
    .B(_2961_),
    .Y(_2962_));
 sky130_fd_sc_hd__nand2_1 _3800_ (.A(_2962_),
    .B(_2778_),
    .Y(_2963_));
 sky130_fd_sc_hd__buf_2 _3801_ (.A(_1674_),
    .X(_2964_));
 sky130_fd_sc_hd__buf_2 _3802_ (.A(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__a32o_1 _3803_ (.A1(_2955_),
    .A2(_2793_),
    .A3(_2963_),
    .B1(net26),
    .B2(_2965_),
    .X(_2966_));
 sky130_fd_sc_hd__or2b_1 _3804_ (.A(_2943_),
    .B_N(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__or2b_1 _3805_ (.A(_2966_),
    .B_N(_2943_),
    .X(_2968_));
 sky130_fd_sc_hd__nand2_2 _3806_ (.A(_2967_),
    .B(_2968_),
    .Y(_2969_));
 sky130_fd_sc_hd__mux2_1 _3807_ (.A0(_2757_),
    .A1(_2745_),
    .S(_2782_),
    .X(_2970_));
 sky130_fd_sc_hd__nand2_1 _3808_ (.A(_2037_),
    .B(net23),
    .Y(_2971_));
 sky130_fd_sc_hd__mux2_1 _3809_ (.A0(_2971_),
    .A1(_2947_),
    .S(_2329_),
    .X(_2972_));
 sky130_fd_sc_hd__mux2_1 _3810_ (.A0(_2972_),
    .A1(_2754_),
    .S(_2782_),
    .X(_2973_));
 sky130_fd_sc_hd__mux2_1 _3811_ (.A0(_2970_),
    .A1(_2973_),
    .S(_2789_),
    .X(_2974_));
 sky130_fd_sc_hd__mux2_1 _3812_ (.A0(_2748_),
    .A1(_2771_),
    .S(_2782_),
    .X(_2975_));
 sky130_fd_sc_hd__mux2_1 _3813_ (.A0(_2774_),
    .A1(_2764_),
    .S(_2782_),
    .X(_2976_));
 sky130_fd_sc_hd__mux2_1 _3814_ (.A0(_2975_),
    .A1(_2976_),
    .S(_1729_),
    .X(_2977_));
 sky130_fd_sc_hd__mux2_1 _3815_ (.A0(_2974_),
    .A1(_2977_),
    .S(_1135_),
    .X(_2978_));
 sky130_fd_sc_hd__nand2_1 _3816_ (.A(_2978_),
    .B(_2780_),
    .Y(_2979_));
 sky130_fd_sc_hd__or2_1 _3817_ (.A(_2758_),
    .B(_2767_),
    .X(_2980_));
 sky130_fd_sc_hd__o21a_1 _3818_ (.A1(_2090_),
    .A2(_2785_),
    .B1(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__nor2_1 _3819_ (.A(_2782_),
    .B(_2786_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _3820_ (.A(_2982_),
    .B(_2951_),
    .Y(_2983_));
 sky130_fd_sc_hd__o21ai_1 _3821_ (.A1(_2951_),
    .A2(_2981_),
    .B1(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__nand2_1 _3822_ (.A(_2984_),
    .B(_2953_),
    .Y(_2985_));
 sky130_fd_sc_hd__a21oi_1 _3823_ (.A1(_2985_),
    .A2(_2778_),
    .B1(_2794_),
    .Y(_2986_));
 sky130_fd_sc_hd__a22o_1 _3824_ (.A1(net23),
    .A2(_2964_),
    .B1(_2979_),
    .B2(_2986_),
    .X(_2987_));
 sky130_fd_sc_hd__inv_2 _3825_ (.A(_2987_),
    .Y(_2988_));
 sky130_fd_sc_hd__mux2_1 _3826_ (.A0(_2813_),
    .A1(_2801_),
    .S(_2840_),
    .X(_2989_));
 sky130_fd_sc_hd__nand2_1 _3827_ (.A(_1927_),
    .B(net55),
    .Y(_2990_));
 sky130_fd_sc_hd__mux2_1 _3828_ (.A0(_2990_),
    .A1(_2922_),
    .S(_2339_),
    .X(_2991_));
 sky130_fd_sc_hd__mux2_1 _3829_ (.A0(_2991_),
    .A1(_2810_),
    .S(_2840_),
    .X(_2992_));
 sky130_fd_sc_hd__mux2_1 _3830_ (.A0(_2989_),
    .A1(_2992_),
    .S(_2847_),
    .X(_2993_));
 sky130_fd_sc_hd__mux2_1 _3831_ (.A0(_2804_),
    .A1(_2827_),
    .S(_2814_),
    .X(_2994_));
 sky130_fd_sc_hd__mux2_1 _3832_ (.A0(_2830_),
    .A1(_2820_),
    .S(_2814_),
    .X(_2995_));
 sky130_fd_sc_hd__mux2_1 _3833_ (.A0(_2994_),
    .A1(_2995_),
    .S(_1762_),
    .X(_2996_));
 sky130_fd_sc_hd__mux2_1 _3834_ (.A0(_2993_),
    .A1(_2996_),
    .S(_2839_),
    .X(_2997_));
 sky130_fd_sc_hd__nand2_1 _3835_ (.A(_2997_),
    .B(_2934_),
    .Y(_2998_));
 sky130_fd_sc_hd__or2_1 _3836_ (.A(_2840_),
    .B(_2823_),
    .X(_2999_));
 sky130_fd_sc_hd__o21a_1 _3837_ (.A1(_2120_),
    .A2(_2843_),
    .B1(_2999_),
    .X(_3000_));
 sky130_fd_sc_hd__nor2_1 _3838_ (.A(_2840_),
    .B(_2844_),
    .Y(_3001_));
 sky130_fd_sc_hd__nand2_1 _3839_ (.A(_3001_),
    .B(_2921_),
    .Y(_3002_));
 sky130_fd_sc_hd__o21ai_2 _3840_ (.A1(_2921_),
    .A2(_3000_),
    .B1(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__a21o_1 _3841_ (.A1(_3003_),
    .A2(_2941_),
    .B1(_2934_),
    .X(_3004_));
 sky130_fd_sc_hd__a32o_1 _3842_ (.A1(_2998_),
    .A2(_2838_),
    .A3(_3004_),
    .B1(net55),
    .B2(_2851_),
    .X(_3005_));
 sky130_fd_sc_hd__or2_1 _3843_ (.A(_2988_),
    .B(_3005_),
    .X(_3006_));
 sky130_fd_sc_hd__nand2_1 _3844_ (.A(_3005_),
    .B(_2988_),
    .Y(_3007_));
 sky130_fd_sc_hd__nand2_1 _3845_ (.A(_3006_),
    .B(_3007_),
    .Y(_3008_));
 sky130_fd_sc_hd__nor2_1 _3846_ (.A(_2969_),
    .B(_3008_),
    .Y(_3009_));
 sky130_fd_sc_hd__and2b_1 _3847_ (.A_N(_2920_),
    .B(_3009_),
    .X(_3010_));
 sky130_fd_sc_hd__nand2_1 _3848_ (.A(_2742_),
    .B(net1),
    .Y(_3011_));
 sky130_fd_sc_hd__nand2_1 _3849_ (.A(_2037_),
    .B(net12),
    .Y(_3012_));
 sky130_fd_sc_hd__mux2_1 _3850_ (.A0(_3011_),
    .A1(_3012_),
    .S(_2329_),
    .X(_3013_));
 sky130_fd_sc_hd__mux2_1 _3851_ (.A0(_3013_),
    .A1(_2972_),
    .S(_2758_),
    .X(_3014_));
 sky130_fd_sc_hd__mux2_1 _3852_ (.A0(_3014_),
    .A1(_2759_),
    .S(_1729_),
    .X(_3015_));
 sky130_fd_sc_hd__mux2_1 _3853_ (.A0(_2775_),
    .A1(_2750_),
    .S(_2760_),
    .X(_3016_));
 sky130_fd_sc_hd__mux2_1 _3854_ (.A0(_3015_),
    .A1(_3016_),
    .S(_1124_),
    .X(_3017_));
 sky130_fd_sc_hd__nand2_1 _3855_ (.A(_3017_),
    .B(_2779_),
    .Y(_3018_));
 sky130_fd_sc_hd__nand2_1 _3856_ (.A(_2788_),
    .B(_1729_),
    .Y(_3019_));
 sky130_fd_sc_hd__o21ai_1 _3857_ (.A1(_2951_),
    .A2(_2768_),
    .B1(_3019_),
    .Y(_3020_));
 sky130_fd_sc_hd__nand2_1 _3858_ (.A(_3020_),
    .B(_2873_),
    .Y(_3021_));
 sky130_fd_sc_hd__a21oi_1 _3859_ (.A1(_3021_),
    .A2(_2778_),
    .B1(_2794_),
    .Y(_3022_));
 sky130_fd_sc_hd__a22o_1 _3860_ (.A1(net1),
    .A2(_1674_),
    .B1(_3018_),
    .B2(_3022_),
    .X(_3023_));
 sky130_fd_sc_hd__inv_2 _3861_ (.A(_3023_),
    .Y(_3024_));
 sky130_fd_sc_hd__nand2_1 _3862_ (.A(_1927_),
    .B(net44),
    .Y(_3025_));
 sky130_fd_sc_hd__inv_2 _3863_ (.A(net33),
    .Y(_3026_));
 sky130_fd_sc_hd__or3_1 _3864_ (.A(_3026_),
    .B(_2329_),
    .C(_1905_),
    .X(_3027_));
 sky130_fd_sc_hd__o21a_1 _3865_ (.A1(_2441_),
    .A2(_3025_),
    .B1(_3027_),
    .X(_3028_));
 sky130_fd_sc_hd__mux2_1 _3866_ (.A0(_3028_),
    .A1(_2991_),
    .S(_2814_),
    .X(_3029_));
 sky130_fd_sc_hd__mux2_1 _3867_ (.A0(_3029_),
    .A1(_2815_),
    .S(_1762_),
    .X(_3030_));
 sky130_fd_sc_hd__mux2_1 _3868_ (.A0(_2831_),
    .A1(_2806_),
    .S(_2816_),
    .X(_3031_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(_3030_),
    .A1(_3031_),
    .S(_1245_),
    .X(_3032_));
 sky130_fd_sc_hd__nand2_1 _3870_ (.A(_3032_),
    .B(_2834_),
    .Y(_3033_));
 sky130_fd_sc_hd__nand2_1 _3871_ (.A(_2846_),
    .B(_2921_),
    .Y(_3034_));
 sky130_fd_sc_hd__o21ai_2 _3872_ (.A1(_2921_),
    .A2(_2824_),
    .B1(_3034_),
    .Y(_3035_));
 sky130_fd_sc_hd__a21o_1 _3873_ (.A1(_3035_),
    .A2(_2941_),
    .B1(_2834_),
    .X(_3036_));
 sky130_fd_sc_hd__nor2_1 _3874_ (.A(_3026_),
    .B(_2697_),
    .Y(_3037_));
 sky130_fd_sc_hd__a31o_1 _3875_ (.A1(_3033_),
    .A2(_2838_),
    .A3(_3036_),
    .B1(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__nor2_1 _3876_ (.A(_3024_),
    .B(_3038_),
    .Y(_3039_));
 sky130_fd_sc_hd__inv_2 _3877_ (.A(_3039_),
    .Y(_3040_));
 sky130_fd_sc_hd__nand2_1 _3878_ (.A(_3038_),
    .B(_3024_),
    .Y(_3041_));
 sky130_fd_sc_hd__and2_1 _3879_ (.A(_3040_),
    .B(_3041_),
    .X(_3042_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3880_ (.A(_3042_),
    .X(_3043_));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(_3000_),
    .A1(_2995_),
    .S(_2847_),
    .X(_3044_));
 sky130_fd_sc_hd__clkbuf_4 _3882_ (.A(_2941_),
    .X(_3045_));
 sky130_fd_sc_hd__nand2_1 _3883_ (.A(_3001_),
    .B(_2847_),
    .Y(_3046_));
 sky130_fd_sc_hd__or2_1 _3884_ (.A(_3045_),
    .B(_3046_),
    .X(_3047_));
 sky130_fd_sc_hd__o21ai_2 _3885_ (.A1(_2839_),
    .A2(_3044_),
    .B1(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__buf_2 _3886_ (.A(_2941_),
    .X(_3049_));
 sky130_fd_sc_hd__or3_1 _3887_ (.A(_2921_),
    .B(_2120_),
    .C(_3028_),
    .X(_3050_));
 sky130_fd_sc_hd__o21ai_1 _3888_ (.A1(_2847_),
    .A2(_2992_),
    .B1(_3050_),
    .Y(_3051_));
 sky130_fd_sc_hd__mux2_1 _3889_ (.A0(_2989_),
    .A1(_2994_),
    .S(_2921_),
    .X(_3052_));
 sky130_fd_sc_hd__nor2_1 _3890_ (.A(_3049_),
    .B(_3052_),
    .Y(_3053_));
 sky130_fd_sc_hd__a211o_1 _3891_ (.A1(_3049_),
    .A2(_3051_),
    .B1(_2177_),
    .C1(_3053_),
    .X(_3054_));
 sky130_fd_sc_hd__o211ai_4 _3892_ (.A1(_2934_),
    .A2(_3048_),
    .B1(_2838_),
    .C1(_3054_),
    .Y(_3055_));
 sky130_fd_sc_hd__nand2_1 _3893_ (.A(_2939_),
    .B(_2847_),
    .Y(_3056_));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(_2929_),
    .A1(_2938_),
    .S(_2921_),
    .X(_3057_));
 sky130_fd_sc_hd__nand2_1 _3895_ (.A(_3057_),
    .B(_3045_),
    .Y(_3058_));
 sky130_fd_sc_hd__o21ai_2 _3896_ (.A1(_3045_),
    .A2(_3056_),
    .B1(_3058_),
    .Y(_3059_));
 sky130_fd_sc_hd__mux2_1 _3897_ (.A0(_3025_),
    .A1(_2990_),
    .S(_2339_),
    .X(_3060_));
 sky130_fd_sc_hd__or4_1 _3898_ (.A(_3026_),
    .B(_2814_),
    .C(_2441_),
    .D(_1905_),
    .X(_3061_));
 sky130_fd_sc_hd__o21ai_1 _3899_ (.A1(_2120_),
    .A2(_3060_),
    .B1(_3061_),
    .Y(_3062_));
 sky130_fd_sc_hd__mux2_1 _3900_ (.A0(_2925_),
    .A1(_3062_),
    .S(_2847_),
    .X(_3063_));
 sky130_fd_sc_hd__mux2_1 _3901_ (.A0(_2926_),
    .A1(_2930_),
    .S(_2921_),
    .X(_3064_));
 sky130_fd_sc_hd__nor2_1 _3902_ (.A(_2941_),
    .B(_3064_),
    .Y(_3065_));
 sky130_fd_sc_hd__a211o_1 _3903_ (.A1(_3045_),
    .A2(_3063_),
    .B1(_2177_),
    .C1(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__o211ai_2 _3904_ (.A1(_2934_),
    .A2(_3059_),
    .B1(_2838_),
    .C1(_3066_),
    .Y(_3067_));
 sky130_fd_sc_hd__mux2_1 _3905_ (.A0(_2944_),
    .A1(_2957_),
    .S(_1729_),
    .X(_3068_));
 sky130_fd_sc_hd__nand2_1 _3906_ (.A(_2958_),
    .B(_2789_),
    .Y(_3069_));
 sky130_fd_sc_hd__mux2_1 _3907_ (.A0(_3068_),
    .A1(_3069_),
    .S(_1135_),
    .X(_3070_));
 sky130_fd_sc_hd__inv_2 _3908_ (.A(_3070_),
    .Y(_3071_));
 sky130_fd_sc_hd__mux2_1 _3909_ (.A0(_3012_),
    .A1(_2971_),
    .S(_2809_),
    .X(_3072_));
 sky130_fd_sc_hd__nand2_1 _3910_ (.A(_3072_),
    .B(_2782_),
    .Y(_3073_));
 sky130_fd_sc_hd__o21ai_1 _3911_ (.A1(_2441_),
    .A2(_3011_),
    .B1(_2090_),
    .Y(_3074_));
 sky130_fd_sc_hd__nor2_1 _3912_ (.A(_2789_),
    .B(_2949_),
    .Y(_3075_));
 sky130_fd_sc_hd__a31o_1 _3913_ (.A1(_2789_),
    .A2(_3073_),
    .A3(_3074_),
    .B1(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__mux2_1 _3914_ (.A0(_2950_),
    .A1(_2945_),
    .S(_1729_),
    .X(_3077_));
 sky130_fd_sc_hd__nor2_1 _3915_ (.A(_2961_),
    .B(_3077_),
    .Y(_3078_));
 sky130_fd_sc_hd__a211o_1 _3916_ (.A1(_3076_),
    .A2(_2961_),
    .B1(_2778_),
    .C1(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__o211ai_2 _3917_ (.A1(_2780_),
    .A2(_3071_),
    .B1(_2793_),
    .C1(_3079_),
    .Y(_3080_));
 sky130_fd_sc_hd__a21bo_1 _3918_ (.A1(_3055_),
    .A2(_3067_),
    .B1_N(_3080_),
    .X(_3081_));
 sky130_fd_sc_hd__nand2_1 _3919_ (.A(_3043_),
    .B(_3081_),
    .Y(_3082_));
 sky130_fd_sc_hd__nand2_1 _3920_ (.A(_3082_),
    .B(_3040_),
    .Y(_3083_));
 sky130_fd_sc_hd__mux2_1 _3921_ (.A0(_2864_),
    .A1(_2871_),
    .S(_2760_),
    .X(_3084_));
 sky130_fd_sc_hd__mux2_1 _3922_ (.A0(_2948_),
    .A1(_3072_),
    .S(_2090_),
    .X(_3085_));
 sky130_fd_sc_hd__mux2_1 _3923_ (.A0(_2868_),
    .A1(_3085_),
    .S(_2760_),
    .X(_3086_));
 sky130_fd_sc_hd__mux2_1 _3924_ (.A0(_3084_),
    .A1(_3086_),
    .S(_2873_),
    .X(_3087_));
 sky130_fd_sc_hd__nand2_1 _3925_ (.A(_3087_),
    .B(_2780_),
    .Y(_3088_));
 sky130_fd_sc_hd__nand2_1 _3926_ (.A(_2879_),
    .B(_2951_),
    .Y(_3089_));
 sky130_fd_sc_hd__o21ai_1 _3927_ (.A1(_2951_),
    .A2(_2860_),
    .B1(_3089_),
    .Y(_3090_));
 sky130_fd_sc_hd__nand2_1 _3928_ (.A(_3090_),
    .B(_2953_),
    .Y(_3091_));
 sky130_fd_sc_hd__a21oi_1 _3929_ (.A1(_3091_),
    .A2(_2778_),
    .B1(_2794_),
    .Y(_3092_));
 sky130_fd_sc_hd__a22o_1 _3930_ (.A1(net12),
    .A2(_2964_),
    .B1(_3088_),
    .B2(_3092_),
    .X(_3093_));
 sky130_fd_sc_hd__inv_2 _3931_ (.A(_3093_),
    .Y(_3094_));
 sky130_fd_sc_hd__mux2_1 _3932_ (.A0(_2923_),
    .A1(_3060_),
    .S(_2120_),
    .X(_3095_));
 sky130_fd_sc_hd__mux2_1 _3933_ (.A0(_2900_),
    .A1(_3095_),
    .S(_2816_),
    .X(_3096_));
 sky130_fd_sc_hd__mux2_1 _3934_ (.A0(_2904_),
    .A1(_2894_),
    .S(_1762_),
    .X(_3097_));
 sky130_fd_sc_hd__mux2_1 _3935_ (.A0(_3096_),
    .A1(_3097_),
    .S(_2839_),
    .X(_3098_));
 sky130_fd_sc_hd__nand2_1 _3936_ (.A(_3098_),
    .B(_2934_),
    .Y(_3099_));
 sky130_fd_sc_hd__mux2_1 _3937_ (.A0(_2912_),
    .A1(_2889_),
    .S(_2847_),
    .X(_3100_));
 sky130_fd_sc_hd__a21o_1 _3938_ (.A1(_3100_),
    .A2(_2941_),
    .B1(_2934_),
    .X(_3101_));
 sky130_fd_sc_hd__a32o_1 _3939_ (.A1(_3099_),
    .A2(_3101_),
    .A3(_2838_),
    .B1(net44),
    .B2(_2851_),
    .X(_3102_));
 sky130_fd_sc_hd__or2_1 _3940_ (.A(_3094_),
    .B(_3102_),
    .X(_3103_));
 sky130_fd_sc_hd__nand2_1 _3941_ (.A(_3102_),
    .B(_3094_),
    .Y(_3104_));
 sky130_fd_sc_hd__and2_1 _3942_ (.A(_3103_),
    .B(_3104_),
    .X(_3105_));
 sky130_fd_sc_hd__clkbuf_2 _3943_ (.A(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(_3083_),
    .B(_3106_),
    .Y(_3107_));
 sky130_fd_sc_hd__nand2_1 _3945_ (.A(_3107_),
    .B(_3103_),
    .Y(_3108_));
 sky130_fd_sc_hd__o21a_1 _3946_ (.A1(_2969_),
    .A2(_3006_),
    .B1(_2967_),
    .X(_3109_));
 sky130_fd_sc_hd__o21a_1 _3947_ (.A1(_2853_),
    .A2(_2919_),
    .B1(_2917_),
    .X(_3110_));
 sky130_fd_sc_hd__o21ai_1 _3948_ (.A1(_3109_),
    .A2(_2920_),
    .B1(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__a21o_1 _3949_ (.A1(_3010_),
    .A2(_3108_),
    .B1(_3111_),
    .X(_3112_));
 sky130_fd_sc_hd__nand2_1 _3950_ (.A(_2946_),
    .B(_2953_),
    .Y(_3113_));
 sky130_fd_sc_hd__or2_1 _3951_ (.A(_2953_),
    .B(_2960_),
    .X(_3114_));
 sky130_fd_sc_hd__nand2_2 _3952_ (.A(_2793_),
    .B(_2779_),
    .Y(_3115_));
 sky130_fd_sc_hd__inv_2 _3953_ (.A(_3115_),
    .Y(_3116_));
 sky130_fd_sc_hd__a32o_1 _3954_ (.A1(_3113_),
    .A2(_3114_),
    .A3(_3116_),
    .B1(net3),
    .B2(_2964_),
    .X(_3117_));
 sky130_fd_sc_hd__inv_2 _3955_ (.A(_3117_),
    .Y(_3118_));
 sky130_fd_sc_hd__or2_1 _3956_ (.A(_2941_),
    .B(_2940_),
    .X(_3119_));
 sky130_fd_sc_hd__nand2_2 _3957_ (.A(_2837_),
    .B(_2834_),
    .Y(_3120_));
 sky130_fd_sc_hd__inv_2 _3958_ (.A(_3120_),
    .Y(_3121_));
 sky130_fd_sc_hd__buf_2 _3959_ (.A(_3121_),
    .X(_3122_));
 sky130_fd_sc_hd__nand2_1 _3960_ (.A(_2932_),
    .B(_3045_),
    .Y(_3123_));
 sky130_fd_sc_hd__a32o_1 _3961_ (.A1(_3119_),
    .A2(_3122_),
    .A3(_3123_),
    .B1(net35),
    .B2(_2851_),
    .X(_3124_));
 sky130_fd_sc_hd__or2_1 _3962_ (.A(_3118_),
    .B(_3124_),
    .X(_3125_));
 sky130_fd_sc_hd__nand2_1 _3963_ (.A(_3124_),
    .B(_3118_),
    .Y(_3126_));
 sky130_fd_sc_hd__nand2_2 _3964_ (.A(_3125_),
    .B(_3126_),
    .Y(_3127_));
 sky130_fd_sc_hd__or2_1 _3965_ (.A(_2953_),
    .B(_2984_),
    .X(_3128_));
 sky130_fd_sc_hd__nand2_1 _3966_ (.A(_2977_),
    .B(_2961_),
    .Y(_3129_));
 sky130_fd_sc_hd__a32o_1 _3967_ (.A1(_3128_),
    .A2(_3129_),
    .A3(_3116_),
    .B1(net2),
    .B2(_2964_),
    .X(_3130_));
 sky130_fd_sc_hd__inv_2 _3968_ (.A(_3130_),
    .Y(_3131_));
 sky130_fd_sc_hd__or2_1 _3969_ (.A(_2941_),
    .B(_3003_),
    .X(_3132_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(_2996_),
    .B(_3049_),
    .Y(_3133_));
 sky130_fd_sc_hd__buf_2 _3971_ (.A(_2851_),
    .X(_3134_));
 sky130_fd_sc_hd__a32o_1 _3972_ (.A1(_3132_),
    .A2(_3133_),
    .A3(_3122_),
    .B1(net34),
    .B2(_3134_),
    .X(_3135_));
 sky130_fd_sc_hd__or2_1 _3973_ (.A(_3131_),
    .B(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__nand2_1 _3974_ (.A(_3135_),
    .B(_3131_),
    .Y(_3137_));
 sky130_fd_sc_hd__nand2_1 _3975_ (.A(_3136_),
    .B(_3137_),
    .Y(_3138_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(_3127_),
    .B(_3138_),
    .Y(_3139_));
 sky130_fd_sc_hd__nand2_1 _3977_ (.A(_2776_),
    .B(_2953_),
    .Y(_3140_));
 sky130_fd_sc_hd__a21oi_1 _3978_ (.A1(_2790_),
    .A2(_1135_),
    .B1(_3115_),
    .Y(_3141_));
 sky130_fd_sc_hd__a22o_1 _3979_ (.A1(net4),
    .A2(_2964_),
    .B1(_3140_),
    .B2(_3141_),
    .X(_3142_));
 sky130_fd_sc_hd__inv_2 _3980_ (.A(_3142_),
    .Y(_3143_));
 sky130_fd_sc_hd__nand2_1 _3981_ (.A(_2832_),
    .B(_3045_),
    .Y(_3144_));
 sky130_fd_sc_hd__nand2_1 _3982_ (.A(_2848_),
    .B(_2839_),
    .Y(_3145_));
 sky130_fd_sc_hd__a32o_1 _3983_ (.A1(_3144_),
    .A2(_3121_),
    .A3(_3145_),
    .B1(net36),
    .B2(_2851_),
    .X(_3146_));
 sky130_fd_sc_hd__or2_1 _3984_ (.A(_3143_),
    .B(_3146_),
    .X(_3147_));
 sky130_fd_sc_hd__nand2_1 _3985_ (.A(_3146_),
    .B(_3143_),
    .Y(_3148_));
 sky130_fd_sc_hd__nand2_1 _3986_ (.A(_3147_),
    .B(_3148_),
    .Y(_3149_));
 sky130_fd_sc_hd__nand2_1 _3987_ (.A(_2865_),
    .B(_2953_),
    .Y(_3150_));
 sky130_fd_sc_hd__a21oi_1 _3988_ (.A1(_2880_),
    .A2(_1135_),
    .B1(_3115_),
    .Y(_3151_));
 sky130_fd_sc_hd__a22o_1 _3989_ (.A1(net5),
    .A2(_2964_),
    .B1(_3150_),
    .B2(_3151_),
    .X(_3152_));
 sky130_fd_sc_hd__inv_2 _3990_ (.A(_3152_),
    .Y(_3153_));
 sky130_fd_sc_hd__nand2_1 _3991_ (.A(_2897_),
    .B(_2941_),
    .Y(_3154_));
 sky130_fd_sc_hd__nand2_1 _3992_ (.A(_2913_),
    .B(_2839_),
    .Y(_3155_));
 sky130_fd_sc_hd__a32o_1 _3993_ (.A1(_3154_),
    .A2(_3121_),
    .A3(_3155_),
    .B1(net37),
    .B2(_2851_),
    .X(_3156_));
 sky130_fd_sc_hd__or2_1 _3994_ (.A(_3153_),
    .B(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__nand2_1 _3995_ (.A(_3156_),
    .B(_3153_),
    .Y(_3158_));
 sky130_fd_sc_hd__nand2_2 _3996_ (.A(_3157_),
    .B(_3158_),
    .Y(_3159_));
 sky130_fd_sc_hd__nor2_1 _3997_ (.A(_3149_),
    .B(_3159_),
    .Y(_3160_));
 sky130_fd_sc_hd__nand2_1 _3998_ (.A(_3139_),
    .B(_3160_),
    .Y(_3161_));
 sky130_fd_sc_hd__mux2_1 _3999_ (.A0(_3077_),
    .A1(_3068_),
    .S(_1135_),
    .X(_3162_));
 sky130_fd_sc_hd__nand2_1 _4000_ (.A(_3162_),
    .B(_2780_),
    .Y(_3163_));
 sky130_fd_sc_hd__or2_1 _4001_ (.A(_1135_),
    .B(_3069_),
    .X(_3164_));
 sky130_fd_sc_hd__a21oi_1 _4002_ (.A1(_3164_),
    .A2(_2778_),
    .B1(_2794_),
    .Y(_3165_));
 sky130_fd_sc_hd__a22o_1 _4003_ (.A1(net30),
    .A2(_2964_),
    .B1(_3163_),
    .B2(_3165_),
    .X(_3166_));
 sky130_fd_sc_hd__inv_2 _4004_ (.A(_3166_),
    .Y(_3167_));
 sky130_fd_sc_hd__nand2_1 _4005_ (.A(_3064_),
    .B(_3045_),
    .Y(_3168_));
 sky130_fd_sc_hd__o21ai_1 _4006_ (.A1(_3045_),
    .A2(_3057_),
    .B1(_3168_),
    .Y(_3169_));
 sky130_fd_sc_hd__nand2_1 _4007_ (.A(_3169_),
    .B(_2934_),
    .Y(_3170_));
 sky130_fd_sc_hd__o21ai_1 _4008_ (.A1(_2839_),
    .A2(_3056_),
    .B1(_2177_),
    .Y(_3171_));
 sky130_fd_sc_hd__a32o_1 _4009_ (.A1(_3170_),
    .A2(_2838_),
    .A3(_3171_),
    .B1(net62),
    .B2(_3134_),
    .X(_3172_));
 sky130_fd_sc_hd__or2_1 _4010_ (.A(_3167_),
    .B(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__nand2_1 _4011_ (.A(_3172_),
    .B(_3167_),
    .Y(_3174_));
 sky130_fd_sc_hd__nand2_2 _4012_ (.A(_3173_),
    .B(_3174_),
    .Y(_3175_));
 sky130_fd_sc_hd__mux2_1 _4013_ (.A0(_2981_),
    .A1(_2976_),
    .S(_2789_),
    .X(_3176_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(_2970_),
    .A1(_2975_),
    .S(_2951_),
    .X(_3177_));
 sky130_fd_sc_hd__mux2_1 _4015_ (.A0(_3176_),
    .A1(_3177_),
    .S(_2961_),
    .X(_3178_));
 sky130_fd_sc_hd__nand2_1 _4016_ (.A(_3178_),
    .B(_2780_),
    .Y(_3179_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(_2982_),
    .B(_2789_),
    .Y(_3180_));
 sky130_fd_sc_hd__nor2_1 _4018_ (.A(_1135_),
    .B(_3180_),
    .Y(_3181_));
 sky130_fd_sc_hd__o21a_1 _4019_ (.A1(_2780_),
    .A2(_3181_),
    .B1(_2793_),
    .X(_3182_));
 sky130_fd_sc_hd__a22o_1 _4020_ (.A1(net29),
    .A2(_2965_),
    .B1(_3179_),
    .B2(_3182_),
    .X(_3183_));
 sky130_fd_sc_hd__inv_2 _4021_ (.A(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__mux2_1 _4022_ (.A0(_3044_),
    .A1(_3052_),
    .S(_3045_),
    .X(_3185_));
 sky130_fd_sc_hd__nand2_1 _4023_ (.A(_3185_),
    .B(_2934_),
    .Y(_3186_));
 sky130_fd_sc_hd__nor2_1 _4024_ (.A(_2839_),
    .B(_3046_),
    .Y(_3187_));
 sky130_fd_sc_hd__inv_2 _4025_ (.A(_3187_),
    .Y(_3188_));
 sky130_fd_sc_hd__nand2_1 _4026_ (.A(_3188_),
    .B(_2177_),
    .Y(_3189_));
 sky130_fd_sc_hd__a32o_1 _4027_ (.A1(_3186_),
    .A2(_2838_),
    .A3(_3189_),
    .B1(net61),
    .B2(_3134_),
    .X(_3190_));
 sky130_fd_sc_hd__or2_1 _4028_ (.A(_3184_),
    .B(_3190_),
    .X(_3191_));
 sky130_fd_sc_hd__nand2_1 _4029_ (.A(_3190_),
    .B(_3184_),
    .Y(_3192_));
 sky130_fd_sc_hd__nand2_1 _4030_ (.A(_3191_),
    .B(_3192_),
    .Y(_3193_));
 sky130_fd_sc_hd__nor2_1 _4031_ (.A(_3175_),
    .B(_3193_),
    .Y(_3194_));
 sky130_fd_sc_hd__nand2_1 _4032_ (.A(_3016_),
    .B(_2961_),
    .Y(_3195_));
 sky130_fd_sc_hd__or2_1 _4033_ (.A(_2953_),
    .B(_3020_),
    .X(_3196_));
 sky130_fd_sc_hd__a32o_1 _4034_ (.A1(_3195_),
    .A2(_3196_),
    .A3(_3116_),
    .B1(net31),
    .B2(_2965_),
    .X(_3197_));
 sky130_fd_sc_hd__inv_2 _4035_ (.A(_3197_),
    .Y(_3198_));
 sky130_fd_sc_hd__nand2_1 _4036_ (.A(_3031_),
    .B(_3049_),
    .Y(_3199_));
 sky130_fd_sc_hd__or2_1 _4037_ (.A(_3045_),
    .B(_3035_),
    .X(_3200_));
 sky130_fd_sc_hd__a32o_1 _4038_ (.A1(_3199_),
    .A2(_3200_),
    .A3(_3122_),
    .B1(net63),
    .B2(_3134_),
    .X(_3201_));
 sky130_fd_sc_hd__or2_1 _4039_ (.A(_3198_),
    .B(_3201_),
    .X(_3202_));
 sky130_fd_sc_hd__nand2_1 _4040_ (.A(_3201_),
    .B(_3198_),
    .Y(_3203_));
 sky130_fd_sc_hd__nand2_2 _4041_ (.A(_3202_),
    .B(_3203_),
    .Y(_3204_));
 sky130_fd_sc_hd__or2_1 _4042_ (.A(_2961_),
    .B(_3090_),
    .X(_3205_));
 sky130_fd_sc_hd__nand2_1 _4043_ (.A(_3084_),
    .B(_2961_),
    .Y(_3206_));
 sky130_fd_sc_hd__a32o_1 _4044_ (.A1(_3205_),
    .A2(_3206_),
    .A3(_3116_),
    .B1(net32),
    .B2(_2965_),
    .X(_3207_));
 sky130_fd_sc_hd__inv_2 _4045_ (.A(_3207_),
    .Y(_3208_));
 sky130_fd_sc_hd__or2_1 _4046_ (.A(_3049_),
    .B(_3100_),
    .X(_3209_));
 sky130_fd_sc_hd__nand2_1 _4047_ (.A(_3097_),
    .B(_3049_),
    .Y(_3210_));
 sky130_fd_sc_hd__a32o_1 _4048_ (.A1(_3209_),
    .A2(_3122_),
    .A3(_3210_),
    .B1(net64),
    .B2(_3134_),
    .X(_3211_));
 sky130_fd_sc_hd__or2_1 _4049_ (.A(_3208_),
    .B(_3211_),
    .X(_3212_));
 sky130_fd_sc_hd__nand2_1 _4050_ (.A(_3211_),
    .B(_3208_),
    .Y(_3213_));
 sky130_fd_sc_hd__nand2_2 _4051_ (.A(_3212_),
    .B(_3213_),
    .Y(_3214_));
 sky130_fd_sc_hd__nor2_1 _4052_ (.A(_3204_),
    .B(_3214_),
    .Y(_3215_));
 sky130_fd_sc_hd__nand2_1 _4053_ (.A(_3194_),
    .B(_3215_),
    .Y(_3216_));
 sky130_fd_sc_hd__nor2_1 _4054_ (.A(_3161_),
    .B(_3216_),
    .Y(_3217_));
 sky130_fd_sc_hd__o21ai_1 _4055_ (.A1(_3175_),
    .A2(_3191_),
    .B1(_3173_),
    .Y(_3218_));
 sky130_fd_sc_hd__o21ai_1 _4056_ (.A1(_3202_),
    .A2(_3214_),
    .B1(_3212_),
    .Y(_3219_));
 sky130_fd_sc_hd__a21o_1 _4057_ (.A1(_3218_),
    .A2(_3215_),
    .B1(_3219_),
    .X(_3220_));
 sky130_fd_sc_hd__inv_2 _4058_ (.A(_3161_),
    .Y(_3221_));
 sky130_fd_sc_hd__nand2_1 _4059_ (.A(_3220_),
    .B(_3221_),
    .Y(_3222_));
 sky130_fd_sc_hd__inv_2 _4060_ (.A(_3160_),
    .Y(_3223_));
 sky130_fd_sc_hd__o21a_1 _4061_ (.A1(_3136_),
    .A2(_3127_),
    .B1(_3125_),
    .X(_3224_));
 sky130_fd_sc_hd__o221a_1 _4062_ (.A1(_3159_),
    .A2(_3147_),
    .B1(_3223_),
    .B2(_3224_),
    .C1(_3157_),
    .X(_3225_));
 sky130_fd_sc_hd__nand2_1 _4063_ (.A(_3222_),
    .B(_3225_),
    .Y(_3226_));
 sky130_fd_sc_hd__a21o_1 _4064_ (.A1(_3112_),
    .A2(_3217_),
    .B1(_3226_),
    .X(_3227_));
 sky130_fd_sc_hd__o2bb2a_1 _4065_ (.A1_N(net11),
    .A2_N(_2965_),
    .B1(_3115_),
    .B2(_2962_),
    .X(_3228_));
 sky130_fd_sc_hd__a32o_1 _4066_ (.A1(_2940_),
    .A2(_3049_),
    .A3(_3122_),
    .B1(net43),
    .B2(_3134_),
    .X(_3229_));
 sky130_fd_sc_hd__or2_1 _4067_ (.A(_3228_),
    .B(_3229_),
    .X(_3230_));
 sky130_fd_sc_hd__nand2_1 _4068_ (.A(_3229_),
    .B(_3228_),
    .Y(_3231_));
 sky130_fd_sc_hd__nand2_2 _4069_ (.A(_3230_),
    .B(_3231_),
    .Y(_3232_));
 sky130_fd_sc_hd__o2bb2a_1 _4070_ (.A1_N(net10),
    .A2_N(_2965_),
    .B1(_3115_),
    .B2(_2985_),
    .X(_3233_));
 sky130_fd_sc_hd__a32o_1 _4071_ (.A1(_3003_),
    .A2(_3049_),
    .A3(_3122_),
    .B1(net42),
    .B2(_3134_),
    .X(_3234_));
 sky130_fd_sc_hd__or2_1 _4072_ (.A(_3233_),
    .B(_3234_),
    .X(_3235_));
 sky130_fd_sc_hd__nand2_1 _4073_ (.A(_3234_),
    .B(_3233_),
    .Y(_3236_));
 sky130_fd_sc_hd__nand2_2 _4074_ (.A(_3235_),
    .B(_3236_),
    .Y(_3237_));
 sky130_fd_sc_hd__nor2_1 _4075_ (.A(_3232_),
    .B(_3237_),
    .Y(_3238_));
 sky130_fd_sc_hd__inv_2 _4076_ (.A(net13),
    .Y(_3239_));
 sky130_fd_sc_hd__o22a_1 _4077_ (.A1(_3239_),
    .A2(_1685_),
    .B1(_3115_),
    .B2(_2791_),
    .X(_3240_));
 sky130_fd_sc_hd__inv_2 _4078_ (.A(net45),
    .Y(_3241_));
 sky130_fd_sc_hd__o22a_1 _4079_ (.A1(_3241_),
    .A2(_2697_),
    .B1(_3120_),
    .B2(_2849_),
    .X(_3242_));
 sky130_fd_sc_hd__inv_2 _4080_ (.A(_3242_),
    .Y(_3243_));
 sky130_fd_sc_hd__or2_1 _4081_ (.A(_3240_),
    .B(_3243_),
    .X(_3244_));
 sky130_fd_sc_hd__nand2_1 _4082_ (.A(_3243_),
    .B(_3240_),
    .Y(_3245_));
 sky130_fd_sc_hd__nand2_1 _4083_ (.A(_3244_),
    .B(_3245_),
    .Y(_3246_));
 sky130_fd_sc_hd__o22a_1 _4084_ (.A1(_2705_),
    .A2(_1685_),
    .B1(_3115_),
    .B2(_2881_),
    .X(_3247_));
 sky130_fd_sc_hd__o22a_1 _4085_ (.A1(_2686_),
    .A2(_2697_),
    .B1(_3120_),
    .B2(_2914_),
    .X(_3248_));
 sky130_fd_sc_hd__inv_2 _4086_ (.A(_3248_),
    .Y(_3249_));
 sky130_fd_sc_hd__or2_1 _4087_ (.A(_3247_),
    .B(_3249_),
    .X(_3250_));
 sky130_fd_sc_hd__nand2_1 _4088_ (.A(_3249_),
    .B(_3247_),
    .Y(_3251_));
 sky130_fd_sc_hd__nand2_2 _4089_ (.A(_3250_),
    .B(_3251_),
    .Y(_3252_));
 sky130_fd_sc_hd__nor2_1 _4090_ (.A(_3246_),
    .B(_3252_),
    .Y(_3253_));
 sky130_fd_sc_hd__nand2_1 _4091_ (.A(_3238_),
    .B(_3253_),
    .Y(_3254_));
 sky130_fd_sc_hd__o2bb2a_1 _4092_ (.A1_N(net8),
    .A2_N(_2964_),
    .B1(_3115_),
    .B2(_3021_),
    .X(_3255_));
 sky130_fd_sc_hd__a32o_1 _4093_ (.A1(_3035_),
    .A2(_3049_),
    .A3(_3122_),
    .B1(net40),
    .B2(_2851_),
    .X(_3256_));
 sky130_fd_sc_hd__or2_1 _4094_ (.A(_3255_),
    .B(_3256_),
    .X(_3257_));
 sky130_fd_sc_hd__nand2_1 _4095_ (.A(_3256_),
    .B(_3255_),
    .Y(_3258_));
 sky130_fd_sc_hd__nand2_2 _4096_ (.A(_3257_),
    .B(_3258_),
    .Y(_3259_));
 sky130_fd_sc_hd__o2bb2a_1 _4097_ (.A1_N(net9),
    .A2_N(_2965_),
    .B1(_3115_),
    .B2(_3091_),
    .X(_3260_));
 sky130_fd_sc_hd__a32o_1 _4098_ (.A1(_3100_),
    .A2(_3049_),
    .A3(_3122_),
    .B1(net41),
    .B2(_2851_),
    .X(_3261_));
 sky130_fd_sc_hd__or2_1 _4099_ (.A(_3260_),
    .B(_3261_),
    .X(_3262_));
 sky130_fd_sc_hd__nand2_1 _4100_ (.A(_3261_),
    .B(_3260_),
    .Y(_3263_));
 sky130_fd_sc_hd__nand2_2 _4101_ (.A(_3262_),
    .B(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__nor2_1 _4102_ (.A(_3259_),
    .B(_3264_),
    .Y(_3265_));
 sky130_fd_sc_hd__a22o_1 _4103_ (.A1(net7),
    .A2(_2964_),
    .B1(_3071_),
    .B2(_3116_),
    .X(_3266_));
 sky130_fd_sc_hd__inv_2 _4104_ (.A(_3266_),
    .Y(_3267_));
 sky130_fd_sc_hd__a22o_1 _4105_ (.A1(net39),
    .A2(_3134_),
    .B1(_3059_),
    .B2(_3122_),
    .X(_3268_));
 sky130_fd_sc_hd__or2_1 _4106_ (.A(_3267_),
    .B(_3268_),
    .X(_3269_));
 sky130_fd_sc_hd__nand2_1 _4107_ (.A(_3268_),
    .B(_3267_),
    .Y(_3270_));
 sky130_fd_sc_hd__nand2_2 _4108_ (.A(_3269_),
    .B(_3270_),
    .Y(_3271_));
 sky130_fd_sc_hd__mux2_1 _4109_ (.A0(_3176_),
    .A1(_3180_),
    .S(_1135_),
    .X(_3272_));
 sky130_fd_sc_hd__inv_2 _4110_ (.A(_3272_),
    .Y(_3273_));
 sky130_fd_sc_hd__a22o_1 _4111_ (.A1(net6),
    .A2(_2965_),
    .B1(_3273_),
    .B2(_3116_),
    .X(_3274_));
 sky130_fd_sc_hd__inv_2 _4112_ (.A(_3274_),
    .Y(_3275_));
 sky130_fd_sc_hd__a22o_1 _4113_ (.A1(net38),
    .A2(_3134_),
    .B1(_3048_),
    .B2(_3122_),
    .X(_3276_));
 sky130_fd_sc_hd__or2_1 _4114_ (.A(_3275_),
    .B(_3276_),
    .X(_3277_));
 sky130_fd_sc_hd__nand2_1 _4115_ (.A(_3276_),
    .B(_3275_),
    .Y(_3278_));
 sky130_fd_sc_hd__nand2_1 _4116_ (.A(_3277_),
    .B(_3278_),
    .Y(_3279_));
 sky130_fd_sc_hd__nor2_1 _4117_ (.A(_3271_),
    .B(_3279_),
    .Y(_3280_));
 sky130_fd_sc_hd__nand2_1 _4118_ (.A(_3265_),
    .B(_3280_),
    .Y(_3281_));
 sky130_fd_sc_hd__nor2_1 _4119_ (.A(_3254_),
    .B(_3281_),
    .Y(_3282_));
 sky130_fd_sc_hd__nand2_1 _4120_ (.A(_3227_),
    .B(_3282_),
    .Y(_3283_));
 sky130_fd_sc_hd__inv_2 _4121_ (.A(_3253_),
    .Y(_3284_));
 sky130_fd_sc_hd__o21a_1 _4122_ (.A1(_3235_),
    .A2(_3232_),
    .B1(_3230_),
    .X(_3285_));
 sky130_fd_sc_hd__inv_2 _4123_ (.A(_3265_),
    .Y(_3286_));
 sky130_fd_sc_hd__o21a_1 _4124_ (.A1(_3277_),
    .A2(_3271_),
    .B1(_3269_),
    .X(_3287_));
 sky130_fd_sc_hd__o221a_1 _4125_ (.A1(_3264_),
    .A2(_3257_),
    .B1(_3286_),
    .B2(_3287_),
    .C1(_3262_),
    .X(_3288_));
 sky130_fd_sc_hd__o21a_1 _4126_ (.A1(_3244_),
    .A2(_3252_),
    .B1(_3250_),
    .X(_3289_));
 sky130_fd_sc_hd__o221a_1 _4127_ (.A1(_3284_),
    .A2(_3285_),
    .B1(_3254_),
    .B2(_3288_),
    .C1(_3289_),
    .X(_3290_));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(_3283_),
    .B(_3290_),
    .Y(_3291_));
 sky130_fd_sc_hd__a22o_1 _4129_ (.A1(net15),
    .A2(_2965_),
    .B1(_3181_),
    .B2(_3116_),
    .X(_3292_));
 sky130_fd_sc_hd__inv_2 _4130_ (.A(net47),
    .Y(_3293_));
 sky130_fd_sc_hd__o22a_1 _4131_ (.A1(_3293_),
    .A2(_2697_),
    .B1(_3120_),
    .B2(_3188_),
    .X(_3294_));
 sky130_fd_sc_hd__or2_1 _4132_ (.A(_3292_),
    .B(_3294_),
    .X(_3295_));
 sky130_fd_sc_hd__nand2_1 _4133_ (.A(_3294_),
    .B(_3292_),
    .Y(_3296_));
 sky130_fd_sc_hd__nand2_1 _4134_ (.A(_3295_),
    .B(_3296_),
    .Y(_3297_));
 sky130_fd_sc_hd__nor2_1 _4135_ (.A(_1652_),
    .B(_3297_),
    .Y(_3298_));
 sky130_fd_sc_hd__nand2_1 _4136_ (.A(_3291_),
    .B(_3298_),
    .Y(_3299_));
 sky130_fd_sc_hd__o21a_1 _4137_ (.A1(_1652_),
    .A2(_3296_),
    .B1(_3134_),
    .X(_3300_));
 sky130_fd_sc_hd__nand2_2 _4138_ (.A(_3299_),
    .B(_3300_),
    .Y(_3301_));
 sky130_fd_sc_hd__inv_2 _4139_ (.A(net25),
    .Y(_3302_));
 sky130_fd_sc_hd__nand2_1 _4140_ (.A(_3301_),
    .B(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__or3_1 _4141_ (.A(_2951_),
    .B(_2090_),
    .C(_3013_),
    .X(_3304_));
 sky130_fd_sc_hd__o21ai_1 _4142_ (.A1(_2789_),
    .A2(_2973_),
    .B1(_3304_),
    .Y(_3305_));
 sky130_fd_sc_hd__nor2_1 _4143_ (.A(_2961_),
    .B(_3177_),
    .Y(_3306_));
 sky130_fd_sc_hd__a211o_1 _4144_ (.A1(_2961_),
    .A2(_3305_),
    .B1(_2778_),
    .C1(_3306_),
    .X(_3307_));
 sky130_fd_sc_hd__o211ai_2 _4145_ (.A1(_2780_),
    .A2(_3273_),
    .B1(_2793_),
    .C1(_3307_),
    .Y(_3308_));
 sky130_fd_sc_hd__a21bo_1 _4146_ (.A1(_3080_),
    .A2(_3308_),
    .B1_N(_3067_),
    .X(_3309_));
 sky130_fd_sc_hd__a21bo_1 _4147_ (.A1(_3040_),
    .A2(_3309_),
    .B1_N(_3041_),
    .X(_3310_));
 sky130_fd_sc_hd__a21bo_1 _4148_ (.A1(_3310_),
    .A2(_3103_),
    .B1_N(_3104_),
    .X(_3311_));
 sky130_fd_sc_hd__o21a_1 _4149_ (.A1(_3007_),
    .A2(_2969_),
    .B1(_2968_),
    .X(_0036_));
 sky130_fd_sc_hd__o21a_1 _4150_ (.A1(_2854_),
    .A2(_2919_),
    .B1(_2918_),
    .X(_0037_));
 sky130_fd_sc_hd__o21ai_1 _4151_ (.A1(_0036_),
    .A2(_2920_),
    .B1(_0037_),
    .Y(_0038_));
 sky130_fd_sc_hd__a21o_1 _4152_ (.A1(_3010_),
    .A2(_3311_),
    .B1(_0038_),
    .X(_0039_));
 sky130_fd_sc_hd__nand2_1 _4153_ (.A(_0039_),
    .B(_3217_),
    .Y(_0040_));
 sky130_fd_sc_hd__o21a_1 _4154_ (.A1(_3192_),
    .A2(_3175_),
    .B1(_3174_),
    .X(_0041_));
 sky130_fd_sc_hd__o21a_1 _4155_ (.A1(_3203_),
    .A2(_3214_),
    .B1(_3213_),
    .X(_0042_));
 sky130_fd_sc_hd__o31ai_1 _4156_ (.A1(_3214_),
    .A2(_3204_),
    .A3(_0041_),
    .B1(_0042_),
    .Y(_0043_));
 sky130_fd_sc_hd__nand2_1 _4157_ (.A(_0043_),
    .B(_3221_),
    .Y(_0044_));
 sky130_fd_sc_hd__o21a_1 _4158_ (.A1(_3137_),
    .A2(_3127_),
    .B1(_3126_),
    .X(_0045_));
 sky130_fd_sc_hd__o221a_1 _4159_ (.A1(_3159_),
    .A2(_3148_),
    .B1(_3223_),
    .B2(_0045_),
    .C1(_3158_),
    .X(_0046_));
 sky130_fd_sc_hd__nand3_2 _4160_ (.A(_0040_),
    .B(_0044_),
    .C(_0046_),
    .Y(_0047_));
 sky130_fd_sc_hd__nand2_1 _4161_ (.A(_0047_),
    .B(_3282_),
    .Y(_0048_));
 sky130_fd_sc_hd__o21a_1 _4162_ (.A1(_3236_),
    .A2(_3232_),
    .B1(_3231_),
    .X(_0049_));
 sky130_fd_sc_hd__o21a_1 _4163_ (.A1(_3278_),
    .A2(_3271_),
    .B1(_3270_),
    .X(_0050_));
 sky130_fd_sc_hd__o221a_1 _4164_ (.A1(_3264_),
    .A2(_3258_),
    .B1(_3286_),
    .B2(_0050_),
    .C1(_3263_),
    .X(_0051_));
 sky130_fd_sc_hd__o21a_1 _4165_ (.A1(_3245_),
    .A2(_3252_),
    .B1(_3251_),
    .X(_0052_));
 sky130_fd_sc_hd__o221a_1 _4166_ (.A1(_3284_),
    .A2(_0049_),
    .B1(_3254_),
    .B2(_0051_),
    .C1(_0052_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_1 _4167_ (.A(_0048_),
    .B(_0053_),
    .Y(_0054_));
 sky130_fd_sc_hd__nand2_1 _4168_ (.A(_0054_),
    .B(_3298_),
    .Y(_0055_));
 sky130_fd_sc_hd__o21ai_1 _4169_ (.A1(_1652_),
    .A2(_3295_),
    .B1(_2965_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _4170_ (.A(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__nand2_4 _4171_ (.A(_0055_),
    .B(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _4172_ (.A(net57),
    .Y(_0059_));
 sky130_fd_sc_hd__nand2_1 _4173_ (.A(_0058_),
    .B(_0059_),
    .Y(_0060_));
 sky130_fd_sc_hd__nand2_1 _4174_ (.A(_3303_),
    .B(_0060_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _4175_ (.A(net65),
    .Y(_0062_));
 sky130_fd_sc_hd__and3_1 _4176_ (.A(_2737_),
    .B(_0062_),
    .C(net66),
    .X(_0063_));
 sky130_fd_sc_hd__nand2_2 _4177_ (.A(_0061_),
    .B(_0063_),
    .Y(_0064_));
 sky130_fd_sc_hd__and3_1 _4178_ (.A(_2737_),
    .B(net66),
    .C(net65),
    .X(_0065_));
 sky130_fd_sc_hd__nand3_2 _4179_ (.A(_3303_),
    .B(_0060_),
    .C(_0065_),
    .Y(_0066_));
 sky130_fd_sc_hd__nand2_8 _4180_ (.A(_0064_),
    .B(_0066_),
    .Y(_0067_));
 sky130_fd_sc_hd__nor2_1 _4181_ (.A(_0893_),
    .B(net131),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _4182_ (.A(net132),
    .Y(_0069_));
 sky130_fd_sc_hd__nand2_2 _4183_ (.A(_0067_),
    .B(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__nand2_1 _4184_ (.A(_2741_),
    .B(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(_0071_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand2_1 _4186_ (.A(_2738_),
    .B(_0062_),
    .Y(_0073_));
 sky130_fd_sc_hd__or2_4 _4187_ (.A(_2737_),
    .B(_0073_),
    .X(_0074_));
 sky130_fd_sc_hd__nor2_4 _4188_ (.A(_0074_),
    .B(net138),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _4189_ (.A(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__nand2_2 _4190_ (.A(_0072_),
    .B(_0076_),
    .Y(_0077_));
 sky130_fd_sc_hd__buf_4 _4191_ (.A(_0077_),
    .X(_0078_));
 sky130_fd_sc_hd__clkbuf_4 _4192_ (.A(_1696_),
    .X(_0079_));
 sky130_fd_sc_hd__o31a_1 _4193_ (.A1(_0893_),
    .A2(_2717_),
    .A3(_0078_),
    .B1(_0079_),
    .X(_0000_));
 sky130_fd_sc_hd__nand2_1 _4194_ (.A(net119),
    .B(net116),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _4195_ (.A(net117),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _4196_ (.A(_0077_),
    .Y(_0081_));
 sky130_fd_sc_hd__nand2_1 _4197_ (.A(_1663_),
    .B(net16),
    .Y(_0082_));
 sky130_fd_sc_hd__clkbuf_4 _4198_ (.A(_0805_),
    .X(_0083_));
 sky130_fd_sc_hd__nand3_2 _4199_ (.A(_1608_),
    .B(net48),
    .C(_1652_),
    .Y(_0084_));
 sky130_fd_sc_hd__nand3_2 _4200_ (.A(_0082_),
    .B(_0083_),
    .C(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _4201_ (.A(_0085_),
    .Y(_0086_));
 sky130_fd_sc_hd__nand2_1 _4202_ (.A(_1663_),
    .B(_0992_),
    .Y(_0087_));
 sky130_fd_sc_hd__nand3_1 _4203_ (.A(_1608_),
    .B(_0970_),
    .C(_1652_),
    .Y(_0088_));
 sky130_fd_sc_hd__nand2_4 _4204_ (.A(_0087_),
    .B(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__nand2_1 _4205_ (.A(_1663_),
    .B(_1080_),
    .Y(_0090_));
 sky130_fd_sc_hd__o21ai_4 _4206_ (.A1(net50),
    .A2(_1663_),
    .B1(_0090_),
    .Y(_0091_));
 sky130_fd_sc_hd__nand3_2 _4207_ (.A(_0086_),
    .B(_0089_),
    .C(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _4208_ (.A(_1663_),
    .B(_1157_),
    .Y(_0093_));
 sky130_fd_sc_hd__nand3_1 _4209_ (.A(_1608_),
    .B(_1014_),
    .C(_1652_),
    .Y(_0094_));
 sky130_fd_sc_hd__nand2_2 _4210_ (.A(_0093_),
    .B(_0094_),
    .Y(_0095_));
 sky130_fd_sc_hd__nand3_1 _4211_ (.A(_0089_),
    .B(_0095_),
    .C(_0083_),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _4212_ (.A(_0091_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _4213_ (.A(_0096_),
    .B(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__nand2_1 _4214_ (.A(_0092_),
    .B(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__nand2_1 _4215_ (.A(_0082_),
    .B(_0084_),
    .Y(_0100_));
 sky130_fd_sc_hd__nand2_1 _4216_ (.A(_0089_),
    .B(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__nor2_1 _4217_ (.A(_2719_),
    .B(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _4218_ (.A(_0102_),
    .Y(_0103_));
 sky130_fd_sc_hd__nand2_1 _4219_ (.A(_0099_),
    .B(_0103_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand3_2 _4220_ (.A(_0092_),
    .B(_0098_),
    .C(_0102_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2_1 _4221_ (.A(_0104_),
    .B(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ai_1 _4222_ (.A1(_0706_),
    .A2(_0816_),
    .B1(_0100_),
    .Y(_0107_));
 sky130_fd_sc_hd__nor2_1 _4223_ (.A(_0695_),
    .B(_0816_),
    .Y(_0108_));
 sky130_fd_sc_hd__nand2_1 _4224_ (.A(_0095_),
    .B(_0108_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand3_1 _4225_ (.A(_0107_),
    .B(_2725_),
    .C(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__nand2_1 _4226_ (.A(_0085_),
    .B(_2719_),
    .Y(_0111_));
 sky130_fd_sc_hd__nand2_1 _4227_ (.A(_0111_),
    .B(_0089_),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _4228_ (.A(_0089_),
    .Y(_0113_));
 sky130_fd_sc_hd__nand3_1 _4229_ (.A(_0085_),
    .B(_0113_),
    .C(_2719_),
    .Y(_0114_));
 sky130_fd_sc_hd__nand2_2 _4230_ (.A(_0112_),
    .B(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__nor2_1 _4231_ (.A(_0110_),
    .B(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _4232_ (.A(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__nand2_1 _4233_ (.A(_0106_),
    .B(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__nand3_2 _4234_ (.A(_0104_),
    .B(_0116_),
    .C(_0105_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_1 _4235_ (.A(_0118_),
    .B(_0119_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand2_1 _4236_ (.A(_0107_),
    .B(_0109_),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _4237_ (.A(net147),
    .Y(_0122_));
 sky130_fd_sc_hd__buf_6 _4238_ (.A(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__nand2_1 _4239_ (.A(_0121_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__nor2_1 _4240_ (.A(_0124_),
    .B(_0115_),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _4241_ (.A(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_2 _4242_ (.A(_0120_),
    .B(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__or2_1 _4243_ (.A(_0871_),
    .B(_2730_),
    .X(_0128_));
 sky130_fd_sc_hd__inv_2 _4244_ (.A(_0128_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_1 _4245_ (.A(_0121_),
    .B(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand3_1 _4246_ (.A(_0107_),
    .B(_0109_),
    .C(_0128_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand2_1 _4247_ (.A(_0130_),
    .B(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__mux2_1 _4248_ (.A0(\M000[22] ),
    .A1(net171),
    .S(_0684_),
    .X(_0133_));
 sky130_fd_sc_hd__or2_1 _4249_ (.A(_2718_),
    .B(net172),
    .X(_0134_));
 sky130_fd_sc_hd__o21ai_1 _4250_ (.A1(_0761_),
    .A2(_2728_),
    .B1(_0134_),
    .Y(_0135_));
 sky130_fd_sc_hd__mux2_2 _4251_ (.A0(_0135_),
    .A1(net146),
    .S(_0860_),
    .X(_0136_));
 sky130_fd_sc_hd__nand2_4 _4252_ (.A(_0136_),
    .B(_0122_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _4253_ (.A(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__buf_6 _4254_ (.A(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(_0132_),
    .B(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _4256_ (.A(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__nand3_2 _4257_ (.A(_0115_),
    .B(_0124_),
    .C(_0110_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _4258_ (.A(_0124_),
    .B(_0110_),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _4259_ (.A(_0115_),
    .Y(_0144_));
 sky130_fd_sc_hd__nand2_1 _4260_ (.A(_0143_),
    .B(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__nand3_4 _4261_ (.A(_0141_),
    .B(_0142_),
    .C(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _4262_ (.A(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__nand2_1 _4263_ (.A(_0127_),
    .B(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__nand3_4 _4264_ (.A(_0118_),
    .B(_0119_),
    .C(_0125_),
    .Y(_0149_));
 sky130_fd_sc_hd__nand2_1 _4265_ (.A(_0148_),
    .B(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nor2_1 _4266_ (.A(_0103_),
    .B(_0099_),
    .Y(_0151_));
 sky130_fd_sc_hd__nand2_1 _4267_ (.A(_1663_),
    .B(_0904_),
    .Y(_0152_));
 sky130_fd_sc_hd__o21ai_2 _4268_ (.A1(net51),
    .A2(_1663_),
    .B1(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _4269_ (.A(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__nand2_1 _4270_ (.A(_0092_),
    .B(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _4271_ (.A(_0096_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand2_1 _4272_ (.A(_0153_),
    .B(_0091_),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _4273_ (.A(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__nand2_1 _4274_ (.A(_0156_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__nand2_1 _4275_ (.A(_0155_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__nand2_1 _4276_ (.A(_0151_),
    .B(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__nor2_1 _4277_ (.A(_0157_),
    .B(_0096_),
    .Y(_0162_));
 sky130_fd_sc_hd__a21oi_1 _4278_ (.A1(_0092_),
    .A2(_0154_),
    .B1(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand2_1 _4279_ (.A(_0163_),
    .B(_0105_),
    .Y(_0164_));
 sky130_fd_sc_hd__nand3_1 _4280_ (.A(_0119_),
    .B(_0161_),
    .C(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand2_1 _4281_ (.A(_0164_),
    .B(_0161_),
    .Y(_0166_));
 sky130_fd_sc_hd__nor2_1 _4282_ (.A(_0117_),
    .B(_0106_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand2_2 _4283_ (.A(_0166_),
    .B(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2_2 _4284_ (.A(_0165_),
    .B(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_1 _4285_ (.A(_0150_),
    .B(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _4286_ (.A(_0169_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand3_1 _4287_ (.A(_0171_),
    .B(_0148_),
    .C(_0149_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _4288_ (.A(_0170_),
    .B(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _4289_ (.A(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__nand2_1 _4290_ (.A(_0127_),
    .B(_0149_),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_2 _4291_ (.A(_0175_),
    .B(_0146_),
    .Y(_0176_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(\M000[21] ),
    .A1(\M000[22] ),
    .S(_0684_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(net172),
    .A1(_0177_),
    .S(_0761_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _4294_ (.A(net173),
    .B(_0849_),
    .Y(_0179_));
 sky130_fd_sc_hd__o21ai_2 _4295_ (.A1(_0849_),
    .A2(_0135_),
    .B1(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _4296_ (.A(net174),
    .Y(_0181_));
 sky130_fd_sc_hd__nand3_2 _4297_ (.A(_0136_),
    .B(_0123_),
    .C(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__buf_2 _4298_ (.A(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_4 _4299_ (.A(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__buf_4 _4300_ (.A(_0139_),
    .X(_0185_));
 sky130_fd_sc_hd__xor2_1 _4301_ (.A(_0185_),
    .B(_0132_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_0145_),
    .B(_0142_),
    .Y(_0187_));
 sky130_fd_sc_hd__nand2_1 _4303_ (.A(_0187_),
    .B(_0140_),
    .Y(_0188_));
 sky130_fd_sc_hd__nand3_1 _4304_ (.A(_0146_),
    .B(_0186_),
    .C(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _4305_ (.A(_0184_),
    .B(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__nand3_4 _4306_ (.A(_0127_),
    .B(_0149_),
    .C(_0147_),
    .Y(_0191_));
 sky130_fd_sc_hd__nand3_2 _4307_ (.A(_0176_),
    .B(_0190_),
    .C(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _4308_ (.A(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_1 _4309_ (.A(_0174_),
    .B(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _4310_ (.A(_0173_),
    .B(_0192_),
    .Y(_0195_));
 sky130_fd_sc_hd__nand2_1 _4311_ (.A(_0194_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _4312_ (.A(_0132_),
    .Y(_0197_));
 sky130_fd_sc_hd__clkbuf_4 _4313_ (.A(_0137_),
    .X(_0198_));
 sky130_fd_sc_hd__nand2_1 _4314_ (.A(_0197_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _4315_ (.A(_0199_),
    .B(_0140_),
    .Y(_0200_));
 sky130_fd_sc_hd__nand2_1 _4316_ (.A(_0178_),
    .B(_0860_),
    .Y(_0201_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_0083_),
    .B(net164),
    .Y(_0202_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(_0684_),
    .B(\M000[21] ),
    .Y(_0203_));
 sky130_fd_sc_hd__and2_1 _4319_ (.A(_0202_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(_0177_),
    .B(_2718_),
    .Y(_0205_));
 sky130_fd_sc_hd__o21ai_1 _4321_ (.A1(_2718_),
    .A2(net165),
    .B1(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(net166),
    .B(_0849_),
    .Y(_0207_));
 sky130_fd_sc_hd__nand2_1 _4323_ (.A(_0201_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _4324_ (.A(net167),
    .Y(_0209_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(_0209_),
    .B(_0122_),
    .Y(_0210_));
 sky130_fd_sc_hd__o21ai_1 _4326_ (.A1(_0122_),
    .A2(_0180_),
    .B1(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__or2_1 _4327_ (.A(_0137_),
    .B(net168),
    .X(_0212_));
 sky130_fd_sc_hd__a21o_1 _4328_ (.A1(_0181_),
    .A2(_0123_),
    .B1(_0136_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _4329_ (.A(_0212_),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__inv_2 _4330_ (.A(net175),
    .Y(_0215_));
 sky130_fd_sc_hd__buf_2 _4331_ (.A(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__nand3_1 _4332_ (.A(_0200_),
    .B(_0214_),
    .C(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(_0146_),
    .B(_0188_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_0136_),
    .B(_2732_),
    .Y(_0219_));
 sky130_fd_sc_hd__o21ai_2 _4335_ (.A1(_2732_),
    .A2(_0180_),
    .B1(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__nand3_2 _4336_ (.A(_0197_),
    .B(_0185_),
    .C(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_0218_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__nand3b_2 _4338_ (.A_N(_0221_),
    .B(_0146_),
    .C(_0188_),
    .Y(_0223_));
 sky130_fd_sc_hd__nand3b_2 _4339_ (.A_N(_0217_),
    .B(_0222_),
    .C(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _4340_ (.A(_0176_),
    .B(_0191_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand2_1 _4341_ (.A(_0225_),
    .B(_0223_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand3b_1 _4342_ (.A_N(_0224_),
    .B(_0226_),
    .C(_0192_),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _4343_ (.A(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_2 _4344_ (.A(_0196_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_2 _4345_ (.A(_0223_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand3_2 _4346_ (.A(_0176_),
    .B(_0191_),
    .C(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__nand3_1 _4347_ (.A(_0231_),
    .B(_0170_),
    .C(_0172_),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _4348_ (.A(_0231_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _4349_ (.A(_0233_),
    .B(_0173_),
    .Y(_0234_));
 sky130_fd_sc_hd__nand2_1 _4350_ (.A(_0232_),
    .B(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand3_2 _4351_ (.A(_0220_),
    .B(_0139_),
    .C(net168),
    .Y(_0236_));
 sky130_fd_sc_hd__clkbuf_4 _4352_ (.A(net169),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _4353_ (.A(_0218_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _4354_ (.A(_0200_),
    .B(_0183_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand3_1 _4355_ (.A(_0238_),
    .B(_0221_),
    .C(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__nor2_1 _4356_ (.A(_0237_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand3_2 _4357_ (.A(_0226_),
    .B(_0241_),
    .C(_0192_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2_1 _4358_ (.A(_0235_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_1 _4359_ (.A(_0229_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__nand2_1 _4360_ (.A(_0226_),
    .B(_0192_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand2_2 _4361_ (.A(_0245_),
    .B(_0224_),
    .Y(_0246_));
 sky130_fd_sc_hd__nor2_1 _4362_ (.A(net168),
    .B(_0138_),
    .Y(_0247_));
 sky130_fd_sc_hd__nand2_1 _4363_ (.A(_0209_),
    .B(_2732_),
    .Y(_0248_));
 sky130_fd_sc_hd__mux2_1 _4364_ (.A0(net181),
    .A1(net164),
    .S(_0684_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _4365_ (.A(_0249_),
    .B(_0761_),
    .Y(_0250_));
 sky130_fd_sc_hd__o21ai_1 _4366_ (.A1(_0761_),
    .A2(net165),
    .B1(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__or2_1 _4367_ (.A(_0860_),
    .B(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__o21ai_1 _4368_ (.A1(_0849_),
    .A2(net166),
    .B1(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_1 _4369_ (.A(_0253_),
    .B(_0122_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _4370_ (.A(_0248_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__or2_1 _4371_ (.A(_0255_),
    .B(_0137_),
    .X(_0256_));
 sky130_fd_sc_hd__nor2b_1 _4372_ (.A(_0247_),
    .B_N(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__nand3_2 _4373_ (.A(_0214_),
    .B(_0257_),
    .C(_0215_),
    .Y(_0258_));
 sky130_fd_sc_hd__buf_4 _4374_ (.A(_0258_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _4375_ (.A(_0238_),
    .B(_0183_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand3_1 _4376_ (.A(_0187_),
    .B(_0185_),
    .C(_0220_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_1 _4377_ (.A(_0260_),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__nand2_1 _4378_ (.A(_0239_),
    .B(_0221_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _4379_ (.A(_0263_),
    .B(_0237_),
    .Y(_0264_));
 sky130_fd_sc_hd__nand3_1 _4380_ (.A(_0262_),
    .B(_0217_),
    .C(_0264_),
    .Y(_0265_));
 sky130_fd_sc_hd__nor2_1 _4381_ (.A(_0259_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand3_4 _4382_ (.A(_0246_),
    .B(_0242_),
    .C(_0266_),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_2 _4383_ (.A(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2_1 _4384_ (.A(_0244_),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__nand3_1 _4385_ (.A(_0229_),
    .B(_0267_),
    .C(_0243_),
    .Y(_0270_));
 sky130_fd_sc_hd__nand2_1 _4386_ (.A(_0246_),
    .B(_0242_),
    .Y(_0271_));
 sky130_fd_sc_hd__nand3_1 _4387_ (.A(_0260_),
    .B(_0261_),
    .C(_0217_),
    .Y(_0272_));
 sky130_fd_sc_hd__clkinv_4 _4388_ (.A(net169),
    .Y(_0273_));
 sky130_fd_sc_hd__o21ai_2 _4389_ (.A1(_0139_),
    .A2(net168),
    .B1(_0256_),
    .Y(_0274_));
 sky130_fd_sc_hd__nand3_1 _4390_ (.A(_0212_),
    .B(net175),
    .C(_0213_),
    .Y(_0275_));
 sky130_fd_sc_hd__o21ai_2 _4391_ (.A1(net175),
    .A2(_0274_),
    .B1(net176),
    .Y(_0276_));
 sky130_fd_sc_hd__nand3_2 _4392_ (.A(_0263_),
    .B(_0273_),
    .C(_0276_),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_2 _4393_ (.A(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand3_2 _4394_ (.A(_0272_),
    .B(_0224_),
    .C(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand2_1 _4395_ (.A(_0271_),
    .B(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_2 _4396_ (.A(_0272_),
    .B(_0224_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand2_1 _4397_ (.A(_0281_),
    .B(_0277_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand3_1 _4398_ (.A(_0239_),
    .B(_0221_),
    .C(_0237_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand3_1 _4399_ (.A(_0186_),
    .B(_0214_),
    .C(_0216_),
    .Y(_0284_));
 sky130_fd_sc_hd__nand3_1 _4400_ (.A(_0283_),
    .B(_0259_),
    .C(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_2 _4401_ (.A(\M000[18] ),
    .Y(_0286_));
 sky130_fd_sc_hd__nand2_1 _4402_ (.A(_0083_),
    .B(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__o21a_1 _4403_ (.A1(_0083_),
    .A2(net181),
    .B1(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _4404_ (.A0(_0249_),
    .A1(net182),
    .S(_0761_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _4405_ (.A(_2725_),
    .B(_0251_),
    .X(_0290_));
 sky130_fd_sc_hd__o21a_1 _4406_ (.A1(_0860_),
    .A2(_0289_),
    .B1(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_1 _4407_ (.A(_0253_),
    .B(_2732_),
    .Y(_0292_));
 sky130_fd_sc_hd__o21ai_1 _4408_ (.A1(_2732_),
    .A2(_0291_),
    .B1(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _4409_ (.A(_0293_),
    .B(_0139_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _4410_ (.A(_0137_),
    .B(_0255_),
    .Y(_0295_));
 sky130_fd_sc_hd__a21o_1 _4411_ (.A1(_0294_),
    .A2(_0295_),
    .B1(_0182_),
    .X(_0296_));
 sky130_fd_sc_hd__o21ai_2 _4412_ (.A1(_0215_),
    .A2(_0274_),
    .B1(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__nand3_1 _4413_ (.A(_0297_),
    .B(_0276_),
    .C(_0273_),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_2 _4414_ (.A(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__buf_6 _4415_ (.A(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__nand3_1 _4416_ (.A(_0285_),
    .B(_0300_),
    .C(_0277_),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_2 _4417_ (.A(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand3_1 _4418_ (.A(_0282_),
    .B(_0302_),
    .C(_0279_),
    .Y(_0303_));
 sky130_fd_sc_hd__inv_2 _4419_ (.A(_0303_),
    .Y(_0304_));
 sky130_fd_sc_hd__nand3_4 _4420_ (.A(_0280_),
    .B(_0267_),
    .C(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__a21oi_1 _4421_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _4422_ (.A(_0279_),
    .Y(_0307_));
 sky130_fd_sc_hd__nand3_1 _4423_ (.A(_0246_),
    .B(_0242_),
    .C(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__nor2_1 _4424_ (.A(_0308_),
    .B(_0244_),
    .Y(_0309_));
 sky130_fd_sc_hd__nor2_1 _4425_ (.A(_0227_),
    .B(_0235_),
    .Y(_0310_));
 sky130_fd_sc_hd__nor2_1 _4426_ (.A(_0149_),
    .B(_0169_),
    .Y(_0311_));
 sky130_fd_sc_hd__nand2_1 _4427_ (.A(_0163_),
    .B(_0151_),
    .Y(_0312_));
 sky130_fd_sc_hd__nand2_1 _4428_ (.A(_1674_),
    .B(net20),
    .Y(_0313_));
 sky130_fd_sc_hd__o21ai_4 _4429_ (.A1(_1355_),
    .A2(_1663_),
    .B1(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__nand2_1 _4430_ (.A(_0159_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_2 _4431_ (.A(_0314_),
    .Y(_0316_));
 sky130_fd_sc_hd__nand2_1 _4432_ (.A(_0162_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _4433_ (.A(_0315_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__nand2_1 _4434_ (.A(_0312_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__nor2_1 _4435_ (.A(_0105_),
    .B(_0160_),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_2 _4436_ (.A(_0318_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_1 _4437_ (.A(_0320_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__nand2_1 _4438_ (.A(_0319_),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_2 _4439_ (.A(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_2 _4440_ (.A(_0168_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(_0324_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_1 _4442_ (.A(_0323_),
    .B(_0168_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand3_2 _4443_ (.A(_0311_),
    .B(_0326_),
    .C(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_2 _4444_ (.A(_0149_),
    .Y(_0329_));
 sky130_fd_sc_hd__nand2_1 _4445_ (.A(_0171_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _4446_ (.A(_0326_),
    .B(_0327_),
    .Y(_0331_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(_0330_),
    .B(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__nand2_1 _4448_ (.A(_0328_),
    .B(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__nor2_2 _4449_ (.A(_0169_),
    .B(_0191_),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_2 _4450_ (.A(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _4451_ (.A(_0333_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand3_4 _4452_ (.A(_0328_),
    .B(_0332_),
    .C(_0334_),
    .Y(_0337_));
 sky130_fd_sc_hd__nand2_1 _4453_ (.A(_0336_),
    .B(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _4454_ (.A(_0338_),
    .B(_0234_),
    .Y(_0339_));
 sky130_fd_sc_hd__a21oi_1 _4455_ (.A1(_0170_),
    .A2(_0172_),
    .B1(_0231_),
    .Y(_0340_));
 sky130_fd_sc_hd__nand3_2 _4456_ (.A(_0340_),
    .B(_0336_),
    .C(_0337_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand3_2 _4457_ (.A(_0310_),
    .B(_0339_),
    .C(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _4458_ (.A(_0339_),
    .B(_0341_),
    .Y(_0343_));
 sky130_fd_sc_hd__nand2_1 _4459_ (.A(_0343_),
    .B(_0229_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand3_2 _4460_ (.A(_0309_),
    .B(_0342_),
    .C(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nand2_1 _4461_ (.A(_0344_),
    .B(_0342_),
    .Y(_0346_));
 sky130_fd_sc_hd__nand3b_1 _4462_ (.A_N(_0308_),
    .B(_0229_),
    .C(_0243_),
    .Y(_0347_));
 sky130_fd_sc_hd__nand2_1 _4463_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand3_2 _4464_ (.A(_0306_),
    .B(_0345_),
    .C(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _4465_ (.A(_0345_),
    .B(_0348_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _4466_ (.A(_0269_),
    .B(_0270_),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_2 _4467_ (.A(_0305_),
    .Y(_0352_));
 sky130_fd_sc_hd__nand2_2 _4468_ (.A(_0351_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _4469_ (.A(_0350_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _4470_ (.A(_0349_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__nand2_1 _4471_ (.A(_0280_),
    .B(_0267_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_1 _4472_ (.A(_0356_),
    .B(_0303_),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_2 _4473_ (.A(_0285_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _4474_ (.A(_0297_),
    .B(_0273_),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_1 _4475_ (.A(_0276_),
    .B(net169),
    .Y(_0360_));
 sky130_fd_sc_hd__nand2_1 _4476_ (.A(_0359_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _4477_ (.A(_0361_),
    .B(_0258_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2_1 _4478_ (.A(_0297_),
    .B(net169),
    .Y(_0363_));
 sky130_fd_sc_hd__a21o_1 _4479_ (.A1(_0294_),
    .A2(_0295_),
    .B1(_0215_),
    .X(_0364_));
 sky130_fd_sc_hd__or2_1 _4480_ (.A(_0123_),
    .B(_0291_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_0083_),
    .B(\M000[18] ),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_0695_),
    .B(net181),
    .Y(_0367_));
 sky130_fd_sc_hd__nand2_1 _4483_ (.A(_0286_),
    .B(_0684_),
    .Y(_0368_));
 sky130_fd_sc_hd__o21a_1 _4484_ (.A1(_0684_),
    .A2(\M000[17] ),
    .B1(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__nor2_1 _4485_ (.A(_2719_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a31o_1 _4486_ (.A1(_2719_),
    .A2(_0366_),
    .A3(_0367_),
    .B1(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _4487_ (.A(_0371_),
    .B(_2725_),
    .Y(_0372_));
 sky130_fd_sc_hd__o21a_1 _4488_ (.A1(_2725_),
    .A2(_0289_),
    .B1(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _4489_ (.A(_2732_),
    .B(_0373_),
    .X(_0374_));
 sky130_fd_sc_hd__nand3_1 _4490_ (.A(_0365_),
    .B(_0139_),
    .C(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__o211ai_2 _4491_ (.A1(_2732_),
    .A2(_0291_),
    .B1(_0292_),
    .C1(_0137_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand3_1 _4492_ (.A(_0375_),
    .B(_0376_),
    .C(_0215_),
    .Y(_0377_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(_0364_),
    .B(net183),
    .Y(_0378_));
 sky130_fd_sc_hd__nand2_1 _4494_ (.A(_0378_),
    .B(_0273_),
    .Y(_0379_));
 sky130_fd_sc_hd__nand2_1 _4495_ (.A(_0363_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_2 _4496_ (.A(_0258_),
    .Y(_0381_));
 sky130_fd_sc_hd__buf_4 _4497_ (.A(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _4498_ (.A(_0380_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__nand2_2 _4499_ (.A(_0362_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__o2111ai_4 _4500_ (.A1(_0278_),
    .A2(_0358_),
    .B1(_0281_),
    .C1(_0300_),
    .D1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__inv_2 _4501_ (.A(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__nand3_4 _4502_ (.A(_0357_),
    .B(_0305_),
    .C(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__inv_2 _4503_ (.A(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__nand3_1 _4504_ (.A(_0269_),
    .B(_0305_),
    .C(_0270_),
    .Y(_0389_));
 sky130_fd_sc_hd__nand3_1 _4505_ (.A(_0388_),
    .B(_0353_),
    .C(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__nand2_1 _4506_ (.A(_0355_),
    .B(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(_0353_),
    .B(_0389_),
    .Y(_0392_));
 sky130_fd_sc_hd__nor2_1 _4508_ (.A(_0387_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__nand3_2 _4509_ (.A(_0393_),
    .B(_0349_),
    .C(_0354_),
    .Y(_0394_));
 sky130_fd_sc_hd__nand2_1 _4510_ (.A(_0391_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_0392_),
    .B(_0388_),
    .Y(_0396_));
 sky130_fd_sc_hd__nand3_1 _4512_ (.A(_0353_),
    .B(_0387_),
    .C(_0389_),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _4513_ (.A(_0396_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_1 _4514_ (.A(_0357_),
    .B(_0305_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _4515_ (.A(_0399_),
    .B(_0385_),
    .Y(_0400_));
 sky130_fd_sc_hd__buf_2 _4516_ (.A(net177),
    .X(_0401_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_0285_),
    .B(_0277_),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_2 _4518_ (.A(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__o21ai_1 _4519_ (.A1(_0401_),
    .A2(_0384_),
    .B1(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__nand3_1 _4520_ (.A(_0361_),
    .B(_0380_),
    .C(_0382_),
    .Y(_0405_));
 sky130_fd_sc_hd__buf_4 _4521_ (.A(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__nand3_1 _4522_ (.A(_0406_),
    .B(_0402_),
    .C(_0300_),
    .Y(_0407_));
 sky130_fd_sc_hd__nand2_1 _4523_ (.A(_0404_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nand2_1 _4524_ (.A(_0380_),
    .B(_0258_),
    .Y(_0409_));
 sky130_fd_sc_hd__nand3_1 _4525_ (.A(_0364_),
    .B(_0236_),
    .C(_0377_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand3_1 _4526_ (.A(_0375_),
    .B(_0376_),
    .C(_0182_),
    .Y(_0411_));
 sky130_fd_sc_hd__nand3_1 _4527_ (.A(_0365_),
    .B(_0374_),
    .C(_0137_),
    .Y(_0412_));
 sky130_fd_sc_hd__nand2_1 _4528_ (.A(_0373_),
    .B(_2732_),
    .Y(_0413_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(\M000[16] ),
    .A1(\M000[17] ),
    .S(_0695_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(_0414_),
    .A1(_0369_),
    .S(_2719_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_1 _4531_ (.A(_0415_),
    .B(_2725_),
    .Y(_0416_));
 sky130_fd_sc_hd__o21ai_1 _4532_ (.A1(_2725_),
    .A2(_0371_),
    .B1(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__nand2_1 _4533_ (.A(_0417_),
    .B(_0123_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_0413_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _4535_ (.A(_0139_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand3_1 _4536_ (.A(_0412_),
    .B(_0215_),
    .C(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__nand3_1 _4537_ (.A(_0411_),
    .B(_0421_),
    .C(_0273_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand3_1 _4538_ (.A(_0381_),
    .B(_0410_),
    .C(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__nand2_1 _4539_ (.A(_0409_),
    .B(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand3_4 _4540_ (.A(_0384_),
    .B(_0424_),
    .C(_0299_),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_4 _4541_ (.A(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__buf_6 _4542_ (.A(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _4543_ (.A(_0408_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__clkbuf_4 _4544_ (.A(_0300_),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_1 _4545_ (.A(_0281_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand3_1 _4546_ (.A(_0282_),
    .B(_0279_),
    .C(_0401_),
    .Y(_0431_));
 sky130_fd_sc_hd__o211ai_2 _4547_ (.A1(_0403_),
    .A2(_0406_),
    .B1(_0430_),
    .C1(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__nand3b_2 _4548_ (.A_N(_0428_),
    .B(_0432_),
    .C(_0385_),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_2 _4549_ (.A(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__nand3_2 _4550_ (.A(_0400_),
    .B(_0434_),
    .C(_0387_),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_2 _4551_ (.A(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(_0398_),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__nand2_1 _4553_ (.A(_0395_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nand2_1 _4554_ (.A(_0392_),
    .B(_0387_),
    .Y(_0439_));
 sky130_fd_sc_hd__nand2_1 _4555_ (.A(_0390_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _4556_ (.A(_0435_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand3_2 _4557_ (.A(_0441_),
    .B(_0391_),
    .C(_0394_),
    .Y(_0442_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_0438_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _4559_ (.A(_0400_),
    .B(_0387_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _4560_ (.A(_0444_),
    .B(_0433_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_0445_),
    .B(_0435_),
    .Y(_0446_));
 sky130_fd_sc_hd__inv_2 _4562_ (.A(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_1 _4563_ (.A(_0432_),
    .B(_0385_),
    .Y(_0448_));
 sky130_fd_sc_hd__nand2_1 _4564_ (.A(_0448_),
    .B(_0428_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _4565_ (.A(_0408_),
    .B(_0425_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand3_1 _4566_ (.A(_0427_),
    .B(_0404_),
    .C(_0407_),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_1 _4567_ (.A(_0450_),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__a21o_1 _4568_ (.A1(_0424_),
    .A2(_0299_),
    .B1(_0384_),
    .X(_0453_));
 sky130_fd_sc_hd__nand3_1 _4569_ (.A(_0409_),
    .B(_0401_),
    .C(_0423_),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_2 _4570_ (.A(\M000[15] ),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _4571_ (.A(_0083_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__o21a_1 _4572_ (.A1(_0083_),
    .A2(\M000[16] ),
    .B1(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _4573_ (.A0(_0414_),
    .A1(_0457_),
    .S(_0761_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _4574_ (.A0(_0458_),
    .A1(_0415_),
    .S(_0871_),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_1 _4575_ (.A(_0459_),
    .B(_0123_),
    .Y(_0460_));
 sky130_fd_sc_hd__nand2_1 _4576_ (.A(_0417_),
    .B(_2732_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2_1 _4577_ (.A(_0460_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_1 _4578_ (.A(_0462_),
    .B(_0139_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_1 _4579_ (.A(_0419_),
    .B(_0137_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand2_1 _4580_ (.A(_0463_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__or2_1 _4581_ (.A(_0183_),
    .B(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__nand3_1 _4582_ (.A(_0412_),
    .B(_0183_),
    .C(_0420_),
    .Y(_0467_));
 sky130_fd_sc_hd__nand3_1 _4583_ (.A(_0466_),
    .B(_0273_),
    .C(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__nand3_1 _4584_ (.A(_0411_),
    .B(_0421_),
    .C(_0236_),
    .Y(_0469_));
 sky130_fd_sc_hd__nand3_1 _4585_ (.A(_0468_),
    .B(_0382_),
    .C(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand3_1 _4586_ (.A(_0410_),
    .B(_0258_),
    .C(_0422_),
    .Y(_0471_));
 sky130_fd_sc_hd__nand3_1 _4587_ (.A(_0299_),
    .B(_0470_),
    .C(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _4588_ (.A(_0454_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_2 _4589_ (.A(_0405_),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_1 _4590_ (.A(_0473_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand3_4 _4591_ (.A(_0453_),
    .B(_0475_),
    .C(_0426_),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_6 _4592_ (.A(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_0452_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_2 _4594_ (.A(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand3_1 _4595_ (.A(_0449_),
    .B(_0433_),
    .C(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_2 _4596_ (.A(_0480_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand2_1 _4597_ (.A(_0447_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nand3_1 _4598_ (.A(_0396_),
    .B(_0435_),
    .C(_0397_),
    .Y(_0483_));
 sky130_fd_sc_hd__nand2_1 _4599_ (.A(_0437_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__nor2_1 _4600_ (.A(_0482_),
    .B(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_2 _4601_ (.A(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__nand2_1 _4602_ (.A(_0443_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__nand3_2 _4603_ (.A(_0485_),
    .B(_0438_),
    .C(_0442_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_1 _4604_ (.A(_0487_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2_1 _4605_ (.A(_0446_),
    .B(_0480_),
    .Y(_0490_));
 sky130_fd_sc_hd__clkbuf_4 _4606_ (.A(_0476_),
    .X(_0491_));
 sky130_fd_sc_hd__inv_2 _4607_ (.A(_0448_),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_2 _4608_ (.A(_0408_),
    .Y(_0493_));
 sky130_fd_sc_hd__clkbuf_4 _4609_ (.A(_0425_),
    .X(_0494_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(_0493_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__nand3_1 _4611_ (.A(_0492_),
    .B(_0428_),
    .C(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__nor2_1 _4612_ (.A(_0491_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand3_2 _4613_ (.A(_0445_),
    .B(_0497_),
    .C(_0435_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2_1 _4614_ (.A(_0449_),
    .B(_0433_),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_2 _4615_ (.A(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _4616_ (.A(_0453_),
    .B(_0475_),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_2 _4617_ (.A(_0501_),
    .Y(_0502_));
 sky130_fd_sc_hd__nand2_1 _4618_ (.A(_0502_),
    .B(_0425_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand3_1 _4619_ (.A(_0466_),
    .B(_0236_),
    .C(_0467_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_1 _4620_ (.A(_0459_),
    .B(_2733_),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_2 _4621_ (.A(\M000[14] ),
    .Y(_0506_));
 sky130_fd_sc_hd__mux2_1 _4622_ (.A0(_0506_),
    .A1(_0455_),
    .S(_0695_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _4623_ (.A(_0507_),
    .B(_0761_),
    .Y(_0508_));
 sky130_fd_sc_hd__o21a_1 _4624_ (.A1(_0772_),
    .A2(_0457_),
    .B1(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _4625_ (.A0(_0458_),
    .A1(_0509_),
    .S(_2725_),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _4626_ (.A(_0510_),
    .B(_0123_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _4627_ (.A(_0505_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__nand2_1 _4628_ (.A(_0512_),
    .B(_0139_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(_0462_),
    .B(_0137_),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_1 _4630_ (.A(_0513_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _4631_ (.A(_0515_),
    .B(_0215_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _4632_ (.A(_0465_),
    .B(_0183_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_1 _4633_ (.A(_0516_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _4634_ (.A(_0518_),
    .B(_0273_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand3_1 _4635_ (.A(_0504_),
    .B(_0382_),
    .C(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand3_1 _4636_ (.A(_0468_),
    .B(_0469_),
    .C(_0259_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand3_1 _4637_ (.A(_0299_),
    .B(_0520_),
    .C(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand3_1 _4638_ (.A(_0470_),
    .B(_0471_),
    .C(_0401_),
    .Y(_0523_));
 sky130_fd_sc_hd__nand2_1 _4639_ (.A(_0522_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__nand3_1 _4640_ (.A(_0454_),
    .B(_0406_),
    .C(_0472_),
    .Y(_0525_));
 sky130_fd_sc_hd__o21ai_2 _4641_ (.A1(_0406_),
    .A2(_0524_),
    .B1(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_1 _4642_ (.A(_0526_),
    .B(_0426_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_2 _4643_ (.A(_0503_),
    .B(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__inv_2 _4644_ (.A(_0452_),
    .Y(_0529_));
 sky130_fd_sc_hd__nand3_1 _4645_ (.A(_0528_),
    .B(_0529_),
    .C(_0477_),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _4646_ (.A(_0530_),
    .Y(_0531_));
 sky130_fd_sc_hd__nand2_1 _4647_ (.A(_0500_),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_2 _4648_ (.A(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__nand3_2 _4649_ (.A(_0490_),
    .B(_0498_),
    .C(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__nor2_1 _4650_ (.A(_0484_),
    .B(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__inv_2 _4651_ (.A(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__nand2_1 _4652_ (.A(_0489_),
    .B(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand3_2 _4653_ (.A(_0487_),
    .B(_0488_),
    .C(_0535_),
    .Y(_0538_));
 sky130_fd_sc_hd__nand2_1 _4654_ (.A(_0537_),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__nand2_1 _4655_ (.A(_0490_),
    .B(_0498_),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(_0540_),
    .B(_0532_),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _4657_ (.A(_0499_),
    .B(_0478_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand3_2 _4658_ (.A(_0502_),
    .B(_0526_),
    .C(_0427_),
    .Y(_0543_));
 sky130_fd_sc_hd__clkbuf_4 _4659_ (.A(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__nand3_1 _4660_ (.A(_0542_),
    .B(_0480_),
    .C(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__clkinv_4 _4661_ (.A(_0543_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _4662_ (.A(_0499_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _4663_ (.A(_0545_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__a21o_1 _4664_ (.A1(_0520_),
    .A2(_0521_),
    .B1(_0300_),
    .X(_0549_));
 sky130_fd_sc_hd__a21o_1 _4665_ (.A1(_0504_),
    .A2(_0519_),
    .B1(_0382_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _4666_ (.A0(\M000[13] ),
    .A1(\M000[14] ),
    .S(_0695_),
    .X(_0551_));
 sky130_fd_sc_hd__nand2_1 _4667_ (.A(_0507_),
    .B(_2719_),
    .Y(_0552_));
 sky130_fd_sc_hd__o21a_1 _4668_ (.A1(_2719_),
    .A2(_0551_),
    .B1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__inv_2 _4669_ (.A(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__nand2_1 _4670_ (.A(_0554_),
    .B(_2725_),
    .Y(_0555_));
 sky130_fd_sc_hd__o21ai_1 _4671_ (.A1(_2726_),
    .A2(_0509_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nand2_1 _4672_ (.A(_0510_),
    .B(_2733_),
    .Y(_0557_));
 sky130_fd_sc_hd__o21ai_1 _4673_ (.A1(_2733_),
    .A2(_0556_),
    .B1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_0558_),
    .B(_0139_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _4675_ (.A(_0512_),
    .B(_0198_),
    .Y(_0560_));
 sky130_fd_sc_hd__nand2_1 _4676_ (.A(_0559_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _4677_ (.A(_0561_),
    .B(_0216_),
    .Y(_0562_));
 sky130_fd_sc_hd__nand2_1 _4678_ (.A(_0515_),
    .B(_0183_),
    .Y(_0563_));
 sky130_fd_sc_hd__nand2_1 _4679_ (.A(_0562_),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _4680_ (.A(_0564_),
    .B(_0273_),
    .Y(_0565_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_0518_),
    .B(_0237_),
    .Y(_0566_));
 sky130_fd_sc_hd__nand2_1 _4682_ (.A(_0565_),
    .B(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__nand2_1 _4683_ (.A(_0567_),
    .B(_0382_),
    .Y(_0568_));
 sky130_fd_sc_hd__nand3_1 _4684_ (.A(_0550_),
    .B(_0300_),
    .C(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__nand3_1 _4685_ (.A(_0549_),
    .B(_0569_),
    .C(_0474_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(_0524_),
    .B(_0406_),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_0570_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(_0526_),
    .B(_0425_),
    .Y(_0573_));
 sky130_fd_sc_hd__o21ai_4 _4689_ (.A1(_0425_),
    .A2(_0572_),
    .B1(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__nand2_1 _4690_ (.A(_0574_),
    .B(_0477_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _4691_ (.A(_0528_),
    .B(_0476_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _4692_ (.A(_0575_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nand2_1 _4693_ (.A(_0529_),
    .B(_0476_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand2_1 _4694_ (.A(_0578_),
    .B(_0478_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand3_2 _4695_ (.A(_0577_),
    .B(_0546_),
    .C(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__inv_2 _4696_ (.A(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nand2_1 _4697_ (.A(_0548_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_2 _4698_ (.A(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_2 _4699_ (.A(_0541_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__inv_2 _4700_ (.A(_0498_),
    .Y(_0585_));
 sky130_fd_sc_hd__nand2_1 _4701_ (.A(_0484_),
    .B(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand3_1 _4702_ (.A(_0437_),
    .B(_0498_),
    .C(_0483_),
    .Y(_0587_));
 sky130_fd_sc_hd__nand2_1 _4703_ (.A(_0586_),
    .B(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_2 _4704_ (.A(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2_1 _4705_ (.A(_0584_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_2 _4706_ (.A(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_0539_),
    .B(_0591_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand3_4 _4708_ (.A(_0537_),
    .B(_0538_),
    .C(_0590_),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _4709_ (.A(_0592_),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _4710_ (.A(_0541_),
    .B(_0534_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_1 _4711_ (.A(_0595_),
    .B(_0582_),
    .Y(_0596_));
 sky130_fd_sc_hd__nand2_1 _4712_ (.A(_0579_),
    .B(_0544_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _4713_ (.A(_0597_),
    .B(_0530_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand3_4 _4714_ (.A(_0574_),
    .B(_0528_),
    .C(_0477_),
    .Y(_0599_));
 sky130_fd_sc_hd__nand2_1 _4715_ (.A(_0598_),
    .B(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_2 _4716_ (.A(_0600_),
    .B(_0580_),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_2 _4717_ (.A(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _4718_ (.A(_0574_),
    .B(_0476_),
    .Y(_0603_));
 sky130_fd_sc_hd__nand2_1 _4719_ (.A(_0572_),
    .B(_0425_),
    .Y(_0604_));
 sky130_fd_sc_hd__or2_1 _4720_ (.A(_0259_),
    .B(_0567_),
    .X(_0605_));
 sky130_fd_sc_hd__nand3_1 _4721_ (.A(_0504_),
    .B(_0259_),
    .C(_0519_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand3_1 _4722_ (.A(_0605_),
    .B(_0401_),
    .C(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(_0558_),
    .B(_0198_),
    .Y(_0608_));
 sky130_fd_sc_hd__clkbuf_4 _4724_ (.A(_0123_),
    .X(_0609_));
 sky130_fd_sc_hd__inv_2 _4725_ (.A(\M000[12] ),
    .Y(_0610_));
 sky130_fd_sc_hd__nand2_1 _4726_ (.A(_0083_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__o21a_1 _4727_ (.A1(_0083_),
    .A2(\M000[13] ),
    .B1(_0611_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _4728_ (.A0(_0551_),
    .A1(_0612_),
    .S(_0772_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _4729_ (.A0(_0613_),
    .A1(_0553_),
    .S(_0871_),
    .X(_0614_));
 sky130_fd_sc_hd__nand2_1 _4730_ (.A(_0614_),
    .B(_0123_),
    .Y(_0615_));
 sky130_fd_sc_hd__o21ai_1 _4731_ (.A1(_0609_),
    .A2(_0556_),
    .B1(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _4732_ (.A(_0616_),
    .B(_0185_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_0608_),
    .B(_0617_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(_0618_),
    .B(_0216_),
    .Y(_0619_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_0561_),
    .B(_0183_),
    .Y(_0620_));
 sky130_fd_sc_hd__nand2_1 _4736_ (.A(_0619_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__nand2_1 _4737_ (.A(_0621_),
    .B(_0273_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0564_),
    .B(_0237_),
    .Y(_0623_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(_0622_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _4740_ (.A(_0624_),
    .B(_0382_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _4741_ (.A(_0567_),
    .B(_0259_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _4742_ (.A(_0625_),
    .B(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _4743_ (.A(_0627_),
    .B(_0300_),
    .Y(_0628_));
 sky130_fd_sc_hd__nand3_1 _4744_ (.A(_0607_),
    .B(_0474_),
    .C(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__nand3_1 _4745_ (.A(_0605_),
    .B(_0300_),
    .C(_0606_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand3_1 _4746_ (.A(_0520_),
    .B(_0521_),
    .C(_0401_),
    .Y(_0631_));
 sky130_fd_sc_hd__nand3_1 _4747_ (.A(_0630_),
    .B(_0406_),
    .C(_0631_),
    .Y(_0632_));
 sky130_fd_sc_hd__nand3_1 _4748_ (.A(_0629_),
    .B(_0632_),
    .C(_0427_),
    .Y(_0633_));
 sky130_fd_sc_hd__nand3_1 _4749_ (.A(_0604_),
    .B(_0477_),
    .C(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _4750_ (.A(_0603_),
    .B(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__nand3_2 _4751_ (.A(_0577_),
    .B(_0635_),
    .C(_0546_),
    .Y(_0636_));
 sky130_fd_sc_hd__inv_4 _4752_ (.A(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__buf_6 _4753_ (.A(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__nand3_2 _4754_ (.A(_0602_),
    .B(_0548_),
    .C(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__inv_2 _4755_ (.A(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nand3_2 _4756_ (.A(_0596_),
    .B(_0584_),
    .C(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__inv_2 _4757_ (.A(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand2_1 _4758_ (.A(_0584_),
    .B(_0534_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(_0643_),
    .B(_0589_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand3_1 _4760_ (.A(_0584_),
    .B(_0588_),
    .C(_0534_),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _4761_ (.A(_0644_),
    .B(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_2 _4762_ (.A(_0642_),
    .B(_0646_),
    .Y(_0647_));
 sky130_fd_sc_hd__nand2_1 _4763_ (.A(_0594_),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__inv_2 _4764_ (.A(_0647_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand3_2 _4765_ (.A(_0592_),
    .B(_0649_),
    .C(_0593_),
    .Y(_0650_));
 sky130_fd_sc_hd__nand2_1 _4766_ (.A(_0648_),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__nand2_1 _4767_ (.A(_0596_),
    .B(_0584_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_0652_),
    .B(_0639_),
    .Y(_0653_));
 sky130_fd_sc_hd__nand3_1 _4769_ (.A(_0545_),
    .B(_0580_),
    .C(_0547_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_1 _4770_ (.A(_0582_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(_0602_),
    .B(_0638_),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _4772_ (.A(_0655_),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__a21o_1 _4773_ (.A1(_0574_),
    .A2(_0477_),
    .B1(_0528_),
    .X(_0658_));
 sky130_fd_sc_hd__nand3_1 _4774_ (.A(_0603_),
    .B(_0546_),
    .C(_0634_),
    .Y(_0659_));
 sky130_fd_sc_hd__nand3_1 _4775_ (.A(_0658_),
    .B(_0659_),
    .C(_0599_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand3_1 _4776_ (.A(_0603_),
    .B(_0543_),
    .C(_0634_),
    .Y(_0661_));
 sky130_fd_sc_hd__inv_2 _4777_ (.A(_0599_),
    .Y(_0662_));
 sky130_fd_sc_hd__nand3_1 _4778_ (.A(_0604_),
    .B(_0633_),
    .C(_0476_),
    .Y(_0663_));
 sky130_fd_sc_hd__inv_2 _4779_ (.A(\M000[11] ),
    .Y(_0664_));
 sky130_fd_sc_hd__mux2_1 _4780_ (.A0(_0664_),
    .A1(_0610_),
    .S(_0695_),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_0665_),
    .B(_0772_),
    .Y(_0666_));
 sky130_fd_sc_hd__o21a_1 _4782_ (.A1(_0772_),
    .A2(_0612_),
    .B1(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_1 _4783_ (.A0(_0613_),
    .A1(_0667_),
    .S(_2725_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _4784_ (.A0(_0668_),
    .A1(_0614_),
    .S(_2733_),
    .X(_0669_));
 sky130_fd_sc_hd__nand2_1 _4785_ (.A(_0669_),
    .B(_0185_),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _4786_ (.A(_0616_),
    .B(_0198_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _4787_ (.A(_0670_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__nand2_1 _4788_ (.A(_0672_),
    .B(_0216_),
    .Y(_0673_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_0618_),
    .B(_0183_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _4790_ (.A(_0673_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__buf_2 _4791_ (.A(_0273_),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_1 _4792_ (.A(_0675_),
    .B(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_0621_),
    .B(_0237_),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _4794_ (.A(_0677_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__nand2_1 _4795_ (.A(_0679_),
    .B(_0382_),
    .Y(_0680_));
 sky130_fd_sc_hd__nand2_1 _4796_ (.A(_0624_),
    .B(_0259_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _4797_ (.A(_0680_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _4798_ (.A(_0682_),
    .B(_0300_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _4799_ (.A(_0627_),
    .B(_0401_),
    .Y(_0685_));
 sky130_fd_sc_hd__nand3_1 _4800_ (.A(_0683_),
    .B(_0685_),
    .C(_0474_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand3_1 _4801_ (.A(_0607_),
    .B(_0406_),
    .C(_0628_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand3_1 _4802_ (.A(_0686_),
    .B(_0427_),
    .C(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand3_1 _4803_ (.A(_0629_),
    .B(_0632_),
    .C(_0425_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand3_1 _4804_ (.A(_0477_),
    .B(_0688_),
    .C(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__nand3_1 _4805_ (.A(_0663_),
    .B(_0690_),
    .C(_0546_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand3_1 _4806_ (.A(_0661_),
    .B(_0662_),
    .C(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _4807_ (.A(_0660_),
    .B(_0692_),
    .Y(_0693_));
 sky130_fd_sc_hd__nand3_2 _4808_ (.A(_0693_),
    .B(_0601_),
    .C(_0638_),
    .Y(_0694_));
 sky130_fd_sc_hd__inv_2 _4809_ (.A(_0694_),
    .Y(_0696_));
 sky130_fd_sc_hd__nand3_2 _4810_ (.A(_0657_),
    .B(_0639_),
    .C(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__inv_2 _4811_ (.A(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__nand3_1 _4812_ (.A(_0653_),
    .B(_0641_),
    .C(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__inv_2 _4813_ (.A(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand3_1 _4814_ (.A(_0641_),
    .B(_0645_),
    .C(_0644_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand3_2 _4815_ (.A(_0700_),
    .B(_0647_),
    .C(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_1 _4816_ (.A(_0651_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__nand2_1 _4817_ (.A(_0701_),
    .B(_0647_),
    .Y(_0704_));
 sky130_fd_sc_hd__nor2_1 _4818_ (.A(_0699_),
    .B(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__nand3_2 _4819_ (.A(_0648_),
    .B(_0650_),
    .C(_0705_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand2_1 _4820_ (.A(_0703_),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(_0653_),
    .B(_0641_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand2_1 _4822_ (.A(_0709_),
    .B(_0697_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _4823_ (.A(_0693_),
    .B(_0637_),
    .Y(_0711_));
 sky130_fd_sc_hd__buf_6 _4824_ (.A(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_1 _4825_ (.A(_0601_),
    .B(_0638_),
    .Y(_0713_));
 sky130_fd_sc_hd__clkbuf_4 _4826_ (.A(_0636_),
    .X(_0714_));
 sky130_fd_sc_hd__nand3_1 _4827_ (.A(_0600_),
    .B(_0580_),
    .C(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand2_1 _4828_ (.A(_0713_),
    .B(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__nand3_1 _4829_ (.A(_0657_),
    .B(_0639_),
    .C(_0716_),
    .Y(_0718_));
 sky130_fd_sc_hd__nor2_1 _4830_ (.A(_0712_),
    .B(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__nand3_2 _4831_ (.A(_0653_),
    .B(_0719_),
    .C(_0641_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_0657_),
    .B(_0639_),
    .Y(_0721_));
 sky130_fd_sc_hd__a21o_1 _4833_ (.A1(_0607_),
    .A2(_0628_),
    .B1(_0474_),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_1 _4834_ (.A(_0683_),
    .B(_0685_),
    .Y(_0723_));
 sky130_fd_sc_hd__nand2_1 _4835_ (.A(_0723_),
    .B(_0474_),
    .Y(_0724_));
 sky130_fd_sc_hd__nand3_1 _4836_ (.A(_0722_),
    .B(_0425_),
    .C(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2_1 _4837_ (.A(_0669_),
    .B(_0198_),
    .Y(_0726_));
 sky130_fd_sc_hd__mux2_1 _4838_ (.A0(\M000[10] ),
    .A1(\M000[11] ),
    .S(_0695_),
    .X(_0727_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_0727_),
    .B(_0772_),
    .Y(_0729_));
 sky130_fd_sc_hd__o21ai_1 _4840_ (.A1(_0772_),
    .A2(_0665_),
    .B1(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__inv_2 _4841_ (.A(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__nand2_1 _4842_ (.A(_0731_),
    .B(_2726_),
    .Y(_0732_));
 sky130_fd_sc_hd__o21a_1 _4843_ (.A1(_2726_),
    .A2(_0667_),
    .B1(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(_0668_),
    .A1(_0733_),
    .S(_0123_),
    .X(_0734_));
 sky130_fd_sc_hd__nand2_1 _4845_ (.A(_0734_),
    .B(_0185_),
    .Y(_0735_));
 sky130_fd_sc_hd__nand2_1 _4846_ (.A(_0726_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _4847_ (.A(_0736_),
    .B(_0216_),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _4848_ (.A(_0672_),
    .B(_0183_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand2_1 _4849_ (.A(_0737_),
    .B(_0738_),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(_0740_),
    .B(_0676_),
    .Y(_0741_));
 sky130_fd_sc_hd__nand2_1 _4851_ (.A(_0675_),
    .B(_0237_),
    .Y(_0742_));
 sky130_fd_sc_hd__nand2_1 _4852_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__nand2_1 _4853_ (.A(_0743_),
    .B(_0382_),
    .Y(_0744_));
 sky130_fd_sc_hd__nand2_1 _4854_ (.A(_0679_),
    .B(_0259_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_0744_),
    .B(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_1 _4856_ (.A(_0746_),
    .B(_0300_),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(_0682_),
    .B(_0401_),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _4858_ (.A(_0747_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nand2_1 _4859_ (.A(_0749_),
    .B(_0474_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _4860_ (.A(_0723_),
    .B(_0406_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand3_1 _4861_ (.A(_0751_),
    .B(_0752_),
    .C(_0427_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand3_1 _4862_ (.A(_0725_),
    .B(_0753_),
    .C(_0477_),
    .Y(_0754_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(_0688_),
    .B(_0689_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _4864_ (.A(_0755_),
    .B(_0476_),
    .Y(_0756_));
 sky130_fd_sc_hd__nand3_1 _4865_ (.A(_0754_),
    .B(_0546_),
    .C(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__nand2_1 _4866_ (.A(_0690_),
    .B(_0663_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand2_1 _4867_ (.A(_0758_),
    .B(_0543_),
    .Y(_0759_));
 sky130_fd_sc_hd__nand2_1 _4868_ (.A(_0757_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _4869_ (.A(_0760_),
    .B(_0662_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand3_1 _4870_ (.A(_0661_),
    .B(_0691_),
    .C(_0599_),
    .Y(_0763_));
 sky130_fd_sc_hd__nand2_1 _4871_ (.A(_0762_),
    .B(_0763_),
    .Y(_0764_));
 sky130_fd_sc_hd__nand3_1 _4872_ (.A(_0693_),
    .B(_0764_),
    .C(_0638_),
    .Y(_0765_));
 sky130_fd_sc_hd__buf_6 _4873_ (.A(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__or2_1 _4874_ (.A(_0766_),
    .B(_0716_),
    .X(_0767_));
 sky130_fd_sc_hd__or2_2 _4875_ (.A(_0721_),
    .B(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__inv_2 _4876_ (.A(_0768_),
    .Y(_0769_));
 sky130_fd_sc_hd__nand3_4 _4877_ (.A(_0710_),
    .B(_0720_),
    .C(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__inv_2 _4878_ (.A(_0770_),
    .Y(_0771_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(_0704_),
    .B(_0720_),
    .Y(_0773_));
 sky130_fd_sc_hd__nand3_2 _4880_ (.A(_0771_),
    .B(_0702_),
    .C(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__nand2_1 _4881_ (.A(_0708_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(_0702_),
    .B(_0773_),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_1 _4883_ (.A(_0770_),
    .B(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__nand3_2 _4884_ (.A(_0777_),
    .B(_0703_),
    .C(_0707_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(_0775_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _4886_ (.A(_0710_),
    .B(_0720_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand2_1 _4887_ (.A(_0780_),
    .B(_0768_),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_1 _4888_ (.A(_0721_),
    .B(_0694_),
    .Y(_0782_));
 sky130_fd_sc_hd__nand2_1 _4889_ (.A(_0782_),
    .B(_0697_),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2_1 _4890_ (.A(_0784_),
    .B(_0767_),
    .Y(_0785_));
 sky130_fd_sc_hd__nand2_1 _4891_ (.A(_0764_),
    .B(_0714_),
    .Y(_0786_));
 sky130_fd_sc_hd__or2b_1 _4892_ (.A(_0736_),
    .B_N(_0184_),
    .X(_0787_));
 sky130_fd_sc_hd__buf_2 _4893_ (.A(_0185_),
    .X(_0788_));
 sky130_fd_sc_hd__inv_2 _4894_ (.A(\M000[9] ),
    .Y(_0789_));
 sky130_fd_sc_hd__inv_2 _4895_ (.A(\M000[10] ),
    .Y(_0790_));
 sky130_fd_sc_hd__mux2_1 _4896_ (.A0(_0789_),
    .A1(_0790_),
    .S(_0706_),
    .X(_0791_));
 sky130_fd_sc_hd__nand2_1 _4897_ (.A(_0791_),
    .B(_0783_),
    .Y(_0792_));
 sky130_fd_sc_hd__o21a_1 _4898_ (.A1(_0783_),
    .A2(_0727_),
    .B1(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _4899_ (.A0(_0793_),
    .A1(_0730_),
    .S(_0871_),
    .X(_0795_));
 sky130_fd_sc_hd__inv_2 _4900_ (.A(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _4901_ (.A(_0796_),
    .B(_0609_),
    .Y(_0797_));
 sky130_fd_sc_hd__o21ai_1 _4902_ (.A1(_0609_),
    .A2(_0733_),
    .B1(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__nand2_1 _4903_ (.A(_0798_),
    .B(_0185_),
    .Y(_0799_));
 sky130_fd_sc_hd__o21ai_1 _4904_ (.A1(_0788_),
    .A2(_0734_),
    .B1(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_0800_),
    .B(_0216_),
    .Y(_0801_));
 sky130_fd_sc_hd__nand2_1 _4906_ (.A(_0787_),
    .B(_0801_),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _4907_ (.A(_0740_),
    .B(_0237_),
    .Y(_0803_));
 sky130_fd_sc_hd__o21ai_1 _4908_ (.A1(_0237_),
    .A2(_0802_),
    .B1(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__buf_2 _4909_ (.A(_0382_),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_1 _4910_ (.A(_0804_),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__nand2_1 _4911_ (.A(_0743_),
    .B(_0259_),
    .Y(_0808_));
 sky130_fd_sc_hd__nand3_1 _4912_ (.A(_0807_),
    .B(_0808_),
    .C(_0429_),
    .Y(_0809_));
 sky130_fd_sc_hd__or2b_1 _4913_ (.A(_0746_),
    .B_N(_0401_),
    .X(_0810_));
 sky130_fd_sc_hd__clkbuf_4 _4914_ (.A(_0474_),
    .X(_0811_));
 sky130_fd_sc_hd__nand3_1 _4915_ (.A(_0809_),
    .B(_0810_),
    .C(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__nand2_1 _4916_ (.A(_0749_),
    .B(_0406_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand3_1 _4917_ (.A(_0812_),
    .B(_0813_),
    .C(_0427_),
    .Y(_0814_));
 sky130_fd_sc_hd__nand3_1 _4918_ (.A(_0751_),
    .B(_0752_),
    .C(_0494_),
    .Y(_0815_));
 sky130_fd_sc_hd__buf_4 _4919_ (.A(_0477_),
    .X(_0817_));
 sky130_fd_sc_hd__nand3_1 _4920_ (.A(_0814_),
    .B(_0815_),
    .C(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nand3_1 _4921_ (.A(_0725_),
    .B(_0753_),
    .C(_0476_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand3_1 _4922_ (.A(_0818_),
    .B(_0819_),
    .C(_0546_),
    .Y(_0820_));
 sky130_fd_sc_hd__buf_4 _4923_ (.A(_0662_),
    .X(_0821_));
 sky130_fd_sc_hd__nand3_1 _4924_ (.A(_0754_),
    .B(_0544_),
    .C(_0756_),
    .Y(_0822_));
 sky130_fd_sc_hd__nand3_1 _4925_ (.A(_0820_),
    .B(_0821_),
    .C(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__nand3_1 _4926_ (.A(_0757_),
    .B(_0759_),
    .C(_0599_),
    .Y(_0824_));
 sky130_fd_sc_hd__nand3_1 _4927_ (.A(_0823_),
    .B(_0637_),
    .C(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(_0786_),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__inv_2 _4929_ (.A(_0711_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _4930_ (.A(_0826_),
    .B(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__nand3_1 _4931_ (.A(_0637_),
    .B(_0762_),
    .C(_0763_),
    .Y(_0830_));
 sky130_fd_sc_hd__nand3_1 _4932_ (.A(_0660_),
    .B(_0692_),
    .C(_0636_),
    .Y(_0831_));
 sky130_fd_sc_hd__nand3_1 _4933_ (.A(_0711_),
    .B(_0830_),
    .C(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_2 _4934_ (.A(_0829_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__nand3_1 _4935_ (.A(_0712_),
    .B(_0713_),
    .C(_0715_),
    .Y(_0834_));
 sky130_fd_sc_hd__nand2_1 _4936_ (.A(_0834_),
    .B(_0694_),
    .Y(_0835_));
 sky130_fd_sc_hd__inv_2 _4937_ (.A(_0765_),
    .Y(_0836_));
 sky130_fd_sc_hd__nand3_2 _4938_ (.A(_0833_),
    .B(_0835_),
    .C(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__inv_2 _4939_ (.A(_0837_),
    .Y(_0839_));
 sky130_fd_sc_hd__nand3_2 _4940_ (.A(_0785_),
    .B(_0839_),
    .C(_0768_),
    .Y(_0840_));
 sky130_fd_sc_hd__inv_2 _4941_ (.A(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__nand3_4 _4942_ (.A(_0781_),
    .B(_0770_),
    .C(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_2 _4943_ (.A(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__nand2_1 _4944_ (.A(_0776_),
    .B(_0770_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand3_2 _4945_ (.A(_0843_),
    .B(_0774_),
    .C(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _4946_ (.A(_0779_),
    .B(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _4947_ (.A(_0774_),
    .B(_0844_),
    .Y(_0847_));
 sky130_fd_sc_hd__nor2_1 _4948_ (.A(_0842_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__nand3_2 _4949_ (.A(_0848_),
    .B(_0778_),
    .C(_0775_),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _4950_ (.A(_0846_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__nand2_1 _4951_ (.A(_0781_),
    .B(_0770_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_1 _4952_ (.A(_0852_),
    .B(_0840_),
    .Y(_0853_));
 sky130_fd_sc_hd__nand2_1 _4953_ (.A(_0785_),
    .B(_0768_),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_1 _4954_ (.A(_0854_),
    .B(_0837_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_1 _4955_ (.A(_0833_),
    .B(_0766_),
    .Y(_0856_));
 sky130_fd_sc_hd__buf_2 _4956_ (.A(_0259_),
    .X(_0857_));
 sky130_fd_sc_hd__nand2_1 _4957_ (.A(_0804_),
    .B(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__mux2_1 _4958_ (.A0(\M000[8] ),
    .A1(\M000[9] ),
    .S(_0695_),
    .X(_0859_));
 sky130_fd_sc_hd__nand2_1 _4959_ (.A(_0859_),
    .B(_0772_),
    .Y(_0861_));
 sky130_fd_sc_hd__o21ai_1 _4960_ (.A1(_0783_),
    .A2(_0791_),
    .B1(_0861_),
    .Y(_0862_));
 sky130_fd_sc_hd__inv_2 _4961_ (.A(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__nand2_1 _4962_ (.A(_0863_),
    .B(_2726_),
    .Y(_0864_));
 sky130_fd_sc_hd__o21a_1 _4963_ (.A1(_2726_),
    .A2(_0793_),
    .B1(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _4964_ (.A0(_0795_),
    .A1(_0865_),
    .S(_0609_),
    .X(_0866_));
 sky130_fd_sc_hd__nand2_1 _4965_ (.A(_0866_),
    .B(_0185_),
    .Y(_0867_));
 sky130_fd_sc_hd__o21ai_1 _4966_ (.A1(_0185_),
    .A2(_0798_),
    .B1(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__or2_1 _4967_ (.A(_0184_),
    .B(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(_0800_),
    .B(_0184_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_1 _4969_ (.A(_0869_),
    .B(_0870_),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_1 _4970_ (.A(_0872_),
    .B(_0676_),
    .Y(_0873_));
 sky130_fd_sc_hd__buf_2 _4971_ (.A(_0237_),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _4972_ (.A(_0802_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__nand3_1 _4973_ (.A(_0873_),
    .B(_0875_),
    .C(_0806_),
    .Y(_0876_));
 sky130_fd_sc_hd__nand3_1 _4974_ (.A(_0858_),
    .B(_0876_),
    .C(_0429_),
    .Y(_0877_));
 sky130_fd_sc_hd__buf_2 _4975_ (.A(_0401_),
    .X(_0878_));
 sky130_fd_sc_hd__nand3_1 _4976_ (.A(_0807_),
    .B(_0808_),
    .C(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nand3_1 _4977_ (.A(_0877_),
    .B(_0879_),
    .C(_0811_),
    .Y(_0880_));
 sky130_fd_sc_hd__buf_2 _4978_ (.A(_0406_),
    .X(_0881_));
 sky130_fd_sc_hd__nand3_1 _4979_ (.A(_0809_),
    .B(_0810_),
    .C(_0881_),
    .Y(_0883_));
 sky130_fd_sc_hd__nand3_1 _4980_ (.A(_0880_),
    .B(_0883_),
    .C(_0427_),
    .Y(_0884_));
 sky130_fd_sc_hd__nand3_1 _4981_ (.A(_0812_),
    .B(_0813_),
    .C(_0494_),
    .Y(_0885_));
 sky130_fd_sc_hd__nand3_1 _4982_ (.A(_0884_),
    .B(_0885_),
    .C(_0817_),
    .Y(_0886_));
 sky130_fd_sc_hd__nand3_1 _4983_ (.A(_0814_),
    .B(_0815_),
    .C(_0476_),
    .Y(_0887_));
 sky130_fd_sc_hd__nand3_1 _4984_ (.A(_0886_),
    .B(_0887_),
    .C(_0546_),
    .Y(_0888_));
 sky130_fd_sc_hd__nand3_1 _4985_ (.A(_0818_),
    .B(_0819_),
    .C(_0544_),
    .Y(_0889_));
 sky130_fd_sc_hd__nand3_1 _4986_ (.A(_0888_),
    .B(_0889_),
    .C(_0821_),
    .Y(_0890_));
 sky130_fd_sc_hd__buf_2 _4987_ (.A(_0599_),
    .X(_0891_));
 sky130_fd_sc_hd__nand3_1 _4988_ (.A(_0820_),
    .B(_0822_),
    .C(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand3_1 _4989_ (.A(_0890_),
    .B(_0892_),
    .C(_0638_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand3_1 _4990_ (.A(_0823_),
    .B(_0824_),
    .C(_0714_),
    .Y(_0895_));
 sky130_fd_sc_hd__nand3_1 _4991_ (.A(_0828_),
    .B(_0894_),
    .C(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__nand3_1 _4992_ (.A(_0712_),
    .B(_0786_),
    .C(_0825_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand3_1 _4993_ (.A(_0896_),
    .B(_0897_),
    .C(_0836_),
    .Y(_0898_));
 sky130_fd_sc_hd__nand2_2 _4994_ (.A(_0856_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _4995_ (.A(_0835_),
    .B(_0766_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_1 _4996_ (.A(_0900_),
    .B(_0767_),
    .Y(_0901_));
 sky130_fd_sc_hd__and2_1 _4997_ (.A(_0830_),
    .B(_0831_),
    .X(_0902_));
 sky130_fd_sc_hd__nand3_2 _4998_ (.A(_0902_),
    .B(_0826_),
    .C(_0828_),
    .Y(_0903_));
 sky130_fd_sc_hd__inv_2 _4999_ (.A(_0903_),
    .Y(_0905_));
 sky130_fd_sc_hd__buf_4 _5000_ (.A(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__nand3_2 _5001_ (.A(_0899_),
    .B(_0901_),
    .C(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__inv_2 _5002_ (.A(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__nand3_2 _5003_ (.A(_0855_),
    .B(_0908_),
    .C(_0840_),
    .Y(_0909_));
 sky130_fd_sc_hd__inv_2 _5004_ (.A(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand3_2 _5005_ (.A(_0853_),
    .B(_0842_),
    .C(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__inv_2 _5006_ (.A(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__nand2_1 _5007_ (.A(_0776_),
    .B(_0771_),
    .Y(_0913_));
 sky130_fd_sc_hd__nand3_1 _5008_ (.A(_0702_),
    .B(_0770_),
    .C(_0773_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand3_1 _5009_ (.A(_0913_),
    .B(_0842_),
    .C(_0914_),
    .Y(_0916_));
 sky130_fd_sc_hd__nand3_1 _5010_ (.A(_0912_),
    .B(_0845_),
    .C(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__nand2_1 _5011_ (.A(_0851_),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__nand2_1 _5012_ (.A(_0845_),
    .B(_0916_),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_1 _5013_ (.A(_0911_),
    .B(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__nand3_2 _5014_ (.A(_0920_),
    .B(_0846_),
    .C(_0850_),
    .Y(_0921_));
 sky130_fd_sc_hd__nand2_1 _5015_ (.A(_0918_),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(_0896_),
    .B(_0897_),
    .Y(_0923_));
 sky130_fd_sc_hd__inv_2 _5017_ (.A(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__buf_4 _5018_ (.A(_0836_),
    .X(_0925_));
 sky130_fd_sc_hd__nand3_4 _5019_ (.A(_0924_),
    .B(_0925_),
    .C(_0833_),
    .Y(_0927_));
 sky130_fd_sc_hd__nand2_1 _5020_ (.A(_0901_),
    .B(_0903_),
    .Y(_0928_));
 sky130_fd_sc_hd__nand3b_1 _5021_ (.A_N(_0854_),
    .B(_0837_),
    .C(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_1 _5022_ (.A(_0927_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand3_2 _5023_ (.A(_0853_),
    .B(_0930_),
    .C(_0842_),
    .Y(_0931_));
 sky130_fd_sc_hd__inv_2 _5024_ (.A(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__nand2_1 _5025_ (.A(_0919_),
    .B(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand3_1 _5026_ (.A(_0845_),
    .B(_0931_),
    .C(_0916_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _5027_ (.A(_0933_),
    .B(_0934_),
    .Y(_0935_));
 sky130_fd_sc_hd__nand2_1 _5028_ (.A(_0855_),
    .B(_0840_),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2_1 _5029_ (.A(_0936_),
    .B(_0907_),
    .Y(_0938_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_0928_),
    .B(_0837_),
    .Y(_0939_));
 sky130_fd_sc_hd__nand2_1 _5031_ (.A(_0939_),
    .B(_0927_),
    .Y(_0940_));
 sky130_fd_sc_hd__nand2_1 _5032_ (.A(_0940_),
    .B(_0907_),
    .Y(_0941_));
 sky130_fd_sc_hd__inv_2 _5033_ (.A(_0941_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(_0924_),
    .B(_0766_),
    .Y(_0943_));
 sky130_fd_sc_hd__buf_6 _5035_ (.A(_0828_),
    .X(_0944_));
 sky130_fd_sc_hd__inv_2 _5036_ (.A(\M000[7] ),
    .Y(_0945_));
 sky130_fd_sc_hd__inv_2 _5037_ (.A(\M000[8] ),
    .Y(_0946_));
 sky130_fd_sc_hd__mux2_1 _5038_ (.A0(_0945_),
    .A1(_0946_),
    .S(_0695_),
    .X(_0947_));
 sky130_fd_sc_hd__nand2_1 _5039_ (.A(_0947_),
    .B(_0772_),
    .Y(_0949_));
 sky130_fd_sc_hd__o21a_1 _5040_ (.A1(_0772_),
    .A2(_0859_),
    .B1(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__mux2_1 _5041_ (.A0(_0950_),
    .A1(_0862_),
    .S(_0871_),
    .X(_0951_));
 sky130_fd_sc_hd__inv_2 _5042_ (.A(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__nand2_1 _5043_ (.A(_0952_),
    .B(_0609_),
    .Y(_0953_));
 sky130_fd_sc_hd__o21a_1 _5044_ (.A1(_0609_),
    .A2(_0865_),
    .B1(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__inv_2 _5045_ (.A(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _5046_ (.A(_0955_),
    .B(_0788_),
    .Y(_0956_));
 sky130_fd_sc_hd__o21a_1 _5047_ (.A1(_0788_),
    .A2(_0866_),
    .B1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__inv_2 _5048_ (.A(_0957_),
    .Y(_0958_));
 sky130_fd_sc_hd__clkbuf_4 _5049_ (.A(_0216_),
    .X(_0960_));
 sky130_fd_sc_hd__nand2_1 _5050_ (.A(_0958_),
    .B(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__or2_1 _5051_ (.A(_0216_),
    .B(_0868_),
    .X(_0962_));
 sky130_fd_sc_hd__nand2_1 _5052_ (.A(_0961_),
    .B(_0962_),
    .Y(_0963_));
 sky130_fd_sc_hd__nand2_1 _5053_ (.A(_0963_),
    .B(_0676_),
    .Y(_0964_));
 sky130_fd_sc_hd__nand2_1 _5054_ (.A(_0872_),
    .B(_0874_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand3_1 _5055_ (.A(_0964_),
    .B(_0965_),
    .C(_0806_),
    .Y(_0966_));
 sky130_fd_sc_hd__nand3_1 _5056_ (.A(_0873_),
    .B(_0875_),
    .C(_0857_),
    .Y(_0967_));
 sky130_fd_sc_hd__nand3_1 _5057_ (.A(_0966_),
    .B(_0429_),
    .C(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__nand3_1 _5058_ (.A(_0858_),
    .B(_0876_),
    .C(_0878_),
    .Y(_0969_));
 sky130_fd_sc_hd__nand3_1 _5059_ (.A(_0968_),
    .B(_0969_),
    .C(_0811_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand3_1 _5060_ (.A(_0877_),
    .B(_0879_),
    .C(_0881_),
    .Y(_0972_));
 sky130_fd_sc_hd__nand3_1 _5061_ (.A(_0971_),
    .B(_0972_),
    .C(_0427_),
    .Y(_0973_));
 sky130_fd_sc_hd__nand3_1 _5062_ (.A(_0880_),
    .B(_0883_),
    .C(_0494_),
    .Y(_0974_));
 sky130_fd_sc_hd__nand3_1 _5063_ (.A(_0973_),
    .B(_0974_),
    .C(_0817_),
    .Y(_0975_));
 sky130_fd_sc_hd__nand3_1 _5064_ (.A(_0884_),
    .B(_0885_),
    .C(_0491_),
    .Y(_0976_));
 sky130_fd_sc_hd__nand3_1 _5065_ (.A(_0975_),
    .B(_0976_),
    .C(_0546_),
    .Y(_0977_));
 sky130_fd_sc_hd__nand3_1 _5066_ (.A(_0886_),
    .B(_0887_),
    .C(_0544_),
    .Y(_0978_));
 sky130_fd_sc_hd__nand3_1 _5067_ (.A(_0977_),
    .B(_0978_),
    .C(_0821_),
    .Y(_0979_));
 sky130_fd_sc_hd__nand3_1 _5068_ (.A(_0888_),
    .B(_0889_),
    .C(_0891_),
    .Y(_0980_));
 sky130_fd_sc_hd__nand3_1 _5069_ (.A(_0979_),
    .B(_0980_),
    .C(_0638_),
    .Y(_0982_));
 sky130_fd_sc_hd__nand3_1 _5070_ (.A(_0890_),
    .B(_0892_),
    .C(_0714_),
    .Y(_0983_));
 sky130_fd_sc_hd__nand3_1 _5071_ (.A(_0944_),
    .B(_0982_),
    .C(_0983_),
    .Y(_0984_));
 sky130_fd_sc_hd__nand3_1 _5072_ (.A(_0894_),
    .B(_0712_),
    .C(_0895_),
    .Y(_0985_));
 sky130_fd_sc_hd__nand3_1 _5073_ (.A(_0984_),
    .B(_0836_),
    .C(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__nand2_1 _5074_ (.A(_0943_),
    .B(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__nand3_2 _5075_ (.A(_0987_),
    .B(_0906_),
    .C(_0899_),
    .Y(_0988_));
 sky130_fd_sc_hd__inv_2 _5076_ (.A(_0988_),
    .Y(_0989_));
 sky130_fd_sc_hd__nand3_1 _5077_ (.A(_0938_),
    .B(_0942_),
    .C(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__buf_2 _5078_ (.A(_0903_),
    .X(_0991_));
 sky130_fd_sc_hd__nand3b_1 _5079_ (.A_N(_0784_),
    .B(_0767_),
    .C(_0900_),
    .Y(_0993_));
 sky130_fd_sc_hd__nor2_1 _5080_ (.A(_0991_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__nand3_1 _5081_ (.A(_0781_),
    .B(_0994_),
    .C(_0770_),
    .Y(_0995_));
 sky130_fd_sc_hd__nand2_1 _5082_ (.A(_0853_),
    .B(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_0996_),
    .B(_0909_),
    .Y(_0997_));
 sky130_fd_sc_hd__nand3b_1 _5084_ (.A_N(_0990_),
    .B(_0997_),
    .C(_0931_),
    .Y(_0998_));
 sky130_fd_sc_hd__inv_2 _5085_ (.A(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(_0935_),
    .B(_0999_),
    .Y(_1000_));
 sky130_fd_sc_hd__nand2_1 _5087_ (.A(_0922_),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__nand2_1 _5088_ (.A(_0919_),
    .B(_0911_),
    .Y(_1002_));
 sky130_fd_sc_hd__nand2_1 _5089_ (.A(_0917_),
    .B(_1002_),
    .Y(_1004_));
 sky130_fd_sc_hd__nor2_1 _5090_ (.A(_0998_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__nand3_2 _5091_ (.A(_1005_),
    .B(_0918_),
    .C(_0921_),
    .Y(_1006_));
 sky130_fd_sc_hd__nand2_1 _5092_ (.A(_1001_),
    .B(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__nand2_1 _5093_ (.A(_0997_),
    .B(_0931_),
    .Y(_1008_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_1008_),
    .B(_0990_),
    .Y(_1009_));
 sky130_fd_sc_hd__buf_4 _5095_ (.A(_0988_),
    .X(_1010_));
 sky130_fd_sc_hd__nand3_1 _5096_ (.A(_0938_),
    .B(_0942_),
    .C(_0909_),
    .Y(_1011_));
 sky130_fd_sc_hd__nor2_1 _5097_ (.A(_1010_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__nand3_2 _5098_ (.A(_0997_),
    .B(_1012_),
    .C(_0911_),
    .Y(_1013_));
 sky130_fd_sc_hd__nand2_1 _5099_ (.A(_1009_),
    .B(_1013_),
    .Y(_1015_));
 sky130_fd_sc_hd__inv_2 _5100_ (.A(_0899_),
    .Y(_1016_));
 sky130_fd_sc_hd__nand2_1 _5101_ (.A(_1016_),
    .B(_0991_),
    .Y(_1017_));
 sky130_fd_sc_hd__nand3_1 _5102_ (.A(_0943_),
    .B(_0905_),
    .C(_0986_),
    .Y(_1018_));
 sky130_fd_sc_hd__and2_1 _5103_ (.A(_1017_),
    .B(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__nand2_1 _5104_ (.A(_0957_),
    .B(_0184_),
    .Y(_1020_));
 sky130_fd_sc_hd__inv_2 _5105_ (.A(\M000[6] ),
    .Y(_1021_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(_1021_),
    .A1(_0945_),
    .S(_0706_),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(_0947_),
    .A1(_1022_),
    .S(_0783_),
    .X(_1023_));
 sky130_fd_sc_hd__nand2_1 _5108_ (.A(_1023_),
    .B(_2726_),
    .Y(_1024_));
 sky130_fd_sc_hd__o21a_1 _5109_ (.A1(_2726_),
    .A2(_0950_),
    .B1(_1024_),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_1 _5110_ (.A0(_1026_),
    .A1(_0951_),
    .S(_2733_),
    .X(_1027_));
 sky130_fd_sc_hd__mux2_1 _5111_ (.A0(_0954_),
    .A1(_1027_),
    .S(_0788_),
    .X(_1028_));
 sky130_fd_sc_hd__nand2_1 _5112_ (.A(_1028_),
    .B(_0216_),
    .Y(_1029_));
 sky130_fd_sc_hd__nand2_1 _5113_ (.A(_1020_),
    .B(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__inv_2 _5114_ (.A(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__nand2_1 _5115_ (.A(_1031_),
    .B(_0676_),
    .Y(_1032_));
 sky130_fd_sc_hd__nand2_1 _5116_ (.A(_0963_),
    .B(_0874_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand3_1 _5117_ (.A(_1032_),
    .B(_1033_),
    .C(_0806_),
    .Y(_1034_));
 sky130_fd_sc_hd__nand3_1 _5118_ (.A(_0964_),
    .B(_0965_),
    .C(_0857_),
    .Y(_1035_));
 sky130_fd_sc_hd__nand3_1 _5119_ (.A(_1034_),
    .B(_1035_),
    .C(_0429_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand3_1 _5120_ (.A(_0966_),
    .B(_0878_),
    .C(_0967_),
    .Y(_1038_));
 sky130_fd_sc_hd__nand3_1 _5121_ (.A(_1037_),
    .B(_1038_),
    .C(_0811_),
    .Y(_1039_));
 sky130_fd_sc_hd__nand3_1 _5122_ (.A(_0968_),
    .B(_0969_),
    .C(_0881_),
    .Y(_1040_));
 sky130_fd_sc_hd__clkbuf_4 _5123_ (.A(_0427_),
    .X(_1041_));
 sky130_fd_sc_hd__nand3_1 _5124_ (.A(_1039_),
    .B(_1040_),
    .C(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__nand3_1 _5125_ (.A(_0971_),
    .B(_0972_),
    .C(_0494_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand3_1 _5126_ (.A(_1042_),
    .B(_1043_),
    .C(_0817_),
    .Y(_1044_));
 sky130_fd_sc_hd__nand3_1 _5127_ (.A(_0973_),
    .B(_0974_),
    .C(_0491_),
    .Y(_1045_));
 sky130_fd_sc_hd__buf_2 _5128_ (.A(_0546_),
    .X(_1046_));
 sky130_fd_sc_hd__nand3_1 _5129_ (.A(_1044_),
    .B(_1045_),
    .C(_1046_),
    .Y(_1048_));
 sky130_fd_sc_hd__nand3_1 _5130_ (.A(_0975_),
    .B(_0976_),
    .C(_0544_),
    .Y(_1049_));
 sky130_fd_sc_hd__nand3_1 _5131_ (.A(_1048_),
    .B(_1049_),
    .C(_0821_),
    .Y(_1050_));
 sky130_fd_sc_hd__nand3_1 _5132_ (.A(_0977_),
    .B(_0978_),
    .C(_0891_),
    .Y(_1051_));
 sky130_fd_sc_hd__nand3_1 _5133_ (.A(_1050_),
    .B(_1051_),
    .C(_0638_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand3_1 _5134_ (.A(_0979_),
    .B(_0980_),
    .C(_0714_),
    .Y(_1053_));
 sky130_fd_sc_hd__nand3_1 _5135_ (.A(_0944_),
    .B(_1052_),
    .C(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__nand3_1 _5136_ (.A(_0982_),
    .B(_0983_),
    .C(_0712_),
    .Y(_1055_));
 sky130_fd_sc_hd__nand3_1 _5137_ (.A(_1054_),
    .B(_1055_),
    .C(_0836_),
    .Y(_1056_));
 sky130_fd_sc_hd__nand3_1 _5138_ (.A(_0984_),
    .B(_0766_),
    .C(_0985_),
    .Y(_1057_));
 sky130_fd_sc_hd__a21o_1 _5139_ (.A1(_1056_),
    .A2(_1057_),
    .B1(_0903_),
    .X(_1059_));
 sky130_fd_sc_hd__nand2_1 _5140_ (.A(_0987_),
    .B(_0991_),
    .Y(_1060_));
 sky130_fd_sc_hd__nand2_1 _5141_ (.A(_1059_),
    .B(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__inv_6 _5142_ (.A(_0927_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand3_4 _5143_ (.A(_1019_),
    .B(_1061_),
    .C(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__nand2_1 _5144_ (.A(_0942_),
    .B(_0989_),
    .Y(_1064_));
 sky130_fd_sc_hd__nand2_1 _5145_ (.A(_0941_),
    .B(_0988_),
    .Y(_1065_));
 sky130_fd_sc_hd__nand2_2 _5146_ (.A(_1064_),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__nand2_1 _5147_ (.A(_0938_),
    .B(_0909_),
    .Y(_1067_));
 sky130_fd_sc_hd__nand2_1 _5148_ (.A(_1067_),
    .B(_1064_),
    .Y(_1068_));
 sky130_fd_sc_hd__nand2_1 _5149_ (.A(_1068_),
    .B(_0990_),
    .Y(_1070_));
 sky130_fd_sc_hd__or2_1 _5150_ (.A(_1066_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__inv_2 _5151_ (.A(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__nand2_1 _5152_ (.A(_0935_),
    .B(_1072_),
    .Y(_1073_));
 sky130_fd_sc_hd__nor3_1 _5153_ (.A(_1015_),
    .B(_1063_),
    .C(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__inv_2 _5154_ (.A(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__nand2_1 _5155_ (.A(_1007_),
    .B(_1075_),
    .Y(_1076_));
 sky130_fd_sc_hd__inv_2 _5156_ (.A(_1066_),
    .Y(_1077_));
 sky130_fd_sc_hd__inv_2 _5157_ (.A(_1067_),
    .Y(_1078_));
 sky130_fd_sc_hd__inv_2 _5158_ (.A(_1063_),
    .Y(_1079_));
 sky130_fd_sc_hd__buf_6 _5159_ (.A(_1079_),
    .X(_1081_));
 sky130_fd_sc_hd__nand3_2 _5160_ (.A(_1077_),
    .B(_1078_),
    .C(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__inv_2 _5161_ (.A(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__nand3_4 _5162_ (.A(_1009_),
    .B(_1013_),
    .C(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__nor2_1 _5163_ (.A(_1004_),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__nand3_1 _5164_ (.A(_1001_),
    .B(_1006_),
    .C(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__nand2_1 _5165_ (.A(_1076_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__nand3_1 _5166_ (.A(_0933_),
    .B(_1013_),
    .C(_0934_),
    .Y(_1088_));
 sky130_fd_sc_hd__nand2_1 _5167_ (.A(_1000_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__inv_2 _5168_ (.A(_1084_),
    .Y(_1090_));
 sky130_fd_sc_hd__nand2_1 _5169_ (.A(_1089_),
    .B(_1090_),
    .Y(_1092_));
 sky130_fd_sc_hd__nand3_1 _5170_ (.A(_1000_),
    .B(_1084_),
    .C(_1088_),
    .Y(_1093_));
 sky130_fd_sc_hd__nand2_1 _5171_ (.A(_1092_),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__nand2_1 _5172_ (.A(_1015_),
    .B(_1082_),
    .Y(_1095_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(_1061_),
    .B(_0927_),
    .Y(_1096_));
 sky130_fd_sc_hd__or2b_1 _5174_ (.A(_1028_),
    .B_N(_0184_),
    .X(_1097_));
 sky130_fd_sc_hd__mux2_1 _5175_ (.A0(net159),
    .A1(\M000[6] ),
    .S(_0706_),
    .X(_1098_));
 sky130_fd_sc_hd__nand2_1 _5176_ (.A(net160),
    .B(_0783_),
    .Y(_1099_));
 sky130_fd_sc_hd__o21ai_1 _5177_ (.A1(_0783_),
    .A2(_1022_),
    .B1(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__nand2_1 _5178_ (.A(_1023_),
    .B(_0871_),
    .Y(_1101_));
 sky130_fd_sc_hd__o21ai_1 _5179_ (.A1(_0871_),
    .A2(net161),
    .B1(_1101_),
    .Y(_1103_));
 sky130_fd_sc_hd__nand2_1 _5180_ (.A(net162),
    .B(_0609_),
    .Y(_1104_));
 sky130_fd_sc_hd__o21ai_1 _5181_ (.A1(_0609_),
    .A2(_1026_),
    .B1(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__nand2_1 _5182_ (.A(net163),
    .B(_0788_),
    .Y(_1106_));
 sky130_fd_sc_hd__o21ai_1 _5183_ (.A1(_0788_),
    .A2(_1027_),
    .B1(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__nand2_1 _5184_ (.A(_1107_),
    .B(_0960_),
    .Y(_1108_));
 sky130_fd_sc_hd__nand2_1 _5185_ (.A(_1097_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__nand2_1 _5186_ (.A(_1030_),
    .B(_0874_),
    .Y(_1110_));
 sky130_fd_sc_hd__o21ai_1 _5187_ (.A1(_0874_),
    .A2(_1109_),
    .B1(_1110_),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_1 _5188_ (.A(_1111_),
    .B(_0806_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand3_1 _5189_ (.A(_1032_),
    .B(_1033_),
    .C(_0857_),
    .Y(_1114_));
 sky130_fd_sc_hd__nand3_1 _5190_ (.A(_1112_),
    .B(_0429_),
    .C(_1114_),
    .Y(_1115_));
 sky130_fd_sc_hd__nand3_1 _5191_ (.A(_1034_),
    .B(_1035_),
    .C(_0878_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand3_1 _5192_ (.A(_1115_),
    .B(_1116_),
    .C(_0811_),
    .Y(_1117_));
 sky130_fd_sc_hd__nand3_1 _5193_ (.A(_1037_),
    .B(_1038_),
    .C(_0881_),
    .Y(_1118_));
 sky130_fd_sc_hd__nand3_1 _5194_ (.A(_1117_),
    .B(_1118_),
    .C(_1041_),
    .Y(_1119_));
 sky130_fd_sc_hd__nand3_1 _5195_ (.A(_1039_),
    .B(_1040_),
    .C(_0494_),
    .Y(_1120_));
 sky130_fd_sc_hd__nand3_1 _5196_ (.A(_1119_),
    .B(_1120_),
    .C(_0817_),
    .Y(_1121_));
 sky130_fd_sc_hd__nand3_1 _5197_ (.A(_1042_),
    .B(_1043_),
    .C(_0491_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand3_1 _5198_ (.A(_1121_),
    .B(_1122_),
    .C(_1046_),
    .Y(_1123_));
 sky130_fd_sc_hd__nand3_1 _5199_ (.A(_1044_),
    .B(_1045_),
    .C(_0544_),
    .Y(_1125_));
 sky130_fd_sc_hd__nand3_1 _5200_ (.A(_1123_),
    .B(_1125_),
    .C(_0821_),
    .Y(_1126_));
 sky130_fd_sc_hd__nand3_1 _5201_ (.A(_1048_),
    .B(_1049_),
    .C(_0891_),
    .Y(_1127_));
 sky130_fd_sc_hd__nand3_1 _5202_ (.A(_1126_),
    .B(_1127_),
    .C(_0638_),
    .Y(_1128_));
 sky130_fd_sc_hd__nand3_1 _5203_ (.A(_1050_),
    .B(_1051_),
    .C(_0714_),
    .Y(_1129_));
 sky130_fd_sc_hd__nand3_1 _5204_ (.A(_1128_),
    .B(_0944_),
    .C(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__nand3_1 _5205_ (.A(_1052_),
    .B(_1053_),
    .C(_0712_),
    .Y(_1131_));
 sky130_fd_sc_hd__nand3_1 _5206_ (.A(_1130_),
    .B(_1131_),
    .C(_0925_),
    .Y(_1132_));
 sky130_fd_sc_hd__nand3_1 _5207_ (.A(_1054_),
    .B(_1055_),
    .C(_0766_),
    .Y(_1133_));
 sky130_fd_sc_hd__nand3_1 _5208_ (.A(_1132_),
    .B(_1133_),
    .C(_0906_),
    .Y(_1134_));
 sky130_fd_sc_hd__nand3_1 _5209_ (.A(_1056_),
    .B(_1057_),
    .C(_0991_),
    .Y(_1136_));
 sky130_fd_sc_hd__nand3_1 _5210_ (.A(_1062_),
    .B(_1134_),
    .C(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__nand2_2 _5211_ (.A(_1096_),
    .B(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__nand2_1 _5212_ (.A(_1138_),
    .B(_0989_),
    .Y(_1139_));
 sky130_fd_sc_hd__nand2_1 _5213_ (.A(_1056_),
    .B(_1057_),
    .Y(_1140_));
 sky130_fd_sc_hd__nand3_1 _5214_ (.A(_0943_),
    .B(_0991_),
    .C(_0986_),
    .Y(_1141_));
 sky130_fd_sc_hd__o211ai_1 _5215_ (.A1(_0991_),
    .A2(_1140_),
    .B1(_1062_),
    .C1(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__nand3_1 _5216_ (.A(_1017_),
    .B(_1018_),
    .C(_0927_),
    .Y(_1143_));
 sky130_fd_sc_hd__nand2_2 _5217_ (.A(_1142_),
    .B(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__nand2_1 _5218_ (.A(_1144_),
    .B(_1010_),
    .Y(_1145_));
 sky130_fd_sc_hd__nand2_2 _5219_ (.A(_1139_),
    .B(_1145_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand3_2 _5220_ (.A(_1147_),
    .B(_1066_),
    .C(_1079_),
    .Y(_1148_));
 sky130_fd_sc_hd__or2_1 _5221_ (.A(_1070_),
    .B(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__inv_2 _5222_ (.A(_1149_),
    .Y(_1150_));
 sky130_fd_sc_hd__nand3_4 _5223_ (.A(_1095_),
    .B(_1084_),
    .C(_1150_),
    .Y(_1151_));
 sky130_fd_sc_hd__inv_2 _5224_ (.A(_1151_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _5225_ (.A(_1094_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__nand2_1 _5226_ (.A(_1087_),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__a21oi_1 _5227_ (.A1(_1092_),
    .A2(_1093_),
    .B1(_1151_),
    .Y(_1155_));
 sky130_fd_sc_hd__nand3_2 _5228_ (.A(_1155_),
    .B(_1076_),
    .C(_1086_),
    .Y(_1156_));
 sky130_fd_sc_hd__nand2_1 _5229_ (.A(_1154_),
    .B(_1156_),
    .Y(_1158_));
 sky130_fd_sc_hd__nand2_1 _5230_ (.A(_1095_),
    .B(_1084_),
    .Y(_1159_));
 sky130_fd_sc_hd__nand2_1 _5231_ (.A(_1159_),
    .B(_1149_),
    .Y(_1160_));
 sky130_fd_sc_hd__nand2_1 _5232_ (.A(_1077_),
    .B(_1079_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _5233_ (.A(_1161_),
    .B(_1070_),
    .Y(_1162_));
 sky130_fd_sc_hd__nand2_1 _5234_ (.A(_1162_),
    .B(_1082_),
    .Y(_1163_));
 sky130_fd_sc_hd__inv_2 _5235_ (.A(_1148_),
    .Y(_1164_));
 sky130_fd_sc_hd__nand2_1 _5236_ (.A(_1163_),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__nand3_1 _5237_ (.A(_1162_),
    .B(_1148_),
    .C(_1082_),
    .Y(_1166_));
 sky130_fd_sc_hd__nand2_1 _5238_ (.A(_1165_),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__nand2_1 _5239_ (.A(_1147_),
    .B(_1063_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _5240_ (.A(_1138_),
    .B(_1010_),
    .Y(_1170_));
 sky130_fd_sc_hd__nand2_1 _5241_ (.A(_1111_),
    .B(_0857_),
    .Y(_1171_));
 sky130_fd_sc_hd__nand2_1 _5242_ (.A(_1109_),
    .B(_0874_),
    .Y(_1172_));
 sky130_fd_sc_hd__nand2_1 _5243_ (.A(_1107_),
    .B(_0184_),
    .Y(_1173_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(net148),
    .A1(\M000[5] ),
    .S(_0706_),
    .X(_1174_));
 sky130_fd_sc_hd__mux2_1 _5245_ (.A0(net149),
    .A1(net160),
    .S(_2719_),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _5246_ (.A0(_1175_),
    .A1(net161),
    .S(_0871_),
    .X(_1176_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(net162),
    .B(_2733_),
    .Y(_1177_));
 sky130_fd_sc_hd__o21a_1 _5248_ (.A1(_2733_),
    .A2(_1176_),
    .B1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__nand2_1 _5249_ (.A(net163),
    .B(_0198_),
    .Y(_1180_));
 sky130_fd_sc_hd__o21ai_1 _5250_ (.A1(_0198_),
    .A2(_1178_),
    .B1(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__nand2_1 _5251_ (.A(_1181_),
    .B(_0960_),
    .Y(_1182_));
 sky130_fd_sc_hd__nand2_1 _5252_ (.A(_1173_),
    .B(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_1 _5253_ (.A(_1183_),
    .B(_0676_),
    .Y(_1184_));
 sky130_fd_sc_hd__nand3_1 _5254_ (.A(_1172_),
    .B(_1184_),
    .C(_0806_),
    .Y(_1185_));
 sky130_fd_sc_hd__nand3_1 _5255_ (.A(_1171_),
    .B(_1185_),
    .C(_0429_),
    .Y(_1186_));
 sky130_fd_sc_hd__nand3_1 _5256_ (.A(_1112_),
    .B(_0878_),
    .C(_1114_),
    .Y(_1187_));
 sky130_fd_sc_hd__nand3_1 _5257_ (.A(_1186_),
    .B(_1187_),
    .C(_0811_),
    .Y(_1188_));
 sky130_fd_sc_hd__nand3_1 _5258_ (.A(_1115_),
    .B(_1116_),
    .C(_0881_),
    .Y(_1189_));
 sky130_fd_sc_hd__nand3_1 _5259_ (.A(_1188_),
    .B(_1189_),
    .C(_1041_),
    .Y(_1191_));
 sky130_fd_sc_hd__nand3_1 _5260_ (.A(_1117_),
    .B(_1118_),
    .C(_0494_),
    .Y(_1192_));
 sky130_fd_sc_hd__nand3_1 _5261_ (.A(_1191_),
    .B(_1192_),
    .C(_0817_),
    .Y(_1193_));
 sky130_fd_sc_hd__nand3_1 _5262_ (.A(_1119_),
    .B(_1120_),
    .C(_0491_),
    .Y(_1194_));
 sky130_fd_sc_hd__nand3_1 _5263_ (.A(_1193_),
    .B(_1194_),
    .C(_1046_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand3_1 _5264_ (.A(_1121_),
    .B(_1122_),
    .C(_0544_),
    .Y(_1196_));
 sky130_fd_sc_hd__nand3_1 _5265_ (.A(_1195_),
    .B(_1196_),
    .C(_0821_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand3_1 _5266_ (.A(_1123_),
    .B(_1125_),
    .C(_0891_),
    .Y(_1198_));
 sky130_fd_sc_hd__clkbuf_4 _5267_ (.A(_0638_),
    .X(_1199_));
 sky130_fd_sc_hd__nand3_1 _5268_ (.A(_1197_),
    .B(_1198_),
    .C(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nand3_1 _5269_ (.A(_1126_),
    .B(_1127_),
    .C(_0714_),
    .Y(_1202_));
 sky130_fd_sc_hd__nand3_1 _5270_ (.A(_1200_),
    .B(_1202_),
    .C(_0944_),
    .Y(_1203_));
 sky130_fd_sc_hd__nand3_1 _5271_ (.A(_1128_),
    .B(_1129_),
    .C(_0712_),
    .Y(_1204_));
 sky130_fd_sc_hd__nand3_1 _5272_ (.A(_1203_),
    .B(_1204_),
    .C(_0925_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand3_1 _5273_ (.A(_1130_),
    .B(_1131_),
    .C(_0766_),
    .Y(_1206_));
 sky130_fd_sc_hd__nand3_1 _5274_ (.A(_1205_),
    .B(_1206_),
    .C(_0906_),
    .Y(_1207_));
 sky130_fd_sc_hd__nand3_1 _5275_ (.A(_1132_),
    .B(_1133_),
    .C(_0991_),
    .Y(_1208_));
 sky130_fd_sc_hd__nand3_1 _5276_ (.A(_1062_),
    .B(_1207_),
    .C(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand3_1 _5277_ (.A(_1134_),
    .B(_1136_),
    .C(_0927_),
    .Y(_1210_));
 sky130_fd_sc_hd__a21o_1 _5278_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1010_),
    .X(_1211_));
 sky130_fd_sc_hd__nand2_2 _5279_ (.A(_1170_),
    .B(_1211_),
    .Y(_1213_));
 sky130_fd_sc_hd__nand2_1 _5280_ (.A(_1213_),
    .B(_1081_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand2_1 _5281_ (.A(_1169_),
    .B(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand2_1 _5282_ (.A(_1066_),
    .B(_1063_),
    .Y(_1216_));
 sky130_fd_sc_hd__nand2_1 _5283_ (.A(_1161_),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__nand3_4 _5284_ (.A(_1138_),
    .B(_1144_),
    .C(_0989_),
    .Y(_1218_));
 sky130_fd_sc_hd__inv_2 _5285_ (.A(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__nand3_2 _5286_ (.A(_1215_),
    .B(_1217_),
    .C(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__inv_2 _5287_ (.A(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__nand2_2 _5288_ (.A(_1167_),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__inv_2 _5289_ (.A(_1222_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand3_4 _5290_ (.A(_1160_),
    .B(_1224_),
    .C(_1151_),
    .Y(_1225_));
 sky130_fd_sc_hd__inv_2 _5291_ (.A(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__nand3_1 _5292_ (.A(_1092_),
    .B(_1151_),
    .C(_1093_),
    .Y(_1227_));
 sky130_fd_sc_hd__nand3_2 _5293_ (.A(_1226_),
    .B(_1153_),
    .C(_1227_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _5294_ (.A(_1158_),
    .B(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__nand2_1 _5295_ (.A(_1153_),
    .B(_1227_),
    .Y(_1230_));
 sky130_fd_sc_hd__nor2_1 _5296_ (.A(_1225_),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__nand3_2 _5297_ (.A(_1231_),
    .B(_1154_),
    .C(_1156_),
    .Y(_1232_));
 sky130_fd_sc_hd__nand2_1 _5298_ (.A(_1229_),
    .B(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__nand2_1 _5299_ (.A(_1160_),
    .B(_1151_),
    .Y(_1235_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(_1235_),
    .B(_1222_),
    .Y(_1236_));
 sky130_fd_sc_hd__nand2_1 _5301_ (.A(_1217_),
    .B(_1218_),
    .Y(_1237_));
 sky130_fd_sc_hd__nand2_1 _5302_ (.A(_1237_),
    .B(_1148_),
    .Y(_1238_));
 sky130_fd_sc_hd__nand2_1 _5303_ (.A(_1213_),
    .B(_1063_),
    .Y(_1239_));
 sky130_fd_sc_hd__nand3_1 _5304_ (.A(_1209_),
    .B(_1210_),
    .C(_1010_),
    .Y(_1240_));
 sky130_fd_sc_hd__nand3_1 _5305_ (.A(_1186_),
    .B(_1187_),
    .C(_0881_),
    .Y(_1241_));
 sky130_fd_sc_hd__nand3_1 _5306_ (.A(_1171_),
    .B(_1185_),
    .C(_0878_),
    .Y(_1242_));
 sky130_fd_sc_hd__nand3_1 _5307_ (.A(_1172_),
    .B(_1184_),
    .C(_0857_),
    .Y(_1243_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(net139),
    .A1(net148),
    .S(_0706_),
    .X(_1244_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net149),
    .A1(_1244_),
    .S(_0783_),
    .X(_1246_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(net150),
    .A1(_1175_),
    .S(_0871_),
    .X(_1247_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(_1247_),
    .A1(_1176_),
    .S(_2733_),
    .X(_1248_));
 sky130_fd_sc_hd__or2_1 _5312_ (.A(_0788_),
    .B(_1178_),
    .X(_1249_));
 sky130_fd_sc_hd__o21ai_1 _5313_ (.A1(_0198_),
    .A2(_1248_),
    .B1(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__nand2_1 _5314_ (.A(_1250_),
    .B(_0960_),
    .Y(_1251_));
 sky130_fd_sc_hd__nand2_1 _5315_ (.A(_1181_),
    .B(_0184_),
    .Y(_1252_));
 sky130_fd_sc_hd__nand2_1 _5316_ (.A(_1251_),
    .B(_1252_),
    .Y(_1253_));
 sky130_fd_sc_hd__nand2_1 _5317_ (.A(_1253_),
    .B(_0676_),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _5318_ (.A(_1183_),
    .B(_0874_),
    .Y(_1255_));
 sky130_fd_sc_hd__and2_1 _5319_ (.A(_1254_),
    .B(_1255_),
    .X(_1257_));
 sky130_fd_sc_hd__nand2_1 _5320_ (.A(_1257_),
    .B(_0806_),
    .Y(_1258_));
 sky130_fd_sc_hd__nand3_1 _5321_ (.A(_1243_),
    .B(_1258_),
    .C(_0429_),
    .Y(_1259_));
 sky130_fd_sc_hd__nand3_1 _5322_ (.A(_1242_),
    .B(_1259_),
    .C(_0811_),
    .Y(_1260_));
 sky130_fd_sc_hd__nand3_1 _5323_ (.A(_1241_),
    .B(_1260_),
    .C(_1041_),
    .Y(_1261_));
 sky130_fd_sc_hd__nand3_1 _5324_ (.A(_1188_),
    .B(_1189_),
    .C(_0494_),
    .Y(_1262_));
 sky130_fd_sc_hd__nand3_1 _5325_ (.A(_1261_),
    .B(_1262_),
    .C(_0817_),
    .Y(_1263_));
 sky130_fd_sc_hd__nand3_1 _5326_ (.A(_1191_),
    .B(_1192_),
    .C(_0491_),
    .Y(_1264_));
 sky130_fd_sc_hd__nand3_1 _5327_ (.A(_1263_),
    .B(_1264_),
    .C(_1046_),
    .Y(_1265_));
 sky130_fd_sc_hd__nand3_1 _5328_ (.A(_1193_),
    .B(_1194_),
    .C(_0544_),
    .Y(_1266_));
 sky130_fd_sc_hd__nand3_1 _5329_ (.A(_1265_),
    .B(_1266_),
    .C(_0821_),
    .Y(_1268_));
 sky130_fd_sc_hd__nand3_1 _5330_ (.A(_1195_),
    .B(_1196_),
    .C(_0891_),
    .Y(_1269_));
 sky130_fd_sc_hd__nand3_1 _5331_ (.A(_1268_),
    .B(_1269_),
    .C(_1199_),
    .Y(_1270_));
 sky130_fd_sc_hd__nand3_1 _5332_ (.A(_1197_),
    .B(_1198_),
    .C(_0714_),
    .Y(_1271_));
 sky130_fd_sc_hd__nand3_1 _5333_ (.A(_1270_),
    .B(_1271_),
    .C(_0944_),
    .Y(_1272_));
 sky130_fd_sc_hd__nand3_1 _5334_ (.A(_1200_),
    .B(_1202_),
    .C(_0712_),
    .Y(_1273_));
 sky130_fd_sc_hd__nand3_1 _5335_ (.A(_1272_),
    .B(_1273_),
    .C(_0925_),
    .Y(_1274_));
 sky130_fd_sc_hd__nand3_1 _5336_ (.A(_1203_),
    .B(_1204_),
    .C(_0766_),
    .Y(_1275_));
 sky130_fd_sc_hd__nand3_1 _5337_ (.A(_1274_),
    .B(_1275_),
    .C(_0906_),
    .Y(_1276_));
 sky130_fd_sc_hd__nand3_1 _5338_ (.A(_1205_),
    .B(_1206_),
    .C(_0991_),
    .Y(_1277_));
 sky130_fd_sc_hd__nand3_1 _5339_ (.A(_1276_),
    .B(_1062_),
    .C(_1277_),
    .Y(_1279_));
 sky130_fd_sc_hd__nand3_1 _5340_ (.A(_1207_),
    .B(_1208_),
    .C(_0927_),
    .Y(_1280_));
 sky130_fd_sc_hd__nand3_1 _5341_ (.A(_0989_),
    .B(_1279_),
    .C(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__nand3_1 _5342_ (.A(_1081_),
    .B(_1240_),
    .C(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__nand2_1 _5343_ (.A(_1239_),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__nand2_1 _5344_ (.A(_1283_),
    .B(_1219_),
    .Y(_1284_));
 sky130_fd_sc_hd__nand2_1 _5345_ (.A(_1209_),
    .B(_1210_),
    .Y(_1285_));
 sky130_fd_sc_hd__nand3_1 _5346_ (.A(_1096_),
    .B(_1010_),
    .C(_1137_),
    .Y(_1286_));
 sky130_fd_sc_hd__o21ai_1 _5347_ (.A1(_1010_),
    .A2(_1285_),
    .B1(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__nand2_1 _5348_ (.A(_1287_),
    .B(_1081_),
    .Y(_1288_));
 sky130_fd_sc_hd__a21o_1 _5349_ (.A1(_1138_),
    .A2(_0989_),
    .B1(_1144_),
    .X(_1290_));
 sky130_fd_sc_hd__nand3_1 _5350_ (.A(_1288_),
    .B(_1290_),
    .C(_1218_),
    .Y(_1291_));
 sky130_fd_sc_hd__nand2_1 _5351_ (.A(_1284_),
    .B(_1291_),
    .Y(_1292_));
 sky130_fd_sc_hd__nand3_4 _5352_ (.A(_1147_),
    .B(_1213_),
    .C(_1081_),
    .Y(_1293_));
 sky130_fd_sc_hd__inv_4 _5353_ (.A(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__nand3_2 _5354_ (.A(_1238_),
    .B(_1292_),
    .C(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__inv_2 _5355_ (.A(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__nand3_1 _5356_ (.A(_1165_),
    .B(_1220_),
    .C(_1166_),
    .Y(_1297_));
 sky130_fd_sc_hd__nand3_2 _5357_ (.A(_1296_),
    .B(_1222_),
    .C(_1297_),
    .Y(_1298_));
 sky130_fd_sc_hd__inv_2 _5358_ (.A(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand3_4 _5359_ (.A(_1236_),
    .B(_1299_),
    .C(_1225_),
    .Y(_1301_));
 sky130_fd_sc_hd__inv_2 _5360_ (.A(_1301_),
    .Y(_1302_));
 sky130_fd_sc_hd__nand2_1 _5361_ (.A(_1230_),
    .B(_1225_),
    .Y(_1303_));
 sky130_fd_sc_hd__nand3_2 _5362_ (.A(_1302_),
    .B(_1228_),
    .C(_1303_),
    .Y(_1304_));
 sky130_fd_sc_hd__nand2_1 _5363_ (.A(_1233_),
    .B(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__nand2_1 _5364_ (.A(_1228_),
    .B(_1303_),
    .Y(_1306_));
 sky130_fd_sc_hd__nor2_1 _5365_ (.A(_1301_),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__nand3_2 _5366_ (.A(_1307_),
    .B(_1229_),
    .C(_1232_),
    .Y(_1308_));
 sky130_fd_sc_hd__nand2_1 _5367_ (.A(_1305_),
    .B(_1308_),
    .Y(_1309_));
 sky130_fd_sc_hd__nand2_1 _5368_ (.A(_1236_),
    .B(_1225_),
    .Y(_1310_));
 sky130_fd_sc_hd__nand2_1 _5369_ (.A(_1310_),
    .B(_1298_),
    .Y(_1312_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_1283_),
    .B(_1218_),
    .Y(_1313_));
 sky130_fd_sc_hd__a21o_1 _5371_ (.A1(_1263_),
    .A2(_1264_),
    .B1(_1046_),
    .X(_1314_));
 sky130_fd_sc_hd__mux2_1 _5372_ (.A0(_1244_),
    .A1(net140),
    .S(_0783_),
    .X(_1315_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net150),
    .A1(_1315_),
    .S(_2726_),
    .X(_1316_));
 sky130_fd_sc_hd__mux2_1 _5374_ (.A0(net151),
    .A1(_1247_),
    .S(_2733_),
    .X(_1317_));
 sky130_fd_sc_hd__or2_1 _5375_ (.A(_0198_),
    .B(_1317_),
    .X(_1318_));
 sky130_fd_sc_hd__or2_1 _5376_ (.A(_0788_),
    .B(_1248_),
    .X(_1319_));
 sky130_fd_sc_hd__nand2_1 _5377_ (.A(_1318_),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__nand2_1 _5378_ (.A(_1320_),
    .B(_0960_),
    .Y(_1321_));
 sky130_fd_sc_hd__nand2_1 _5379_ (.A(_1250_),
    .B(_0184_),
    .Y(_1323_));
 sky130_fd_sc_hd__nand2_1 _5380_ (.A(_1321_),
    .B(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__inv_2 _5381_ (.A(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_1 _5382_ (.A(_1325_),
    .B(_0676_),
    .Y(_1326_));
 sky130_fd_sc_hd__o21ai_1 _5383_ (.A1(_0676_),
    .A2(_1253_),
    .B1(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__nand2_1 _5384_ (.A(_1327_),
    .B(_0806_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2_1 _5385_ (.A(_1257_),
    .B(_0857_),
    .Y(_1329_));
 sky130_fd_sc_hd__nand2_1 _5386_ (.A(_1328_),
    .B(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__nand2_1 _5387_ (.A(_1330_),
    .B(_0429_),
    .Y(_1331_));
 sky130_fd_sc_hd__nand2_1 _5388_ (.A(_1243_),
    .B(_1258_),
    .Y(_1332_));
 sky130_fd_sc_hd__nand2_1 _5389_ (.A(_1332_),
    .B(_0878_),
    .Y(_1334_));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(_1331_),
    .B(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__nand2_1 _5391_ (.A(_1335_),
    .B(_0811_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand3_1 _5392_ (.A(_1242_),
    .B(_0881_),
    .C(_1259_),
    .Y(_1337_));
 sky130_fd_sc_hd__nand2_1 _5393_ (.A(_1336_),
    .B(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__nand2_1 _5394_ (.A(_1338_),
    .B(_1041_),
    .Y(_1339_));
 sky130_fd_sc_hd__nand2_1 _5395_ (.A(_1241_),
    .B(_1260_),
    .Y(_1340_));
 sky130_fd_sc_hd__nand2_1 _5396_ (.A(_1340_),
    .B(_0494_),
    .Y(_1341_));
 sky130_fd_sc_hd__nand2_1 _5397_ (.A(_1339_),
    .B(_1341_),
    .Y(_1342_));
 sky130_fd_sc_hd__nand2_1 _5398_ (.A(_1342_),
    .B(_0817_),
    .Y(_1343_));
 sky130_fd_sc_hd__nand3_1 _5399_ (.A(_1261_),
    .B(_1262_),
    .C(_0491_),
    .Y(_1345_));
 sky130_fd_sc_hd__nand2_1 _5400_ (.A(_1343_),
    .B(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__nand2_1 _5401_ (.A(_1346_),
    .B(_1046_),
    .Y(_1347_));
 sky130_fd_sc_hd__nand2_1 _5402_ (.A(_1314_),
    .B(_1347_),
    .Y(_1348_));
 sky130_fd_sc_hd__nand2_1 _5403_ (.A(_1348_),
    .B(_0821_),
    .Y(_1349_));
 sky130_fd_sc_hd__nand3_1 _5404_ (.A(_1265_),
    .B(_1266_),
    .C(_0891_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand3_1 _5405_ (.A(_1349_),
    .B(_1199_),
    .C(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__nand2_1 _5406_ (.A(_1268_),
    .B(_1269_),
    .Y(_1352_));
 sky130_fd_sc_hd__or2_1 _5407_ (.A(_1199_),
    .B(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__nand3_1 _5408_ (.A(_1351_),
    .B(_1353_),
    .C(_0944_),
    .Y(_1354_));
 sky130_fd_sc_hd__nand3_1 _5409_ (.A(_1270_),
    .B(_1271_),
    .C(_0712_),
    .Y(_1356_));
 sky130_fd_sc_hd__nand3_1 _5410_ (.A(_1354_),
    .B(_0925_),
    .C(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__nand2_1 _5411_ (.A(_1272_),
    .B(_1273_),
    .Y(_1358_));
 sky130_fd_sc_hd__or2_1 _5412_ (.A(_0925_),
    .B(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__nand3_1 _5413_ (.A(_1357_),
    .B(_1359_),
    .C(_0906_),
    .Y(_1360_));
 sky130_fd_sc_hd__nand3_1 _5414_ (.A(_1274_),
    .B(_1275_),
    .C(_0991_),
    .Y(_1361_));
 sky130_fd_sc_hd__nand3_1 _5415_ (.A(_1360_),
    .B(_1062_),
    .C(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__nand3_1 _5416_ (.A(_1276_),
    .B(_1277_),
    .C(_0927_),
    .Y(_1363_));
 sky130_fd_sc_hd__nand3_1 _5417_ (.A(_1362_),
    .B(_0989_),
    .C(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__nand3_1 _5418_ (.A(_1279_),
    .B(_1280_),
    .C(_1010_),
    .Y(_1365_));
 sky130_fd_sc_hd__nand3_1 _5419_ (.A(_1364_),
    .B(_1081_),
    .C(_1365_),
    .Y(_1367_));
 sky130_fd_sc_hd__nand3_1 _5420_ (.A(_1063_),
    .B(_1281_),
    .C(_1240_),
    .Y(_1368_));
 sky130_fd_sc_hd__nand2_1 _5421_ (.A(_1367_),
    .B(_1368_),
    .Y(_1369_));
 sky130_fd_sc_hd__nand2_1 _5422_ (.A(_1369_),
    .B(_1219_),
    .Y(_1370_));
 sky130_fd_sc_hd__nand2_1 _5423_ (.A(_1313_),
    .B(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__nand2_1 _5424_ (.A(_1371_),
    .B(_1294_),
    .Y(_1372_));
 sky130_fd_sc_hd__a21o_1 _5425_ (.A1(_1213_),
    .A2(_1081_),
    .B1(_1147_),
    .X(_1373_));
 sky130_fd_sc_hd__nand3_1 _5426_ (.A(_1239_),
    .B(_1219_),
    .C(_1282_),
    .Y(_1374_));
 sky130_fd_sc_hd__nand3_1 _5427_ (.A(_1373_),
    .B(_1374_),
    .C(_1293_),
    .Y(_1375_));
 sky130_fd_sc_hd__nand2_1 _5428_ (.A(_1372_),
    .B(_1375_),
    .Y(_1376_));
 sky130_fd_sc_hd__nand2_1 _5429_ (.A(_1238_),
    .B(_1293_),
    .Y(_1378_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(_1378_),
    .B(_1220_),
    .Y(_1379_));
 sky130_fd_sc_hd__nand2_1 _5431_ (.A(_1292_),
    .B(_1294_),
    .Y(_1380_));
 sky130_fd_sc_hd__inv_2 _5432_ (.A(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__nand3_1 _5433_ (.A(_1376_),
    .B(_1379_),
    .C(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__inv_2 _5434_ (.A(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__nand2_1 _5435_ (.A(_1222_),
    .B(_1297_),
    .Y(_1384_));
 sky130_fd_sc_hd__nand2_1 _5436_ (.A(_1384_),
    .B(_1295_),
    .Y(_1385_));
 sky130_fd_sc_hd__nand3_2 _5437_ (.A(_1383_),
    .B(_1298_),
    .C(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__inv_2 _5438_ (.A(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__nand3_4 _5439_ (.A(_1312_),
    .B(_1387_),
    .C(_1301_),
    .Y(_1389_));
 sky130_fd_sc_hd__inv_2 _5440_ (.A(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(_1306_),
    .B(_1301_),
    .Y(_1391_));
 sky130_fd_sc_hd__nand3_1 _5442_ (.A(_1390_),
    .B(_1391_),
    .C(_1304_),
    .Y(_1392_));
 sky130_fd_sc_hd__nand2_1 _5443_ (.A(_1309_),
    .B(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__nand2_1 _5444_ (.A(_1391_),
    .B(_1304_),
    .Y(_1394_));
 sky130_fd_sc_hd__nor2_1 _5445_ (.A(_1389_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__nand3_2 _5446_ (.A(_1395_),
    .B(_1305_),
    .C(_1308_),
    .Y(_1396_));
 sky130_fd_sc_hd__nand2_1 _5447_ (.A(_1393_),
    .B(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(_1394_),
    .B(_1390_),
    .Y(_1398_));
 sky130_fd_sc_hd__nand3_1 _5449_ (.A(_1391_),
    .B(_1304_),
    .C(_1389_),
    .Y(_1400_));
 sky130_fd_sc_hd__nand2_1 _5450_ (.A(_1398_),
    .B(_1400_),
    .Y(_1401_));
 sky130_fd_sc_hd__or2_1 _5451_ (.A(_1294_),
    .B(_1371_),
    .X(_1402_));
 sky130_fd_sc_hd__nand2_1 _5452_ (.A(_1327_),
    .B(_0857_),
    .Y(_1403_));
 sky130_fd_sc_hd__mux2_1 _5453_ (.A0(_1315_),
    .A1(net141),
    .S(_2726_),
    .X(_1404_));
 sky130_fd_sc_hd__mux2_1 _5454_ (.A0(net151),
    .A1(_1404_),
    .S(_0609_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2_1 _5455_ (.A0(_1317_),
    .A1(net152),
    .S(_0788_),
    .X(_1406_));
 sky130_fd_sc_hd__nand2_1 _5456_ (.A(_1406_),
    .B(_0960_),
    .Y(_1407_));
 sky130_fd_sc_hd__o21ai_1 _5457_ (.A1(_0960_),
    .A2(_1320_),
    .B1(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__nand2_1 _5458_ (.A(_1408_),
    .B(_0676_),
    .Y(_1409_));
 sky130_fd_sc_hd__nand2_1 _5459_ (.A(_1325_),
    .B(_0874_),
    .Y(_1411_));
 sky130_fd_sc_hd__nand2_1 _5460_ (.A(_1409_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__nand2_1 _5461_ (.A(_1412_),
    .B(_0806_),
    .Y(_1413_));
 sky130_fd_sc_hd__nand2_1 _5462_ (.A(_1403_),
    .B(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(_1414_),
    .A1(_1330_),
    .S(_0878_),
    .X(_1415_));
 sky130_fd_sc_hd__nand2_1 _5464_ (.A(_1415_),
    .B(_0811_),
    .Y(_1416_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(_1335_),
    .B(_0881_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _5466_ (.A(_1416_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__nand2_1 _5467_ (.A(_1418_),
    .B(_1041_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_1 _5468_ (.A(_1338_),
    .B(_0494_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _5469_ (.A(_1419_),
    .B(_1420_),
    .Y(_1422_));
 sky130_fd_sc_hd__nand2_1 _5470_ (.A(_1422_),
    .B(_0817_),
    .Y(_1423_));
 sky130_fd_sc_hd__nand2_1 _5471_ (.A(_1342_),
    .B(_0491_),
    .Y(_1424_));
 sky130_fd_sc_hd__nand2_1 _5472_ (.A(_1423_),
    .B(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__nand2_1 _5473_ (.A(_1425_),
    .B(_1046_),
    .Y(_1426_));
 sky130_fd_sc_hd__nand2_1 _5474_ (.A(_1346_),
    .B(_0544_),
    .Y(_1427_));
 sky130_fd_sc_hd__nand2_1 _5475_ (.A(_1426_),
    .B(_1427_),
    .Y(_1428_));
 sky130_fd_sc_hd__nand2_1 _5476_ (.A(_1428_),
    .B(_0821_),
    .Y(_1429_));
 sky130_fd_sc_hd__nand2_1 _5477_ (.A(_1348_),
    .B(_0891_),
    .Y(_1430_));
 sky130_fd_sc_hd__nand2_1 _5478_ (.A(_1429_),
    .B(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__nand2_1 _5479_ (.A(_1431_),
    .B(_1199_),
    .Y(_1433_));
 sky130_fd_sc_hd__nand2_1 _5480_ (.A(_1349_),
    .B(_1350_),
    .Y(_1434_));
 sky130_fd_sc_hd__nand2_1 _5481_ (.A(_1434_),
    .B(_0714_),
    .Y(_1435_));
 sky130_fd_sc_hd__nand3_1 _5482_ (.A(_1433_),
    .B(_1435_),
    .C(_0944_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_1434_),
    .B(_1199_),
    .Y(_1437_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_1352_),
    .B(_0714_),
    .Y(_1438_));
 sky130_fd_sc_hd__nand2_1 _5485_ (.A(_1437_),
    .B(_1438_),
    .Y(_1439_));
 sky130_fd_sc_hd__or2_1 _5486_ (.A(_0944_),
    .B(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__nand3_1 _5487_ (.A(_1436_),
    .B(_1440_),
    .C(_0925_),
    .Y(_1441_));
 sky130_fd_sc_hd__a21o_1 _5488_ (.A1(_1354_),
    .A2(_1356_),
    .B1(_0925_),
    .X(_1442_));
 sky130_fd_sc_hd__nand3_1 _5489_ (.A(_1441_),
    .B(_1442_),
    .C(_0906_),
    .Y(_1444_));
 sky130_fd_sc_hd__a21o_1 _5490_ (.A1(_1357_),
    .A2(_1359_),
    .B1(_0906_),
    .X(_1445_));
 sky130_fd_sc_hd__nand3_1 _5491_ (.A(_1444_),
    .B(_1445_),
    .C(_1062_),
    .Y(_1446_));
 sky130_fd_sc_hd__a21o_1 _5492_ (.A1(_1360_),
    .A2(_1361_),
    .B1(_1062_),
    .X(_1447_));
 sky130_fd_sc_hd__nand3_1 _5493_ (.A(_1446_),
    .B(_1447_),
    .C(_0989_),
    .Y(_1448_));
 sky130_fd_sc_hd__nand2_1 _5494_ (.A(_1362_),
    .B(_1363_),
    .Y(_1449_));
 sky130_fd_sc_hd__nand2_1 _5495_ (.A(_1449_),
    .B(_1010_),
    .Y(_1450_));
 sky130_fd_sc_hd__nand3_1 _5496_ (.A(_1448_),
    .B(_1450_),
    .C(_1081_),
    .Y(_1451_));
 sky130_fd_sc_hd__a21o_1 _5497_ (.A1(_1364_),
    .A2(_1365_),
    .B1(_1081_),
    .X(_1452_));
 sky130_fd_sc_hd__nand3_1 _5498_ (.A(_1451_),
    .B(_1219_),
    .C(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__nand2_1 _5499_ (.A(_1369_),
    .B(_1218_),
    .Y(_1455_));
 sky130_fd_sc_hd__nand3_1 _5500_ (.A(_1453_),
    .B(_1455_),
    .C(_1294_),
    .Y(_1456_));
 sky130_fd_sc_hd__nand3_1 _5501_ (.A(_1402_),
    .B(_1456_),
    .C(_1381_),
    .Y(_1457_));
 sky130_fd_sc_hd__nand2_1 _5502_ (.A(_1376_),
    .B(_1380_),
    .Y(_1458_));
 sky130_fd_sc_hd__nand2_1 _5503_ (.A(_1457_),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__nand2_1 _5504_ (.A(_1376_),
    .B(_1381_),
    .Y(_1460_));
 sky130_fd_sc_hd__inv_2 _5505_ (.A(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__nand2_1 _5506_ (.A(_1459_),
    .B(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__inv_2 _5507_ (.A(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__a21o_1 _5508_ (.A1(_1298_),
    .A2(_1385_),
    .B1(_1383_),
    .X(_1464_));
 sky130_fd_sc_hd__nand2_1 _5509_ (.A(_1464_),
    .B(_1386_),
    .Y(_1466_));
 sky130_fd_sc_hd__inv_2 _5510_ (.A(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2_1 _5511_ (.A(_1379_),
    .B(_1380_),
    .Y(_1468_));
 sky130_fd_sc_hd__nand2_1 _5512_ (.A(_1468_),
    .B(_1295_),
    .Y(_1469_));
 sky130_fd_sc_hd__nand2_1 _5513_ (.A(_1469_),
    .B(_1461_),
    .Y(_1470_));
 sky130_fd_sc_hd__nand3_1 _5514_ (.A(_1468_),
    .B(_1460_),
    .C(_1295_),
    .Y(_1471_));
 sky130_fd_sc_hd__and2_1 _5515_ (.A(_1470_),
    .B(_1471_),
    .X(_1472_));
 sky130_fd_sc_hd__inv_2 _5516_ (.A(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__nand2_1 _5517_ (.A(_1467_),
    .B(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _5518_ (.A(_1312_),
    .B(_1301_),
    .Y(_1475_));
 sky130_fd_sc_hd__nand2_1 _5519_ (.A(_1475_),
    .B(_1386_),
    .Y(_1477_));
 sky130_fd_sc_hd__nand2_1 _5520_ (.A(_1477_),
    .B(_1389_),
    .Y(_1478_));
 sky130_fd_sc_hd__nor2_1 _5521_ (.A(_1474_),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__nand3_1 _5522_ (.A(_1401_),
    .B(_1463_),
    .C(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(_1397_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__nand3_1 _5524_ (.A(_1459_),
    .B(_1461_),
    .C(_1469_),
    .Y(_1482_));
 sky130_fd_sc_hd__inv_2 _5525_ (.A(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__nand3_2 _5526_ (.A(_1483_),
    .B(_1464_),
    .C(_1386_),
    .Y(_1484_));
 sky130_fd_sc_hd__inv_2 _5527_ (.A(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__nand3_2 _5528_ (.A(_1485_),
    .B(_1389_),
    .C(_1477_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand2_1 _5529_ (.A(_1394_),
    .B(_1389_),
    .Y(_1488_));
 sky130_fd_sc_hd__nand2_1 _5530_ (.A(_1488_),
    .B(_1392_),
    .Y(_1489_));
 sky130_fd_sc_hd__nor2_1 _5531_ (.A(_1486_),
    .B(_1489_),
    .Y(_1490_));
 sky130_fd_sc_hd__nand3_2 _5532_ (.A(_1490_),
    .B(_1393_),
    .C(_1396_),
    .Y(_1491_));
 sky130_fd_sc_hd__nand2_1 _5533_ (.A(_1481_),
    .B(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_1 _5534_ (.A(_1472_),
    .B(_1462_),
    .Y(_1493_));
 sky130_fd_sc_hd__nand3_1 _5535_ (.A(_1467_),
    .B(_1493_),
    .C(_1482_),
    .Y(_1494_));
 sky130_fd_sc_hd__nand2_1 _5536_ (.A(_1478_),
    .B(_1484_),
    .Y(_1495_));
 sky130_fd_sc_hd__nand3_1 _5537_ (.A(_1401_),
    .B(_1486_),
    .C(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__nor2_1 _5538_ (.A(_1494_),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__inv_2 _5539_ (.A(_1497_),
    .Y(_1499_));
 sky130_fd_sc_hd__nand2_1 _5540_ (.A(_1492_),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__nand3_1 _5541_ (.A(_1481_),
    .B(_1491_),
    .C(_1497_),
    .Y(_1501_));
 sky130_fd_sc_hd__nand2_1 _5542_ (.A(_1500_),
    .B(_1501_),
    .Y(_1502_));
 sky130_fd_sc_hd__and2_1 _5543_ (.A(_1436_),
    .B(_1440_),
    .X(_1503_));
 sky130_fd_sc_hd__inv_2 _5544_ (.A(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__mux2_1 _5545_ (.A0(_1404_),
    .A1(net142),
    .S(_0609_),
    .X(_1505_));
 sky130_fd_sc_hd__mux2_1 _5546_ (.A0(net152),
    .A1(_1505_),
    .S(_0788_),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(_1406_),
    .A1(_1506_),
    .S(_0960_),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _5548_ (.A0(_1507_),
    .A1(_1408_),
    .S(_0874_),
    .X(_1508_));
 sky130_fd_sc_hd__nand2_1 _5549_ (.A(_1508_),
    .B(_0806_),
    .Y(_1510_));
 sky130_fd_sc_hd__nand2_1 _5550_ (.A(_1412_),
    .B(_0857_),
    .Y(_1511_));
 sky130_fd_sc_hd__nand2_1 _5551_ (.A(_1510_),
    .B(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__or2_1 _5552_ (.A(_0878_),
    .B(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__or2_1 _5553_ (.A(_0429_),
    .B(_1414_),
    .X(_1514_));
 sky130_fd_sc_hd__nand2_1 _5554_ (.A(_1513_),
    .B(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__or2_1 _5555_ (.A(_0881_),
    .B(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__nand2_1 _5556_ (.A(_1415_),
    .B(_0881_),
    .Y(_1517_));
 sky130_fd_sc_hd__nand3_1 _5557_ (.A(_1516_),
    .B(_1041_),
    .C(_1517_),
    .Y(_1518_));
 sky130_fd_sc_hd__or2_1 _5558_ (.A(_1041_),
    .B(_1418_),
    .X(_1519_));
 sky130_fd_sc_hd__nand3_1 _5559_ (.A(_1518_),
    .B(_0817_),
    .C(_1519_),
    .Y(_1521_));
 sky130_fd_sc_hd__nand2_1 _5560_ (.A(_1422_),
    .B(_0491_),
    .Y(_1522_));
 sky130_fd_sc_hd__nand3_1 _5561_ (.A(_1521_),
    .B(_1046_),
    .C(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__or2_1 _5562_ (.A(_1046_),
    .B(_1425_),
    .X(_1524_));
 sky130_fd_sc_hd__nand3_1 _5563_ (.A(_1523_),
    .B(_0821_),
    .C(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__nand2_1 _5564_ (.A(_1428_),
    .B(_0891_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand3_1 _5565_ (.A(_1525_),
    .B(_1199_),
    .C(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__or2_1 _5566_ (.A(_1199_),
    .B(_1431_),
    .X(_1528_));
 sky130_fd_sc_hd__nand3_1 _5567_ (.A(_1527_),
    .B(_0944_),
    .C(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__a21o_1 _5568_ (.A1(_1433_),
    .A2(_1435_),
    .B1(_0944_),
    .X(_1530_));
 sky130_fd_sc_hd__nand2_1 _5569_ (.A(_1529_),
    .B(_1530_),
    .Y(_1532_));
 sky130_fd_sc_hd__nand2_1 _5570_ (.A(_1532_),
    .B(_0925_),
    .Y(_1533_));
 sky130_fd_sc_hd__o211ai_1 _5571_ (.A1(_0925_),
    .A2(_1504_),
    .B1(_0906_),
    .C1(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__nand3_1 _5572_ (.A(_1441_),
    .B(_0991_),
    .C(_1442_),
    .Y(_1535_));
 sky130_fd_sc_hd__nand3_1 _5573_ (.A(_1534_),
    .B(_1062_),
    .C(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__and2_1 _5574_ (.A(_1444_),
    .B(_1445_),
    .X(_1537_));
 sky130_fd_sc_hd__nand2_1 _5575_ (.A(_1537_),
    .B(_0927_),
    .Y(_1538_));
 sky130_fd_sc_hd__nand3_1 _5576_ (.A(_1536_),
    .B(_0989_),
    .C(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__nand3_1 _5577_ (.A(_1446_),
    .B(_1010_),
    .C(_1447_),
    .Y(_1540_));
 sky130_fd_sc_hd__nand3_1 _5578_ (.A(_1539_),
    .B(_1081_),
    .C(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__nand3_1 _5579_ (.A(_1448_),
    .B(_1063_),
    .C(_1450_),
    .Y(_1543_));
 sky130_fd_sc_hd__nand3_1 _5580_ (.A(_1541_),
    .B(_1219_),
    .C(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__nand3_1 _5581_ (.A(_1451_),
    .B(_1218_),
    .C(_1452_),
    .Y(_1545_));
 sky130_fd_sc_hd__nand3_1 _5582_ (.A(_1544_),
    .B(_1294_),
    .C(_1545_),
    .Y(_1546_));
 sky130_fd_sc_hd__nand3_1 _5583_ (.A(_1453_),
    .B(_1293_),
    .C(_1455_),
    .Y(_1547_));
 sky130_fd_sc_hd__nand2_1 _5584_ (.A(_1546_),
    .B(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__a21oi_1 _5585_ (.A1(_1402_),
    .A2(_1456_),
    .B1(_1381_),
    .Y(_1549_));
 sky130_fd_sc_hd__a21oi_2 _5586_ (.A1(_1548_),
    .A2(_1381_),
    .B1(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__nand2_4 _5587_ (.A(_1550_),
    .B(_1463_),
    .Y(_1551_));
 sky130_fd_sc_hd__inv_2 _5588_ (.A(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__nand2_1 _5589_ (.A(_1502_),
    .B(_1552_),
    .Y(_1554_));
 sky130_fd_sc_hd__nand2_1 _5590_ (.A(_1492_),
    .B(_1551_),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_1 _5591_ (.A(_1554_),
    .B(_1555_),
    .Y(_1556_));
 sky130_fd_sc_hd__nand2_1 _5592_ (.A(_1489_),
    .B(_1486_),
    .Y(_1557_));
 sky130_fd_sc_hd__nand2_1 _5593_ (.A(_1480_),
    .B(_1557_),
    .Y(_1558_));
 sky130_fd_sc_hd__nand2_1 _5594_ (.A(_1486_),
    .B(_1495_),
    .Y(_1559_));
 sky130_fd_sc_hd__nor2_1 _5595_ (.A(_1551_),
    .B(_1494_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2b_1 _5596_ (.A_N(_1559_),
    .B(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__inv_2 _5597_ (.A(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__nor2_1 _5598_ (.A(_1558_),
    .B(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__inv_2 _5599_ (.A(_1563_),
    .Y(_1565_));
 sky130_fd_sc_hd__inv_2 _5600_ (.A(_1560_),
    .Y(_1566_));
 sky130_fd_sc_hd__nand2_1 _5601_ (.A(_1566_),
    .B(_1559_),
    .Y(_1567_));
 sky130_fd_sc_hd__nand2_1 _5602_ (.A(_1473_),
    .B(_1462_),
    .Y(_1568_));
 sky130_fd_sc_hd__nand2_1 _5603_ (.A(_1472_),
    .B(_1463_),
    .Y(_1569_));
 sky130_fd_sc_hd__nand2_1 _5604_ (.A(_1568_),
    .B(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__nand2_1 _5605_ (.A(_1552_),
    .B(_1570_),
    .Y(_1571_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_1466_),
    .B(_1482_),
    .Y(_1572_));
 sky130_fd_sc_hd__nand2_1 _5607_ (.A(_1572_),
    .B(_1484_),
    .Y(_1573_));
 sky130_fd_sc_hd__nand2_1 _5608_ (.A(_1571_),
    .B(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__nand2_1 _5609_ (.A(_1566_),
    .B(_1574_),
    .Y(_1576_));
 sky130_fd_sc_hd__inv_2 _5610_ (.A(_1570_),
    .Y(_1577_));
 sky130_fd_sc_hd__nand2_1 _5611_ (.A(_1577_),
    .B(_1551_),
    .Y(_1578_));
 sky130_fd_sc_hd__nand2_1 _5612_ (.A(_1571_),
    .B(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__nand2_1 _5613_ (.A(_1576_),
    .B(_1579_),
    .Y(_1580_));
 sky130_fd_sc_hd__a21oi_1 _5614_ (.A1(_1561_),
    .A2(_1567_),
    .B1(_1580_),
    .Y(_1581_));
 sky130_fd_sc_hd__nand2_1 _5615_ (.A(_1562_),
    .B(_1558_),
    .Y(_1582_));
 sky130_fd_sc_hd__nand3_1 _5616_ (.A(_1565_),
    .B(_1581_),
    .C(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__inv_2 _5617_ (.A(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__nand2_1 _5618_ (.A(_1556_),
    .B(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__nand3_1 _5619_ (.A(_1554_),
    .B(_1555_),
    .C(_1583_),
    .Y(_1587_));
 sky130_fd_sc_hd__nand3_1 _5620_ (.A(_1585_),
    .B(_1551_),
    .C(_1587_),
    .Y(_1588_));
 sky130_fd_sc_hd__nand2_1 _5621_ (.A(_1588_),
    .B(_1554_),
    .Y(_1589_));
 sky130_fd_sc_hd__nand2_1 _5622_ (.A(_1491_),
    .B(_1396_),
    .Y(_1590_));
 sky130_fd_sc_hd__nor2_1 _5623_ (.A(_1228_),
    .B(_1158_),
    .Y(_1591_));
 sky130_fd_sc_hd__nand2_1 _5624_ (.A(_0850_),
    .B(_0778_),
    .Y(_1592_));
 sky130_fd_sc_hd__nor2_1 _5625_ (.A(_0486_),
    .B(_0443_),
    .Y(_1593_));
 sky130_fd_sc_hd__nor2_1 _5626_ (.A(_0437_),
    .B(_0395_),
    .Y(_1594_));
 sky130_fd_sc_hd__nor2_1 _5627_ (.A(_0390_),
    .B(_0355_),
    .Y(_1595_));
 sky130_fd_sc_hd__nor2_1 _5628_ (.A(_0353_),
    .B(_0350_),
    .Y(_1596_));
 sky130_fd_sc_hd__nand2_1 _5629_ (.A(_1674_),
    .B(net21),
    .Y(_1598_));
 sky130_fd_sc_hd__o21ai_2 _5630_ (.A1(_1300_),
    .A2(_1674_),
    .B1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__inv_2 _5631_ (.A(_1599_),
    .Y(_1600_));
 sky130_fd_sc_hd__nand2_1 _5632_ (.A(_0317_),
    .B(_1600_),
    .Y(_1601_));
 sky130_fd_sc_hd__nand3_1 _5633_ (.A(_0162_),
    .B(_1599_),
    .C(_0316_),
    .Y(_1602_));
 sky130_fd_sc_hd__nand2_1 _5634_ (.A(_1601_),
    .B(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__inv_2 _5635_ (.A(_1603_),
    .Y(_1604_));
 sky130_fd_sc_hd__nand2_1 _5636_ (.A(_0322_),
    .B(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__nand3_1 _5637_ (.A(_0320_),
    .B(_1603_),
    .C(_0321_),
    .Y(_1606_));
 sky130_fd_sc_hd__nand2_1 _5638_ (.A(_1605_),
    .B(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_0326_),
    .B(_1607_),
    .Y(_1609_));
 sky130_fd_sc_hd__nor2_1 _5640_ (.A(_0168_),
    .B(_0323_),
    .Y(_1610_));
 sky130_fd_sc_hd__inv_2 _5641_ (.A(_1607_),
    .Y(_1611_));
 sky130_fd_sc_hd__nand2_1 _5642_ (.A(_1610_),
    .B(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__nand2_1 _5643_ (.A(_1609_),
    .B(_1612_),
    .Y(_1613_));
 sky130_fd_sc_hd__inv_2 _5644_ (.A(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__nor2_1 _5645_ (.A(_0331_),
    .B(_0330_),
    .Y(_1615_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_1614_),
    .B(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__nand2_1 _5647_ (.A(_0328_),
    .B(_1613_),
    .Y(_1617_));
 sky130_fd_sc_hd__nand2_1 _5648_ (.A(_1616_),
    .B(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__xor2_1 _5649_ (.A(_0337_),
    .B(_1618_),
    .X(_1620_));
 sky130_fd_sc_hd__inv_2 _5650_ (.A(_0341_),
    .Y(_1621_));
 sky130_fd_sc_hd__nand2_1 _5651_ (.A(_1620_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__nor2_1 _5652_ (.A(_0229_),
    .B(_0343_),
    .Y(_1623_));
 sky130_fd_sc_hd__inv_2 _5653_ (.A(_0337_),
    .Y(_1624_));
 sky130_fd_sc_hd__nand3_1 _5654_ (.A(_1624_),
    .B(_1616_),
    .C(_1617_),
    .Y(_1625_));
 sky130_fd_sc_hd__nand2_1 _5655_ (.A(_1618_),
    .B(_0337_),
    .Y(_1626_));
 sky130_fd_sc_hd__nand2_1 _5656_ (.A(_1625_),
    .B(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__nand2_1 _5657_ (.A(_1627_),
    .B(_0341_),
    .Y(_1628_));
 sky130_fd_sc_hd__nand3_1 _5658_ (.A(_1622_),
    .B(_1623_),
    .C(_1628_),
    .Y(_1629_));
 sky130_fd_sc_hd__inv_2 _5659_ (.A(_0338_),
    .Y(_1631_));
 sky130_fd_sc_hd__inv_2 _5660_ (.A(_0189_),
    .Y(_1632_));
 sky130_fd_sc_hd__nand3_1 _5661_ (.A(_0176_),
    .B(_0191_),
    .C(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__nor2_1 _5662_ (.A(_1633_),
    .B(_0174_),
    .Y(_1634_));
 sky130_fd_sc_hd__nand3_1 _5663_ (.A(_1631_),
    .B(_0960_),
    .C(_1634_),
    .Y(_1635_));
 sky130_fd_sc_hd__nand2_1 _5664_ (.A(_1620_),
    .B(_1635_),
    .Y(_1636_));
 sky130_fd_sc_hd__nand2_1 _5665_ (.A(_1634_),
    .B(_0960_),
    .Y(_1637_));
 sky130_fd_sc_hd__nor2_1 _5666_ (.A(_0338_),
    .B(_1637_),
    .Y(_1638_));
 sky130_fd_sc_hd__nand2_1 _5667_ (.A(_1627_),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__nand3_1 _5668_ (.A(_1636_),
    .B(_1639_),
    .C(_0342_),
    .Y(_1640_));
 sky130_fd_sc_hd__nand2_1 _5669_ (.A(_1629_),
    .B(_1640_),
    .Y(_1642_));
 sky130_fd_sc_hd__nand2_1 _5670_ (.A(_1642_),
    .B(_0345_),
    .Y(_1643_));
 sky130_fd_sc_hd__nor2_1 _5671_ (.A(_0347_),
    .B(_0346_),
    .Y(_1644_));
 sky130_fd_sc_hd__nand3_2 _5672_ (.A(_1644_),
    .B(_1629_),
    .C(_1640_),
    .Y(_1645_));
 sky130_fd_sc_hd__nand3_2 _5673_ (.A(_1596_),
    .B(_1643_),
    .C(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__nand2_1 _5674_ (.A(_1643_),
    .B(_1645_),
    .Y(_1647_));
 sky130_fd_sc_hd__nand2_1 _5675_ (.A(_1647_),
    .B(_0349_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand3_2 _5676_ (.A(_1595_),
    .B(_1646_),
    .C(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__nand2_1 _5677_ (.A(_1648_),
    .B(_1646_),
    .Y(_1650_));
 sky130_fd_sc_hd__nand2_1 _5678_ (.A(_1650_),
    .B(_0394_),
    .Y(_1651_));
 sky130_fd_sc_hd__nand3_1 _5679_ (.A(_1594_),
    .B(_1649_),
    .C(_1651_),
    .Y(_1653_));
 sky130_fd_sc_hd__nand2_1 _5680_ (.A(_1649_),
    .B(_1651_),
    .Y(_1654_));
 sky130_fd_sc_hd__nand2_1 _5681_ (.A(_1654_),
    .B(_0442_),
    .Y(_1655_));
 sky130_fd_sc_hd__nand3_1 _5682_ (.A(_1593_),
    .B(_1653_),
    .C(_1655_),
    .Y(_1656_));
 sky130_fd_sc_hd__inv_2 _5683_ (.A(_0395_),
    .Y(_1657_));
 sky130_fd_sc_hd__nor2_1 _5684_ (.A(_0493_),
    .B(_0448_),
    .Y(_1658_));
 sky130_fd_sc_hd__nand3_1 _5685_ (.A(_0400_),
    .B(_0387_),
    .C(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__inv_2 _5686_ (.A(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__nand3_1 _5687_ (.A(_0398_),
    .B(_1041_),
    .C(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__inv_2 _5688_ (.A(_1661_),
    .Y(_1662_));
 sky130_fd_sc_hd__nand2_1 _5689_ (.A(_1657_),
    .B(_1662_),
    .Y(_1664_));
 sky130_fd_sc_hd__nand3_1 _5690_ (.A(_1664_),
    .B(_1649_),
    .C(_1651_),
    .Y(_1665_));
 sky130_fd_sc_hd__nor2_1 _5691_ (.A(_1661_),
    .B(_0395_),
    .Y(_1666_));
 sky130_fd_sc_hd__nand2_1 _5692_ (.A(_1654_),
    .B(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__nand3_1 _5693_ (.A(_1665_),
    .B(_1667_),
    .C(_0488_),
    .Y(_1668_));
 sky130_fd_sc_hd__nand2_1 _5694_ (.A(_1656_),
    .B(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__nand2_1 _5695_ (.A(_1669_),
    .B(_0538_),
    .Y(_1670_));
 sky130_fd_sc_hd__nor2_1 _5696_ (.A(_0536_),
    .B(_0489_),
    .Y(_1671_));
 sky130_fd_sc_hd__nand3_1 _5697_ (.A(_1671_),
    .B(_1656_),
    .C(_1668_),
    .Y(_1672_));
 sky130_fd_sc_hd__nand2_1 _5698_ (.A(_1670_),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__nand2_1 _5699_ (.A(_1673_),
    .B(_0593_),
    .Y(_1675_));
 sky130_fd_sc_hd__inv_2 _5700_ (.A(_0593_),
    .Y(_1676_));
 sky130_fd_sc_hd__nand3_1 _5701_ (.A(_1676_),
    .B(_1670_),
    .C(_1672_),
    .Y(_1677_));
 sky130_fd_sc_hd__nand2_1 _5702_ (.A(_1675_),
    .B(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__or2_1 _5703_ (.A(_0601_),
    .B(_0655_),
    .X(_1679_));
 sky130_fd_sc_hd__nand3b_1 _5704_ (.A_N(_1679_),
    .B(_0584_),
    .C(_0596_),
    .Y(_1680_));
 sky130_fd_sc_hd__nand3b_1 _5705_ (.A_N(_1680_),
    .B(_0646_),
    .C(_1199_),
    .Y(_1681_));
 sky130_fd_sc_hd__nor2_1 _5706_ (.A(_0594_),
    .B(_1681_),
    .Y(_1682_));
 sky130_fd_sc_hd__nand2_1 _5707_ (.A(_1678_),
    .B(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__nand3_1 _5708_ (.A(_1675_),
    .B(_1677_),
    .C(_0650_),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_1 _5709_ (.A(_1683_),
    .B(_1684_),
    .Y(_1686_));
 sky130_fd_sc_hd__inv_2 _5710_ (.A(_0707_),
    .Y(_1687_));
 sky130_fd_sc_hd__nand2_1 _5711_ (.A(_1686_),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__nand3_1 _5712_ (.A(_1683_),
    .B(_1684_),
    .C(_0707_),
    .Y(_1689_));
 sky130_fd_sc_hd__nand2_1 _5713_ (.A(_1688_),
    .B(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__nand2_1 _5714_ (.A(_1592_),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__inv_2 _5715_ (.A(_1690_),
    .Y(_1692_));
 sky130_fd_sc_hd__nand3_2 _5716_ (.A(_0850_),
    .B(_1692_),
    .C(_0778_),
    .Y(_1693_));
 sky130_fd_sc_hd__nand2_1 _5717_ (.A(_1691_),
    .B(_1693_),
    .Y(_1694_));
 sky130_fd_sc_hd__inv_2 _5718_ (.A(_0921_),
    .Y(_1695_));
 sky130_fd_sc_hd__nand2_1 _5719_ (.A(_1694_),
    .B(_1695_),
    .Y(_1697_));
 sky130_fd_sc_hd__nand3_1 _5720_ (.A(_1691_),
    .B(_0921_),
    .C(_1693_),
    .Y(_1698_));
 sky130_fd_sc_hd__nand2_1 _5721_ (.A(_1697_),
    .B(_1698_),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_1 _5722_ (.A(_1699_),
    .B(_1006_),
    .Y(_1700_));
 sky130_fd_sc_hd__nand3b_1 _5723_ (.A_N(_0922_),
    .B(_1694_),
    .C(_1005_),
    .Y(_1701_));
 sky130_fd_sc_hd__nand2_1 _5724_ (.A(_1700_),
    .B(_1701_),
    .Y(_1702_));
 sky130_fd_sc_hd__inv_2 _5725_ (.A(_1087_),
    .Y(_1703_));
 sky130_fd_sc_hd__nand3b_1 _5726_ (.A_N(_1702_),
    .B(_1703_),
    .C(_1155_),
    .Y(_1704_));
 sky130_fd_sc_hd__nand3_1 _5727_ (.A(_1074_),
    .B(_1001_),
    .C(_1006_),
    .Y(_1705_));
 sky130_fd_sc_hd__inv_2 _5728_ (.A(_1705_),
    .Y(_1706_));
 sky130_fd_sc_hd__nand2_1 _5729_ (.A(_1702_),
    .B(_1706_),
    .Y(_1708_));
 sky130_fd_sc_hd__nand3_1 _5730_ (.A(_1705_),
    .B(_1700_),
    .C(_1701_),
    .Y(_1709_));
 sky130_fd_sc_hd__nand3_1 _5731_ (.A(_1156_),
    .B(_1708_),
    .C(_1709_),
    .Y(_1710_));
 sky130_fd_sc_hd__nand3_1 _5732_ (.A(_1591_),
    .B(_1704_),
    .C(_1710_),
    .Y(_1711_));
 sky130_fd_sc_hd__nand2_1 _5733_ (.A(_1710_),
    .B(_1704_),
    .Y(_1712_));
 sky130_fd_sc_hd__nand2_1 _5734_ (.A(_1712_),
    .B(_1232_),
    .Y(_1713_));
 sky130_fd_sc_hd__nand2_1 _5735_ (.A(_1711_),
    .B(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__nand2_1 _5736_ (.A(_1714_),
    .B(_1308_),
    .Y(_1715_));
 sky130_fd_sc_hd__nor2_1 _5737_ (.A(_1712_),
    .B(_1308_),
    .Y(_1716_));
 sky130_fd_sc_hd__inv_2 _5738_ (.A(_1716_),
    .Y(_1717_));
 sky130_fd_sc_hd__nand2_1 _5739_ (.A(_1715_),
    .B(_1717_),
    .Y(_1719_));
 sky130_fd_sc_hd__inv_2 _5740_ (.A(_1719_),
    .Y(_1720_));
 sky130_fd_sc_hd__nand2_1 _5741_ (.A(_1590_),
    .B(_1720_),
    .Y(_1721_));
 sky130_fd_sc_hd__nand3_1 _5742_ (.A(_1491_),
    .B(_1719_),
    .C(_1396_),
    .Y(_1722_));
 sky130_fd_sc_hd__nand2_1 _5743_ (.A(_1721_),
    .B(_1722_),
    .Y(_1723_));
 sky130_fd_sc_hd__inv_2 _5744_ (.A(_1723_),
    .Y(_1724_));
 sky130_fd_sc_hd__inv_2 _5745_ (.A(_1492_),
    .Y(_1725_));
 sky130_fd_sc_hd__nand3_1 _5746_ (.A(_1725_),
    .B(_1552_),
    .C(_1497_),
    .Y(_1726_));
 sky130_fd_sc_hd__nand2_1 _5747_ (.A(_1724_),
    .B(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__nor2_1 _5748_ (.A(_1551_),
    .B(_1501_),
    .Y(_1728_));
 sky130_fd_sc_hd__nand2_1 _5749_ (.A(_1728_),
    .B(_1723_),
    .Y(_1730_));
 sky130_fd_sc_hd__nand2_1 _5750_ (.A(_1727_),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__nor2_1 _5751_ (.A(_1552_),
    .B(_1583_),
    .Y(_1732_));
 sky130_fd_sc_hd__nand3_1 _5752_ (.A(_1731_),
    .B(_1556_),
    .C(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__nand2_1 _5753_ (.A(_1556_),
    .B(_1732_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _5754_ (.A(_1724_),
    .B(_1728_),
    .Y(_1735_));
 sky130_fd_sc_hd__nand2_1 _5755_ (.A(_1726_),
    .B(_1723_),
    .Y(_1736_));
 sky130_fd_sc_hd__nand2_1 _5756_ (.A(_1735_),
    .B(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__nand2_1 _5757_ (.A(_1734_),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__nand2_1 _5758_ (.A(_1733_),
    .B(_1738_),
    .Y(_1739_));
 sky130_fd_sc_hd__o211ai_2 _5759_ (.A1(_1552_),
    .A2(_1580_),
    .B1(_1561_),
    .C1(_1567_),
    .Y(_1741_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(_1581_),
    .B(_1551_),
    .Y(_1742_));
 sky130_fd_sc_hd__nand2_1 _5761_ (.A(_1579_),
    .B(_1573_),
    .Y(_1743_));
 sky130_fd_sc_hd__o21ai_2 _5762_ (.A1(_1579_),
    .A2(_1576_),
    .B1(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__a21oi_1 _5763_ (.A1(_1550_),
    .A2(_1461_),
    .B1(_1459_),
    .Y(_1745_));
 sky130_fd_sc_hd__inv_2 _5764_ (.A(_1745_),
    .Y(_1746_));
 sky130_fd_sc_hd__nand2_1 _5765_ (.A(_1548_),
    .B(_1380_),
    .Y(_1747_));
 sky130_fd_sc_hd__nand3_2 _5766_ (.A(_1544_),
    .B(_1293_),
    .C(_1545_),
    .Y(_1748_));
 sky130_fd_sc_hd__and2_1 _5767_ (.A(_1541_),
    .B(_1543_),
    .X(_1749_));
 sky130_fd_sc_hd__or2_1 _5768_ (.A(_1219_),
    .B(_1749_),
    .X(_1750_));
 sky130_fd_sc_hd__inv_2 _5769_ (.A(_1750_),
    .Y(_1752_));
 sky130_fd_sc_hd__and3_1 _5770_ (.A(_1539_),
    .B(_1063_),
    .C(_1540_),
    .X(_1753_));
 sky130_fd_sc_hd__inv_2 _5771_ (.A(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__a21o_1 _5772_ (.A1(_1536_),
    .A2(_1538_),
    .B1(_0989_),
    .X(_1755_));
 sky130_fd_sc_hd__and2_1 _5773_ (.A(_1532_),
    .B(_0766_),
    .X(_1756_));
 sky130_fd_sc_hd__and3_2 _5774_ (.A(_1527_),
    .B(_0712_),
    .C(_1528_),
    .X(_1757_));
 sky130_fd_sc_hd__and3_2 _5775_ (.A(_1523_),
    .B(_0891_),
    .C(_1524_),
    .X(_1758_));
 sky130_fd_sc_hd__and3_1 _5776_ (.A(_1518_),
    .B(_0491_),
    .C(_1519_),
    .X(_1759_));
 sky130_fd_sc_hd__nand2_2 _5777_ (.A(_1505_),
    .B(_0198_),
    .Y(_1760_));
 sky130_fd_sc_hd__or2_1 _5778_ (.A(net143),
    .B(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__nand2_1 _5779_ (.A(net153),
    .B(_0184_),
    .Y(_1763_));
 sky130_fd_sc_hd__or2_1 _5780_ (.A(_1761_),
    .B(net154),
    .X(_1764_));
 sky130_fd_sc_hd__nand2_1 _5781_ (.A(_1507_),
    .B(_0874_),
    .Y(_1765_));
 sky130_fd_sc_hd__or2_1 _5782_ (.A(_1764_),
    .B(net170),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_2 _5783_ (.A(_1508_),
    .B(_0857_),
    .Y(_1767_));
 sky130_fd_sc_hd__nor2_1 _5784_ (.A(_1766_),
    .B(_1767_),
    .Y(_1768_));
 sky130_fd_sc_hd__inv_2 _5785_ (.A(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__nand2_1 _5786_ (.A(_1512_),
    .B(_0878_),
    .Y(_1770_));
 sky130_fd_sc_hd__nor2_1 _5787_ (.A(_1769_),
    .B(_1770_),
    .Y(_1771_));
 sky130_fd_sc_hd__inv_2 _5788_ (.A(_1771_),
    .Y(_1772_));
 sky130_fd_sc_hd__nor2_2 _5789_ (.A(_0811_),
    .B(_1515_),
    .Y(_1774_));
 sky130_fd_sc_hd__inv_2 _5790_ (.A(_1774_),
    .Y(_1775_));
 sky130_fd_sc_hd__nor2_1 _5791_ (.A(_1772_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__inv_2 _5792_ (.A(_1776_),
    .Y(_1777_));
 sky130_fd_sc_hd__a21o_1 _5793_ (.A1(_1516_),
    .A2(_1517_),
    .B1(_1041_),
    .X(_1778_));
 sky130_fd_sc_hd__nor2_1 _5794_ (.A(_1777_),
    .B(_1778_),
    .Y(_1779_));
 sky130_fd_sc_hd__nand2_1 _5795_ (.A(_1759_),
    .B(_1779_),
    .Y(_1780_));
 sky130_fd_sc_hd__a21o_1 _5796_ (.A1(_1521_),
    .A2(_1522_),
    .B1(_1046_),
    .X(_1781_));
 sky130_fd_sc_hd__nor2_1 _5797_ (.A(_1780_),
    .B(_1781_),
    .Y(_1782_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_1758_),
    .B(_1782_),
    .Y(_1783_));
 sky130_fd_sc_hd__a21o_1 _5799_ (.A1(_1525_),
    .A2(_1526_),
    .B1(_1199_),
    .X(_1785_));
 sky130_fd_sc_hd__nor2_1 _5800_ (.A(_1783_),
    .B(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__and3_1 _5801_ (.A(_1756_),
    .B(_1757_),
    .C(_1786_),
    .X(_1787_));
 sky130_fd_sc_hd__nand2_1 _5802_ (.A(_1503_),
    .B(_0766_),
    .Y(_1788_));
 sky130_fd_sc_hd__a21oi_2 _5803_ (.A1(_1533_),
    .A2(_1788_),
    .B1(_0906_),
    .Y(_1789_));
 sky130_fd_sc_hd__nand2_1 _5804_ (.A(_1787_),
    .B(_1789_),
    .Y(_1790_));
 sky130_fd_sc_hd__and3_1 _5805_ (.A(_1534_),
    .B(_0927_),
    .C(_1535_),
    .X(_1791_));
 sky130_fd_sc_hd__inv_2 _5806_ (.A(_1791_),
    .Y(_1792_));
 sky130_fd_sc_hd__nor2_1 _5807_ (.A(_1790_),
    .B(_1792_),
    .Y(_1793_));
 sky130_fd_sc_hd__inv_2 _5808_ (.A(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__nor2_1 _5809_ (.A(_1755_),
    .B(_1794_),
    .Y(_1796_));
 sky130_fd_sc_hd__inv_2 _5810_ (.A(_1796_),
    .Y(_1797_));
 sky130_fd_sc_hd__nor2_1 _5811_ (.A(_1754_),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__and2_1 _5812_ (.A(_1752_),
    .B(_1798_),
    .X(_1799_));
 sky130_fd_sc_hd__inv_2 _5813_ (.A(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__or2_1 _5814_ (.A(_1748_),
    .B(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__nor2_1 _5815_ (.A(_1747_),
    .B(_1801_),
    .Y(_1802_));
 sky130_fd_sc_hd__nor2_1 _5816_ (.A(_1461_),
    .B(_1550_),
    .Y(_1803_));
 sky130_fd_sc_hd__nand2_1 _5817_ (.A(_1802_),
    .B(_1803_),
    .Y(_1804_));
 sky130_fd_sc_hd__nor2_1 _5818_ (.A(_1746_),
    .B(_1804_),
    .Y(_1805_));
 sky130_fd_sc_hd__nand2_1 _5819_ (.A(_1805_),
    .B(_1570_),
    .Y(_1807_));
 sky130_fd_sc_hd__nor2_1 _5820_ (.A(_1744_),
    .B(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__nand3_2 _5821_ (.A(_1741_),
    .B(_1742_),
    .C(_1808_),
    .Y(_1809_));
 sky130_fd_sc_hd__inv_2 _5822_ (.A(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__nand2_1 _5823_ (.A(_1584_),
    .B(_1551_),
    .Y(_1811_));
 sky130_fd_sc_hd__nand2_1 _5824_ (.A(_1565_),
    .B(_1582_),
    .Y(_1812_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_1812_),
    .B(_1742_),
    .Y(_1813_));
 sky130_fd_sc_hd__nand3_2 _5826_ (.A(_1810_),
    .B(_1811_),
    .C(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__inv_2 _5827_ (.A(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__nand3_2 _5828_ (.A(_1589_),
    .B(_1739_),
    .C(_1815_),
    .Y(_1816_));
 sky130_fd_sc_hd__nor2_1 _5829_ (.A(_1723_),
    .B(_1726_),
    .Y(_1818_));
 sky130_fd_sc_hd__a21oi_1 _5830_ (.A1(_1683_),
    .A2(_1684_),
    .B1(_0707_),
    .Y(_1819_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(_1653_),
    .B(_1655_),
    .Y(_1820_));
 sky130_fd_sc_hd__nor2_1 _5832_ (.A(_0488_),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__nor2_1 _5833_ (.A(_0341_),
    .B(_1627_),
    .Y(_1822_));
 sky130_fd_sc_hd__mux2_2 _5834_ (.A0(net54),
    .A1(net22),
    .S(_1674_),
    .X(_1823_));
 sky130_fd_sc_hd__nor2_1 _5835_ (.A(_1599_),
    .B(_0314_),
    .Y(_1824_));
 sky130_fd_sc_hd__nand2_1 _5836_ (.A(_0162_),
    .B(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__nor2_1 _5837_ (.A(_1823_),
    .B(_1825_),
    .Y(_1826_));
 sky130_fd_sc_hd__nand2_1 _5838_ (.A(_1825_),
    .B(_1823_),
    .Y(_1827_));
 sky130_fd_sc_hd__or2b_1 _5839_ (.A(_1826_),
    .B_N(_1827_),
    .X(_1829_));
 sky130_fd_sc_hd__xor2_1 _5840_ (.A(_1829_),
    .B(_1606_),
    .X(_1830_));
 sky130_fd_sc_hd__nand3_1 _5841_ (.A(_1830_),
    .B(_1611_),
    .C(_1610_),
    .Y(_1831_));
 sky130_fd_sc_hd__inv_2 _5842_ (.A(_1830_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5843_ (.A(_1832_),
    .B(_1612_),
    .Y(_1833_));
 sky130_fd_sc_hd__nand2_1 _5844_ (.A(_1831_),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__inv_2 _5845_ (.A(_1834_),
    .Y(_1835_));
 sky130_fd_sc_hd__inv_2 _5846_ (.A(_1616_),
    .Y(_1836_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_1835_),
    .B(_1836_),
    .Y(_1837_));
 sky130_fd_sc_hd__nand2_1 _5848_ (.A(_1834_),
    .B(_1616_),
    .Y(_1838_));
 sky130_fd_sc_hd__nand2_1 _5849_ (.A(_1837_),
    .B(_1838_),
    .Y(_1840_));
 sky130_fd_sc_hd__inv_2 _5850_ (.A(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__inv_2 _5851_ (.A(_1625_),
    .Y(_1842_));
 sky130_fd_sc_hd__nand2_1 _5852_ (.A(_1841_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__nand2_1 _5853_ (.A(_1840_),
    .B(_1625_),
    .Y(_1844_));
 sky130_fd_sc_hd__nand3_1 _5854_ (.A(_1822_),
    .B(_1843_),
    .C(_1844_),
    .Y(_1845_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_1843_),
    .B(_1844_),
    .Y(_1846_));
 sky130_fd_sc_hd__nand2_1 _5856_ (.A(_1846_),
    .B(_1622_),
    .Y(_1847_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(_1845_),
    .B(_1847_),
    .Y(_1848_));
 sky130_fd_sc_hd__nand2_1 _5858_ (.A(_1848_),
    .B(_1629_),
    .Y(_1849_));
 sky130_fd_sc_hd__nand2_1 _5859_ (.A(_1636_),
    .B(_1639_),
    .Y(_1851_));
 sky130_fd_sc_hd__nand3_1 _5860_ (.A(_1847_),
    .B(_1851_),
    .C(_1623_),
    .Y(_1852_));
 sky130_fd_sc_hd__nand2_1 _5861_ (.A(_1849_),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__nand2_1 _5862_ (.A(_1853_),
    .B(_1645_),
    .Y(_1854_));
 sky130_fd_sc_hd__or2b_1 _5863_ (.A(_1646_),
    .B_N(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__nor2_1 _5864_ (.A(_0345_),
    .B(_1642_),
    .Y(_1856_));
 sky130_fd_sc_hd__nand3_1 _5865_ (.A(_1856_),
    .B(_1852_),
    .C(_1849_),
    .Y(_1857_));
 sky130_fd_sc_hd__nand2_1 _5866_ (.A(_1857_),
    .B(_1854_),
    .Y(_1858_));
 sky130_fd_sc_hd__nand2_1 _5867_ (.A(_1858_),
    .B(_1646_),
    .Y(_1859_));
 sky130_fd_sc_hd__nand2_1 _5868_ (.A(_1855_),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(_1860_),
    .B(_1649_),
    .Y(_1862_));
 sky130_fd_sc_hd__nor2_1 _5870_ (.A(_0394_),
    .B(_1650_),
    .Y(_1863_));
 sky130_fd_sc_hd__nand3_1 _5871_ (.A(_1863_),
    .B(_1859_),
    .C(_1855_),
    .Y(_1864_));
 sky130_fd_sc_hd__nand2_1 _5872_ (.A(_1862_),
    .B(_1864_),
    .Y(_1865_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(_1865_),
    .B(_1653_),
    .Y(_1866_));
 sky130_fd_sc_hd__nor2_1 _5874_ (.A(_0442_),
    .B(_1654_),
    .Y(_1867_));
 sky130_fd_sc_hd__nand3_1 _5875_ (.A(_1867_),
    .B(_1864_),
    .C(_1862_),
    .Y(_1868_));
 sky130_fd_sc_hd__nand3_1 _5876_ (.A(_1821_),
    .B(_1866_),
    .C(_1868_),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_1 _5877_ (.A(_1868_),
    .B(_1866_),
    .Y(_1870_));
 sky130_fd_sc_hd__nand2_1 _5878_ (.A(_1870_),
    .B(_1656_),
    .Y(_1871_));
 sky130_fd_sc_hd__nand2_1 _5879_ (.A(_1869_),
    .B(_1871_),
    .Y(_1873_));
 sky130_fd_sc_hd__nand2_1 _5880_ (.A(_1873_),
    .B(_1672_),
    .Y(_1874_));
 sky130_fd_sc_hd__nor2_1 _5881_ (.A(_0538_),
    .B(_1669_),
    .Y(_1875_));
 sky130_fd_sc_hd__nand3_1 _5882_ (.A(_1875_),
    .B(_1869_),
    .C(_1871_),
    .Y(_1876_));
 sky130_fd_sc_hd__nand2_1 _5883_ (.A(_1874_),
    .B(_1876_),
    .Y(_1877_));
 sky130_fd_sc_hd__nand2_1 _5884_ (.A(_1877_),
    .B(_1677_),
    .Y(_1878_));
 sky130_fd_sc_hd__nor2_1 _5885_ (.A(_0593_),
    .B(_1673_),
    .Y(_1879_));
 sky130_fd_sc_hd__nand2_1 _5886_ (.A(_1879_),
    .B(_1874_),
    .Y(_1880_));
 sky130_fd_sc_hd__nor2_1 _5887_ (.A(_1673_),
    .B(_0650_),
    .Y(_1881_));
 sky130_fd_sc_hd__nand3_1 _5888_ (.A(_1878_),
    .B(_1880_),
    .C(_1881_),
    .Y(_1882_));
 sky130_fd_sc_hd__nand2_1 _5889_ (.A(_1878_),
    .B(_1880_),
    .Y(_1884_));
 sky130_fd_sc_hd__inv_2 _5890_ (.A(_1881_),
    .Y(_1885_));
 sky130_fd_sc_hd__nand2_1 _5891_ (.A(_1884_),
    .B(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__nand3_1 _5892_ (.A(_1819_),
    .B(_1882_),
    .C(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__nand2_1 _5893_ (.A(_1886_),
    .B(_1882_),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_1 _5894_ (.A(_1888_),
    .B(_1688_),
    .Y(_1889_));
 sky130_fd_sc_hd__nand2_1 _5895_ (.A(_1887_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__inv_2 _5896_ (.A(_1686_),
    .Y(_1891_));
 sky130_fd_sc_hd__nor2_1 _5897_ (.A(_1891_),
    .B(_0778_),
    .Y(_1892_));
 sky130_fd_sc_hd__inv_2 _5898_ (.A(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__nand2_1 _5899_ (.A(_1890_),
    .B(_1893_),
    .Y(_1895_));
 sky130_fd_sc_hd__nand3_1 _5900_ (.A(_1887_),
    .B(_1889_),
    .C(_1892_),
    .Y(_1896_));
 sky130_fd_sc_hd__nand2_1 _5901_ (.A(_1895_),
    .B(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__nor2_1 _5902_ (.A(_0845_),
    .B(_0779_),
    .Y(_1898_));
 sky130_fd_sc_hd__nand2_1 _5903_ (.A(_1898_),
    .B(_1692_),
    .Y(_1899_));
 sky130_fd_sc_hd__nand2_1 _5904_ (.A(_1897_),
    .B(_1899_),
    .Y(_1900_));
 sky130_fd_sc_hd__nand3b_1 _5905_ (.A_N(_1899_),
    .B(_1895_),
    .C(_1896_),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2_1 _5906_ (.A(_1900_),
    .B(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(_1902_),
    .B(_1697_),
    .Y(_1903_));
 sky130_fd_sc_hd__a21oi_1 _5908_ (.A1(_1691_),
    .A2(_1693_),
    .B1(_0921_),
    .Y(_1904_));
 sky130_fd_sc_hd__nand3_1 _5909_ (.A(_1904_),
    .B(_1900_),
    .C(_1901_),
    .Y(_1906_));
 sky130_fd_sc_hd__nand2_1 _5910_ (.A(_1903_),
    .B(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__nand2_1 _5911_ (.A(_1907_),
    .B(_1701_),
    .Y(_1908_));
 sky130_fd_sc_hd__a21oi_1 _5912_ (.A1(_1693_),
    .A2(_1691_),
    .B1(_1006_),
    .Y(_1909_));
 sky130_fd_sc_hd__nand3_1 _5913_ (.A(_1903_),
    .B(_1906_),
    .C(_1909_),
    .Y(_1910_));
 sky130_fd_sc_hd__nand2_1 _5914_ (.A(_1908_),
    .B(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__nor2_1 _5915_ (.A(_1086_),
    .B(_1702_),
    .Y(_1912_));
 sky130_fd_sc_hd__inv_2 _5916_ (.A(_1912_),
    .Y(_1913_));
 sky130_fd_sc_hd__nand2_1 _5917_ (.A(_1911_),
    .B(_1913_),
    .Y(_1914_));
 sky130_fd_sc_hd__nand2_1 _5918_ (.A(_1912_),
    .B(_1908_),
    .Y(_1915_));
 sky130_fd_sc_hd__nand2_1 _5919_ (.A(_1914_),
    .B(_1915_),
    .Y(_1917_));
 sky130_fd_sc_hd__nand2_1 _5920_ (.A(_1917_),
    .B(_1704_),
    .Y(_1918_));
 sky130_fd_sc_hd__nor2_1 _5921_ (.A(_1702_),
    .B(_1156_),
    .Y(_1919_));
 sky130_fd_sc_hd__nand3_2 _5922_ (.A(_1914_),
    .B(_1915_),
    .C(_1919_),
    .Y(_1920_));
 sky130_fd_sc_hd__nand2_1 _5923_ (.A(_1918_),
    .B(_1920_),
    .Y(_1921_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(_1921_),
    .B(_1711_),
    .Y(_1922_));
 sky130_fd_sc_hd__nor2_1 _5925_ (.A(_1232_),
    .B(_1712_),
    .Y(_1923_));
 sky130_fd_sc_hd__nand3_1 _5926_ (.A(_1918_),
    .B(_1923_),
    .C(_1920_),
    .Y(_1924_));
 sky130_fd_sc_hd__nand2_1 _5927_ (.A(_1922_),
    .B(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__nand2_1 _5928_ (.A(_1925_),
    .B(_1717_),
    .Y(_1926_));
 sky130_fd_sc_hd__nand2_1 _5929_ (.A(_1922_),
    .B(_1716_),
    .Y(_1928_));
 sky130_fd_sc_hd__nand2_1 _5930_ (.A(_1926_),
    .B(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__nor2_1 _5931_ (.A(_1396_),
    .B(_1719_),
    .Y(_1930_));
 sky130_fd_sc_hd__inv_2 _5932_ (.A(_1930_),
    .Y(_1931_));
 sky130_fd_sc_hd__nand2_1 _5933_ (.A(_1929_),
    .B(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__nand3_2 _5934_ (.A(_1930_),
    .B(_1926_),
    .C(_1928_),
    .Y(_1933_));
 sky130_fd_sc_hd__nor2_1 _5935_ (.A(_1719_),
    .B(_1491_),
    .Y(_1934_));
 sky130_fd_sc_hd__nand3_2 _5936_ (.A(_1932_),
    .B(_1933_),
    .C(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__nand2_1 _5937_ (.A(_1932_),
    .B(_1933_),
    .Y(_1936_));
 sky130_fd_sc_hd__inv_2 _5938_ (.A(_1934_),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _5939_ (.A(_1936_),
    .B(_1937_),
    .Y(_1939_));
 sky130_fd_sc_hd__nand3_1 _5940_ (.A(_1818_),
    .B(_1935_),
    .C(_1939_),
    .Y(_1940_));
 sky130_fd_sc_hd__nand2_1 _5941_ (.A(_1939_),
    .B(_1935_),
    .Y(_1941_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_1941_),
    .B(_1735_),
    .Y(_1942_));
 sky130_fd_sc_hd__nand2_1 _5943_ (.A(_1940_),
    .B(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__inv_2 _5944_ (.A(_1943_),
    .Y(_1944_));
 sky130_fd_sc_hd__nor2_1 _5945_ (.A(_1731_),
    .B(_1734_),
    .Y(_1945_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(_1944_),
    .B(_1945_),
    .Y(_1946_));
 sky130_fd_sc_hd__nand3_1 _5947_ (.A(_1737_),
    .B(_1556_),
    .C(_1732_),
    .Y(_1947_));
 sky130_fd_sc_hd__nand2_1 _5948_ (.A(_1943_),
    .B(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__nand2_1 _5949_ (.A(_1946_),
    .B(_1948_),
    .Y(_1950_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_2736_),
    .B(_2740_),
    .Y(_1951_));
 sky130_fd_sc_hd__nand2_1 _5951_ (.A(_1950_),
    .B(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__o21ai_1 _5952_ (.A1(_0081_),
    .A2(_1816_),
    .B1(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__a21oi_1 _5953_ (.A1(_1588_),
    .A2(_1554_),
    .B1(_1814_),
    .Y(_1954_));
 sky130_fd_sc_hd__nand3_1 _5954_ (.A(_1954_),
    .B(_1950_),
    .C(_1739_),
    .Y(_1955_));
 sky130_fd_sc_hd__nand2_1 _5955_ (.A(_1953_),
    .B(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__nand2_1 _5956_ (.A(_1950_),
    .B(_0081_),
    .Y(_1957_));
 sky130_fd_sc_hd__nand2_1 _5957_ (.A(_1956_),
    .B(_1957_),
    .Y(_1958_));
 sky130_fd_sc_hd__inv_2 _5958_ (.A(_1958_),
    .Y(_1959_));
 sky130_fd_sc_hd__inv_2 _5959_ (.A(_1816_),
    .Y(_1961_));
 sky130_fd_sc_hd__nand3_1 _5960_ (.A(_1961_),
    .B(_0078_),
    .C(_1950_),
    .Y(_1962_));
 sky130_fd_sc_hd__nor2_1 _5961_ (.A(_1731_),
    .B(_1585_),
    .Y(_1963_));
 sky130_fd_sc_hd__nand2_1 _5962_ (.A(_1963_),
    .B(_1943_),
    .Y(_1964_));
 sky130_fd_sc_hd__nand2_1 _5963_ (.A(_1904_),
    .B(_1900_),
    .Y(_1965_));
 sky130_fd_sc_hd__nand2_1 _5964_ (.A(_1965_),
    .B(_1901_),
    .Y(_1966_));
 sky130_fd_sc_hd__nand2_1 _5965_ (.A(_1880_),
    .B(_1876_),
    .Y(_1967_));
 sky130_fd_sc_hd__nand2_2 _5966_ (.A(_1443_),
    .B(_1421_),
    .Y(_1968_));
 sky130_fd_sc_hd__inv_2 _5967_ (.A(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__a41o_1 _5968_ (.A1(_1603_),
    .A2(_0320_),
    .A3(_0321_),
    .A4(_1827_),
    .B1(_1826_),
    .X(_1970_));
 sky130_fd_sc_hd__xor2_1 _5969_ (.A(_1969_),
    .B(_1970_),
    .X(_1972_));
 sky130_fd_sc_hd__nand2_1 _5970_ (.A(_1837_),
    .B(_1831_),
    .Y(_1973_));
 sky130_fd_sc_hd__xnor2_1 _5971_ (.A(_1972_),
    .B(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__xor2_1 _5972_ (.A(_1843_),
    .B(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__nand2_1 _5973_ (.A(_1852_),
    .B(_1845_),
    .Y(_1976_));
 sky130_fd_sc_hd__xnor2_1 _5974_ (.A(_1975_),
    .B(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__nand2_1 _5975_ (.A(_1855_),
    .B(_1857_),
    .Y(_1978_));
 sky130_fd_sc_hd__xnor2_1 _5976_ (.A(_1977_),
    .B(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__a21bo_1 _5977_ (.A1(_1867_),
    .A2(_1862_),
    .B1_N(_1864_),
    .X(_1980_));
 sky130_fd_sc_hd__xnor2_1 _5978_ (.A(_1979_),
    .B(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__xor2_1 _5979_ (.A(_1869_),
    .B(_1981_),
    .X(_1983_));
 sky130_fd_sc_hd__xnor2_1 _5980_ (.A(_1967_),
    .B(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__xor2_1 _5981_ (.A(_1882_),
    .B(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__a21bo_1 _5982_ (.A1(_1889_),
    .A2(_1892_),
    .B1_N(_1887_),
    .X(_1986_));
 sky130_fd_sc_hd__xnor2_1 _5983_ (.A(_1985_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__xnor2_1 _5984_ (.A(_1966_),
    .B(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__nand2_1 _5985_ (.A(_1915_),
    .B(_1910_),
    .Y(_1989_));
 sky130_fd_sc_hd__or2_1 _5986_ (.A(_1988_),
    .B(_1989_),
    .X(_1990_));
 sky130_fd_sc_hd__nand2_1 _5987_ (.A(_1989_),
    .B(_1988_),
    .Y(_1991_));
 sky130_fd_sc_hd__nand2_1 _5988_ (.A(_1990_),
    .B(_1991_),
    .Y(_1992_));
 sky130_fd_sc_hd__inv_2 _5989_ (.A(_1920_),
    .Y(_1994_));
 sky130_fd_sc_hd__nand2_1 _5990_ (.A(_1992_),
    .B(_1994_),
    .Y(_1995_));
 sky130_fd_sc_hd__nand3_1 _5991_ (.A(_1990_),
    .B(_1991_),
    .C(_1920_),
    .Y(_1996_));
 sky130_fd_sc_hd__nand2_1 _5992_ (.A(_1995_),
    .B(_1996_),
    .Y(_1997_));
 sky130_fd_sc_hd__nand2_1 _5993_ (.A(_1928_),
    .B(_1924_),
    .Y(_1998_));
 sky130_fd_sc_hd__nor2_1 _5994_ (.A(_1997_),
    .B(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__and2_1 _5995_ (.A(_1998_),
    .B(_1997_),
    .X(_2000_));
 sky130_fd_sc_hd__o21bai_1 _5996_ (.A1(_1999_),
    .A2(_2000_),
    .B1_N(_1933_),
    .Y(_2001_));
 sky130_fd_sc_hd__or2_1 _5997_ (.A(_1997_),
    .B(_1998_),
    .X(_2002_));
 sky130_fd_sc_hd__nand2_1 _5998_ (.A(_1998_),
    .B(_1997_),
    .Y(_2003_));
 sky130_fd_sc_hd__nand3_1 _5999_ (.A(_2002_),
    .B(_2003_),
    .C(_1933_),
    .Y(_2005_));
 sky130_fd_sc_hd__nand2_1 _6000_ (.A(_2001_),
    .B(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__inv_2 _6001_ (.A(_1935_),
    .Y(_2007_));
 sky130_fd_sc_hd__nand2_1 _6002_ (.A(_2006_),
    .B(_2007_),
    .Y(_2008_));
 sky130_fd_sc_hd__nand3_1 _6003_ (.A(_2001_),
    .B(_1935_),
    .C(_2005_),
    .Y(_2009_));
 sky130_fd_sc_hd__nand2_1 _6004_ (.A(_2008_),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__inv_2 _6005_ (.A(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__nand2_1 _6006_ (.A(_1964_),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__nand3_1 _6007_ (.A(_2010_),
    .B(_1963_),
    .C(_1943_),
    .Y(_2013_));
 sky130_fd_sc_hd__nand2_1 _6008_ (.A(_2012_),
    .B(_2013_),
    .Y(_2014_));
 sky130_fd_sc_hd__inv_2 _6009_ (.A(_2014_),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _6010_ (.A(_2014_),
    .B(_0078_),
    .Y(_2017_));
 sky130_fd_sc_hd__nor2_1 _6011_ (.A(_2017_),
    .B(_1955_),
    .Y(_2018_));
 sky130_fd_sc_hd__a21oi_1 _6012_ (.A1(_1962_),
    .A2(_2016_),
    .B1(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__nor2_1 _6013_ (.A(_0081_),
    .B(_1814_),
    .Y(_2020_));
 sky130_fd_sc_hd__nand2_1 _6014_ (.A(_1589_),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(_1739_),
    .B(_1951_),
    .Y(_2022_));
 sky130_fd_sc_hd__nand2_1 _6016_ (.A(_2021_),
    .B(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__nand2_1 _6017_ (.A(_2023_),
    .B(_1816_),
    .Y(_2024_));
 sky130_fd_sc_hd__nand2_1 _6018_ (.A(_1739_),
    .B(_0081_),
    .Y(_2025_));
 sky130_fd_sc_hd__nand2_1 _6019_ (.A(_2024_),
    .B(_2025_),
    .Y(_2027_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(_1811_),
    .B(_1813_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _6021_ (.A(_1814_),
    .B(_0078_),
    .Y(_2029_));
 sky130_fd_sc_hd__o21ai_1 _6022_ (.A1(_0078_),
    .A2(_2028_),
    .B1(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__inv_2 _6023_ (.A(_0061_),
    .Y(_2031_));
 sky130_fd_sc_hd__nor2_1 _6024_ (.A(net67),
    .B(_0073_),
    .Y(_2032_));
 sky130_fd_sc_hd__a21o_1 _6025_ (.A1(_0061_),
    .A2(_0065_),
    .B1(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__a21oi_4 _6026_ (.A1(_2031_),
    .A2(_0063_),
    .B1(_2033_),
    .Y(_2034_));
 sky130_fd_sc_hd__inv_2 _6027_ (.A(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__o21ai_1 _6028_ (.A1(_2035_),
    .A2(_1809_),
    .B1(_2028_),
    .Y(_2036_));
 sky130_fd_sc_hd__nand2_1 _6029_ (.A(_1741_),
    .B(_1742_),
    .Y(_2038_));
 sky130_fd_sc_hd__nand2_1 _6030_ (.A(_1809_),
    .B(_0077_),
    .Y(_2039_));
 sky130_fd_sc_hd__o21ai_1 _6031_ (.A1(_0077_),
    .A2(_2038_),
    .B1(_2039_),
    .Y(_2040_));
 sky130_fd_sc_hd__a22o_1 _6032_ (.A1(_1808_),
    .A2(_2034_),
    .B1(_1741_),
    .B2(_1742_),
    .X(_2041_));
 sky130_fd_sc_hd__nand2_1 _6033_ (.A(_2040_),
    .B(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__and2_1 _6034_ (.A(_1807_),
    .B(_1744_),
    .X(_2043_));
 sky130_fd_sc_hd__o21ai_1 _6035_ (.A1(_0069_),
    .A2(_1744_),
    .B1(_0067_),
    .Y(_2044_));
 sky130_fd_sc_hd__and2_1 _6036_ (.A(_2741_),
    .B(_0076_),
    .X(_2045_));
 sky130_fd_sc_hd__nand2_1 _6037_ (.A(_2044_),
    .B(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__o21ai_1 _6038_ (.A1(_1808_),
    .A2(_2043_),
    .B1(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__nand2_1 _6039_ (.A(_0081_),
    .B(_1744_),
    .Y(_2049_));
 sky130_fd_sc_hd__nor2_2 _6040_ (.A(_2740_),
    .B(_0067_),
    .Y(_2050_));
 sky130_fd_sc_hd__o21ai_1 _6041_ (.A1(_0075_),
    .A2(_1570_),
    .B1(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__nand2_1 _6042_ (.A(_0072_),
    .B(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__inv_2 _6043_ (.A(_1805_),
    .Y(_2053_));
 sky130_fd_sc_hd__nand2_1 _6044_ (.A(_2053_),
    .B(_1577_),
    .Y(_2054_));
 sky130_fd_sc_hd__nand3_1 _6045_ (.A(_2052_),
    .B(_1807_),
    .C(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__o21ai_1 _6046_ (.A1(_0077_),
    .A2(_1577_),
    .B1(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__a21oi_1 _6047_ (.A1(_2047_),
    .A2(_2049_),
    .B1(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__nand2_1 _6048_ (.A(_2042_),
    .B(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__a21oi_1 _6049_ (.A1(_2030_),
    .A2(_2036_),
    .B1(_2058_),
    .Y(_2060_));
 sky130_fd_sc_hd__inv_2 _6050_ (.A(_1954_),
    .Y(_2061_));
 sky130_fd_sc_hd__nand2_1 _6051_ (.A(_1589_),
    .B(_1951_),
    .Y(_2062_));
 sky130_fd_sc_hd__inv_2 _6052_ (.A(_2020_),
    .Y(_2063_));
 sky130_fd_sc_hd__nand2_1 _6053_ (.A(_2062_),
    .B(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__nand2_1 _6054_ (.A(_2061_),
    .B(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__nand2_1 _6055_ (.A(_1589_),
    .B(_0081_),
    .Y(_2066_));
 sky130_fd_sc_hd__nand3_1 _6056_ (.A(_2060_),
    .B(_2065_),
    .C(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__nor2_1 _6057_ (.A(_2027_),
    .B(_2067_),
    .Y(_2068_));
 sky130_fd_sc_hd__nand3_1 _6058_ (.A(_1959_),
    .B(_2019_),
    .C(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__and3_1 _6059_ (.A(_0158_),
    .B(_1824_),
    .C(_0101_),
    .X(_2071_));
 sky130_fd_sc_hd__or4b_4 _6060_ (.A(_1968_),
    .B(_0113_),
    .C(_1823_),
    .D_N(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__clkbuf_1 _6061_ (.A(net126),
    .X(_2073_));
 sky130_fd_sc_hd__a21oi_1 _6062_ (.A1(_2069_),
    .A2(_2072_),
    .B1(net120),
    .Y(_0035_));
 sky130_fd_sc_hd__nand2_1 _6063_ (.A(_1962_),
    .B(_2016_),
    .Y(_2074_));
 sky130_fd_sc_hd__o21ai_1 _6064_ (.A1(_1955_),
    .A2(_2017_),
    .B1(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__nand3_1 _6065_ (.A(_2047_),
    .B(_2056_),
    .C(_2049_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand3b_1 _6066_ (.A_N(_2076_),
    .B(_2040_),
    .C(_2041_),
    .Y(_2077_));
 sky130_fd_sc_hd__inv_2 _6067_ (.A(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__nand3_1 _6068_ (.A(_2078_),
    .B(_2030_),
    .C(_2036_),
    .Y(_2079_));
 sky130_fd_sc_hd__nand2_1 _6069_ (.A(_2065_),
    .B(_2066_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_2081_),
    .B(_2027_),
    .Y(_2082_));
 sky130_fd_sc_hd__nor2_1 _6071_ (.A(_2079_),
    .B(_2082_),
    .Y(_2083_));
 sky130_fd_sc_hd__nand3_1 _6072_ (.A(_2075_),
    .B(_2083_),
    .C(_1958_),
    .Y(_2084_));
 sky130_fd_sc_hd__nand2_1 _6073_ (.A(_1823_),
    .B(_0314_),
    .Y(_2085_));
 sky130_fd_sc_hd__or4_1 _6074_ (.A(_1969_),
    .B(_0095_),
    .C(_0153_),
    .D(_0091_),
    .X(_2086_));
 sky130_fd_sc_hd__or4_4 _6075_ (.A(_0089_),
    .B(_1600_),
    .C(_2085_),
    .D(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__a21oi_1 _6076_ (.A1(_2084_),
    .A2(_2087_),
    .B1(net120),
    .Y(_0034_));
 sky130_fd_sc_hd__nand2_1 _6077_ (.A(net131),
    .B(_0893_),
    .Y(_2088_));
 sky130_fd_sc_hd__inv_2 _6078_ (.A(net143),
    .Y(_2089_));
 sky130_fd_sc_hd__inv_2 _6079_ (.A(_0067_),
    .Y(_2091_));
 sky130_fd_sc_hd__nor2_2 _6080_ (.A(_0069_),
    .B(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__inv_2 _6081_ (.A(_2050_),
    .Y(_2093_));
 sky130_fd_sc_hd__nor2_4 _6082_ (.A(_0075_),
    .B(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__a2111o_1 _6083_ (.A1(_2740_),
    .A2(_2088_),
    .B1(_2089_),
    .C1(_2092_),
    .D1(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__inv_2 _6084_ (.A(_2094_),
    .Y(_2096_));
 sky130_fd_sc_hd__inv_2 _6085_ (.A(_2092_),
    .Y(_2097_));
 sky130_fd_sc_hd__clkbuf_4 _6086_ (.A(net138),
    .X(_2098_));
 sky130_fd_sc_hd__buf_2 _6087_ (.A(_2740_),
    .X(_2099_));
 sky130_fd_sc_hd__nand2_1 _6088_ (.A(_2098_),
    .B(_2099_),
    .Y(_2100_));
 sky130_fd_sc_hd__a31o_1 _6089_ (.A1(_2096_),
    .A2(_2097_),
    .A3(_2100_),
    .B1(net143),
    .X(_2102_));
 sky130_fd_sc_hd__a21o_1 _6090_ (.A1(_2095_),
    .A2(_2102_),
    .B1(net120),
    .X(_2103_));
 sky130_fd_sc_hd__inv_2 _6091_ (.A(_2103_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _6092_ (.A(_2740_),
    .Y(_2104_));
 sky130_fd_sc_hd__a21oi_1 _6093_ (.A1(_0070_),
    .A2(_0076_),
    .B1(_1761_),
    .Y(_2105_));
 sky130_fd_sc_hd__a31o_1 _6094_ (.A1(_0076_),
    .A2(_0070_),
    .A3(_1760_),
    .B1(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__nand2_1 _6095_ (.A(net180),
    .B(_2098_),
    .Y(_2107_));
 sky130_fd_sc_hd__o31a_1 _6096_ (.A1(_2098_),
    .A2(_1761_),
    .A3(_2035_),
    .B1(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__o21ai_1 _6097_ (.A1(net143),
    .A2(_2035_),
    .B1(net180),
    .Y(_2109_));
 sky130_fd_sc_hd__o21ai_1 _6098_ (.A1(_2104_),
    .A2(_2108_),
    .B1(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__a211o_1 _6099_ (.A1(_2104_),
    .A2(_2106_),
    .B1(net120),
    .C1(_2110_),
    .X(_2112_));
 sky130_fd_sc_hd__inv_2 _6100_ (.A(_2112_),
    .Y(_0013_));
 sky130_fd_sc_hd__nand2_1 _6101_ (.A(net154),
    .B(_1761_),
    .Y(_2113_));
 sky130_fd_sc_hd__nand2_1 _6102_ (.A(_1764_),
    .B(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__mux2_1 _6103_ (.A0(_2114_),
    .A1(net154),
    .S(net138),
    .X(_2115_));
 sky130_fd_sc_hd__mux2_1 _6104_ (.A0(_2115_),
    .A1(net154),
    .S(_0074_),
    .X(_2116_));
 sky130_fd_sc_hd__inv_2 _6105_ (.A(_0070_),
    .Y(_2117_));
 sky130_fd_sc_hd__a22o_1 _6106_ (.A1(_2117_),
    .A2(_2114_),
    .B1(_2092_),
    .B2(net154),
    .X(_2118_));
 sky130_fd_sc_hd__a221o_1 _6107_ (.A1(_2740_),
    .A2(_2115_),
    .B1(_2050_),
    .B2(_2116_),
    .C1(net155),
    .X(_2119_));
 sky130_fd_sc_hd__nor2_1 _6108_ (.A(net120),
    .B(net156),
    .Y(_0024_));
 sky130_fd_sc_hd__or2b_1 _6109_ (.A(net154),
    .B_N(_2119_),
    .X(_2121_));
 sky130_fd_sc_hd__clkbuf_4 _6110_ (.A(net126),
    .X(_2122_));
 sky130_fd_sc_hd__a21oi_1 _6111_ (.A1(_0072_),
    .A2(_0076_),
    .B1(_1766_),
    .Y(_2123_));
 sky130_fd_sc_hd__a211o_1 _6112_ (.A1(_2121_),
    .A2(net170),
    .B1(_2122_),
    .C1(_2123_),
    .X(_2124_));
 sky130_fd_sc_hd__inv_2 _6113_ (.A(_2124_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _6114_ (.A(_1767_),
    .Y(_2125_));
 sky130_fd_sc_hd__nand2_1 _6115_ (.A(_0078_),
    .B(_1768_),
    .Y(_2126_));
 sky130_fd_sc_hd__o211ai_2 _6116_ (.A1(_2125_),
    .A2(_2123_),
    .B1(_0079_),
    .C1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__inv_2 _6117_ (.A(_2127_),
    .Y(_0028_));
 sky130_fd_sc_hd__a221o_1 _6118_ (.A1(_0078_),
    .A2(_1771_),
    .B1(_2126_),
    .B2(net178),
    .C1(_2122_),
    .X(_2128_));
 sky130_fd_sc_hd__inv_2 _6119_ (.A(_2128_),
    .Y(_0029_));
 sky130_fd_sc_hd__nand2_1 _6120_ (.A(_0078_),
    .B(_1771_),
    .Y(_2130_));
 sky130_fd_sc_hd__a21oi_1 _6121_ (.A1(_2130_),
    .A2(_1775_),
    .B1(_1776_),
    .Y(_2131_));
 sky130_fd_sc_hd__a31o_1 _6122_ (.A1(_2045_),
    .A2(_0070_),
    .A3(_1774_),
    .B1(_2035_),
    .X(_2132_));
 sky130_fd_sc_hd__o221ai_2 _6123_ (.A1(_2034_),
    .A2(_1774_),
    .B1(_2131_),
    .B2(_2132_),
    .C1(_0079_),
    .Y(_2133_));
 sky130_fd_sc_hd__inv_2 _6124_ (.A(_2133_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_1 _6125_ (.A(_1778_),
    .B(_1777_),
    .Y(_2134_));
 sky130_fd_sc_hd__or2b_1 _6126_ (.A(_1779_),
    .B_N(_2134_),
    .X(_2135_));
 sky130_fd_sc_hd__inv_2 _6127_ (.A(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__nand2_1 _6128_ (.A(_1778_),
    .B(_2098_),
    .Y(_2137_));
 sky130_fd_sc_hd__o21a_1 _6129_ (.A1(_2098_),
    .A2(_2136_),
    .B1(_2137_),
    .X(_2139_));
 sky130_fd_sc_hd__clkbuf_4 _6130_ (.A(_0075_),
    .X(_2140_));
 sky130_fd_sc_hd__nand2_1 _6131_ (.A(_2135_),
    .B(_2140_),
    .Y(_2141_));
 sky130_fd_sc_hd__o21ai_1 _6132_ (.A1(_2092_),
    .A2(_2094_),
    .B1(_1778_),
    .Y(_2142_));
 sky130_fd_sc_hd__o211a_1 _6133_ (.A1(_0070_),
    .A2(_2136_),
    .B1(_2141_),
    .C1(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__o211ai_2 _6134_ (.A1(_2104_),
    .A2(_2139_),
    .B1(_0079_),
    .C1(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__inv_2 _6135_ (.A(_2144_),
    .Y(_0031_));
 sky130_fd_sc_hd__or2_1 _6136_ (.A(_1779_),
    .B(_1759_),
    .X(_2145_));
 sky130_fd_sc_hd__nand2_1 _6137_ (.A(_2145_),
    .B(_1780_),
    .Y(_2146_));
 sky130_fd_sc_hd__inv_2 _6138_ (.A(_2146_),
    .Y(_2147_));
 sky130_fd_sc_hd__mux2_1 _6139_ (.A0(_2147_),
    .A1(_1759_),
    .S(_2098_),
    .X(_2149_));
 sky130_fd_sc_hd__nor2_1 _6140_ (.A(_2104_),
    .B(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__a21o_1 _6141_ (.A1(_2096_),
    .A2(_2097_),
    .B1(_1759_),
    .X(_2151_));
 sky130_fd_sc_hd__o21ai_1 _6142_ (.A1(_0070_),
    .A2(_2147_),
    .B1(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__a2111o_1 _6143_ (.A1(_2140_),
    .A2(_2146_),
    .B1(net126),
    .C1(_2150_),
    .D1(net133),
    .X(_2153_));
 sky130_fd_sc_hd__inv_2 _6144_ (.A(net134),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2_1 _6145_ (.A(_1781_),
    .B(_1780_),
    .Y(_2154_));
 sky130_fd_sc_hd__or2b_1 _6146_ (.A(_1782_),
    .B_N(_2154_),
    .X(_2155_));
 sky130_fd_sc_hd__mux2_1 _6147_ (.A0(_2155_),
    .A1(_1781_),
    .S(_2098_),
    .X(_2156_));
 sky130_fd_sc_hd__mux2_1 _6148_ (.A0(_2155_),
    .A1(_1781_),
    .S(net132),
    .X(_2157_));
 sky130_fd_sc_hd__a22o_1 _6149_ (.A1(_0075_),
    .A2(_2155_),
    .B1(_2094_),
    .B2(_1781_),
    .X(_2159_));
 sky130_fd_sc_hd__a21o_1 _6150_ (.A1(_0067_),
    .A2(_2157_),
    .B1(_2159_),
    .X(_2160_));
 sky130_fd_sc_hd__a211o_1 _6151_ (.A1(_2099_),
    .A2(_2156_),
    .B1(_2122_),
    .C1(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__inv_2 _6152_ (.A(_2161_),
    .Y(_0033_));
 sky130_fd_sc_hd__nand2_1 _6153_ (.A(_1758_),
    .B(_0076_),
    .Y(_2162_));
 sky130_fd_sc_hd__a21o_1 _6154_ (.A1(_2050_),
    .A2(_2162_),
    .B1(_0071_),
    .X(_2163_));
 sky130_fd_sc_hd__or2_1 _6155_ (.A(_1782_),
    .B(_1758_),
    .X(_2164_));
 sky130_fd_sc_hd__nand2_1 _6156_ (.A(_2164_),
    .B(_1783_),
    .Y(_2165_));
 sky130_fd_sc_hd__nor2_1 _6157_ (.A(_1758_),
    .B(_0078_),
    .Y(_2166_));
 sky130_fd_sc_hd__a311o_1 _6158_ (.A1(_2163_),
    .A2(_2034_),
    .A3(_2165_),
    .B1(_2122_),
    .C1(_2166_),
    .X(_2167_));
 sky130_fd_sc_hd__inv_2 _6159_ (.A(_2167_),
    .Y(_0003_));
 sky130_fd_sc_hd__o21ai_1 _6160_ (.A1(_2140_),
    .A2(_1785_),
    .B1(_2050_),
    .Y(_2169_));
 sky130_fd_sc_hd__a21oi_1 _6161_ (.A1(_0072_),
    .A2(_2169_),
    .B1(_2035_),
    .Y(_2170_));
 sky130_fd_sc_hd__nand2_1 _6162_ (.A(_1785_),
    .B(_1783_),
    .Y(_2171_));
 sky130_fd_sc_hd__or2b_1 _6163_ (.A(_1786_),
    .B_N(_2171_),
    .X(_2172_));
 sky130_fd_sc_hd__a221o_1 _6164_ (.A1(_0081_),
    .A2(_1785_),
    .B1(_2170_),
    .B2(_2172_),
    .C1(_2122_),
    .X(_2173_));
 sky130_fd_sc_hd__inv_2 _6165_ (.A(_2173_),
    .Y(_0004_));
 sky130_fd_sc_hd__or2_1 _6166_ (.A(_1786_),
    .B(_1757_),
    .X(_2174_));
 sky130_fd_sc_hd__nand2_1 _6167_ (.A(_1757_),
    .B(_1786_),
    .Y(_2175_));
 sky130_fd_sc_hd__nand2_1 _6168_ (.A(_2174_),
    .B(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__nand2_1 _6169_ (.A(_2176_),
    .B(_0893_),
    .Y(_2178_));
 sky130_fd_sc_hd__o21ai_1 _6170_ (.A1(_0893_),
    .A2(_1757_),
    .B1(_2178_),
    .Y(_2179_));
 sky130_fd_sc_hd__or2_1 _6171_ (.A(_1757_),
    .B(_0069_),
    .X(_2180_));
 sky130_fd_sc_hd__nand2_1 _6172_ (.A(_0069_),
    .B(_2176_),
    .Y(_2181_));
 sky130_fd_sc_hd__a21oi_1 _6173_ (.A1(_2180_),
    .A2(_2181_),
    .B1(_2091_),
    .Y(_2182_));
 sky130_fd_sc_hd__a2bb2o_1 _6174_ (.A1_N(_1757_),
    .A2_N(_2096_),
    .B1(_2140_),
    .B2(_2176_),
    .X(_2183_));
 sky130_fd_sc_hd__a2111o_1 _6175_ (.A1(_2099_),
    .A2(_2179_),
    .B1(net126),
    .C1(_2182_),
    .D1(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__inv_2 _6176_ (.A(_2184_),
    .Y(_0005_));
 sky130_fd_sc_hd__nand2_1 _6177_ (.A(_1756_),
    .B(_0076_),
    .Y(_2185_));
 sky130_fd_sc_hd__a21o_1 _6178_ (.A1(_2050_),
    .A2(_2185_),
    .B1(_0071_),
    .X(_2186_));
 sky130_fd_sc_hd__xor2_1 _6179_ (.A(_2175_),
    .B(_1756_),
    .X(_2188_));
 sky130_fd_sc_hd__nor2_1 _6180_ (.A(_1756_),
    .B(_0078_),
    .Y(_2189_));
 sky130_fd_sc_hd__a211o_1 _6181_ (.A1(_2186_),
    .A2(_2188_),
    .B1(_2122_),
    .C1(_2189_),
    .X(_2190_));
 sky130_fd_sc_hd__inv_2 _6182_ (.A(_2190_),
    .Y(_0006_));
 sky130_fd_sc_hd__or2_1 _6183_ (.A(_1789_),
    .B(_1787_),
    .X(_2191_));
 sky130_fd_sc_hd__nand2_1 _6184_ (.A(_2191_),
    .B(_1790_),
    .Y(_2192_));
 sky130_fd_sc_hd__nand2_1 _6185_ (.A(_2192_),
    .B(_0893_),
    .Y(_2193_));
 sky130_fd_sc_hd__o21ai_1 _6186_ (.A1(_0893_),
    .A2(_1789_),
    .B1(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__or2_1 _6187_ (.A(_1789_),
    .B(_0069_),
    .X(_2195_));
 sky130_fd_sc_hd__nand2_1 _6188_ (.A(_0069_),
    .B(_2192_),
    .Y(_2196_));
 sky130_fd_sc_hd__a21oi_1 _6189_ (.A1(_2195_),
    .A2(_2196_),
    .B1(_2091_),
    .Y(_2198_));
 sky130_fd_sc_hd__a2bb2o_1 _6190_ (.A1_N(_1789_),
    .A2_N(_2096_),
    .B1(_2140_),
    .B2(_2192_),
    .X(_2199_));
 sky130_fd_sc_hd__a2111o_1 _6191_ (.A1(_2099_),
    .A2(_2194_),
    .B1(net126),
    .C1(_2198_),
    .D1(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__inv_2 _6192_ (.A(_2200_),
    .Y(_0007_));
 sky130_fd_sc_hd__o21ai_1 _6193_ (.A1(_2140_),
    .A2(_1792_),
    .B1(_2050_),
    .Y(_2201_));
 sky130_fd_sc_hd__nand2_1 _6194_ (.A(_0072_),
    .B(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__nand2_1 _6195_ (.A(_1792_),
    .B(_1790_),
    .Y(_2203_));
 sky130_fd_sc_hd__nand2_1 _6196_ (.A(_1794_),
    .B(_2203_),
    .Y(_2204_));
 sky130_fd_sc_hd__a221o_1 _6197_ (.A1(_2202_),
    .A2(_2204_),
    .B1(_0081_),
    .B2(_1792_),
    .C1(_2122_),
    .X(_2205_));
 sky130_fd_sc_hd__inv_2 _6198_ (.A(_2205_),
    .Y(_0008_));
 sky130_fd_sc_hd__nand2_1 _6199_ (.A(_1794_),
    .B(_1755_),
    .Y(_2207_));
 sky130_fd_sc_hd__nand2_1 _6200_ (.A(_1797_),
    .B(_2207_),
    .Y(_2208_));
 sky130_fd_sc_hd__mux2_1 _6201_ (.A0(_2208_),
    .A1(_1755_),
    .S(_2098_),
    .X(_2209_));
 sky130_fd_sc_hd__mux2_1 _6202_ (.A0(_2208_),
    .A1(_1755_),
    .S(net132),
    .X(_2210_));
 sky130_fd_sc_hd__a22o_1 _6203_ (.A1(_2140_),
    .A2(_2208_),
    .B1(_2094_),
    .B2(_1755_),
    .X(_2211_));
 sky130_fd_sc_hd__a221o_1 _6204_ (.A1(_2099_),
    .A2(_2209_),
    .B1(_0067_),
    .B2(_2210_),
    .C1(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__nor2_1 _6205_ (.A(net120),
    .B(_2212_),
    .Y(_0009_));
 sky130_fd_sc_hd__o21ai_1 _6206_ (.A1(_2140_),
    .A2(_1754_),
    .B1(_2050_),
    .Y(_2213_));
 sky130_fd_sc_hd__a21oi_1 _6207_ (.A1(_0072_),
    .A2(_2213_),
    .B1(_2035_),
    .Y(_2214_));
 sky130_fd_sc_hd__nand2_1 _6208_ (.A(_1797_),
    .B(_1754_),
    .Y(_2215_));
 sky130_fd_sc_hd__or2b_1 _6209_ (.A(_1798_),
    .B_N(_2215_),
    .X(_2217_));
 sky130_fd_sc_hd__a221oi_1 _6210_ (.A1(_0081_),
    .A2(_1754_),
    .B1(_2214_),
    .B2(_2217_),
    .C1(net120),
    .Y(_0010_));
 sky130_fd_sc_hd__or2_1 _6211_ (.A(_1798_),
    .B(_1752_),
    .X(_2218_));
 sky130_fd_sc_hd__nand2_1 _6212_ (.A(_1800_),
    .B(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__mux2_1 _6213_ (.A0(_2219_),
    .A1(_1750_),
    .S(net138),
    .X(_2220_));
 sky130_fd_sc_hd__mux2_1 _6214_ (.A0(_2220_),
    .A1(_1750_),
    .S(_0074_),
    .X(_2221_));
 sky130_fd_sc_hd__mux2_1 _6215_ (.A0(_2219_),
    .A1(_1750_),
    .S(net132),
    .X(_2222_));
 sky130_fd_sc_hd__mux2_1 _6216_ (.A0(_2221_),
    .A1(_2222_),
    .S(_0067_),
    .X(_2223_));
 sky130_fd_sc_hd__and2_1 _6217_ (.A(_2220_),
    .B(_2099_),
    .X(_2224_));
 sky130_fd_sc_hd__a211o_1 _6218_ (.A1(_2223_),
    .A2(_2104_),
    .B1(_2122_),
    .C1(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__inv_2 _6219_ (.A(_2225_),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2_1 _6220_ (.A(_1800_),
    .B(_1748_),
    .Y(_2227_));
 sky130_fd_sc_hd__nand2_1 _6221_ (.A(_1801_),
    .B(_2227_),
    .Y(_2228_));
 sky130_fd_sc_hd__mux2_1 _6222_ (.A0(_2228_),
    .A1(_1748_),
    .S(_2098_),
    .X(_2229_));
 sky130_fd_sc_hd__and3_1 _6223_ (.A(_0067_),
    .B(net132),
    .C(_1748_),
    .X(_2230_));
 sky130_fd_sc_hd__a221o_1 _6224_ (.A1(_2117_),
    .A2(_2228_),
    .B1(_2094_),
    .B2(_1748_),
    .C1(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__a21o_1 _6225_ (.A1(_2140_),
    .A2(_2228_),
    .B1(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__a211o_1 _6226_ (.A1(_2099_),
    .A2(_2229_),
    .B1(_2122_),
    .C1(_2232_),
    .X(_2233_));
 sky130_fd_sc_hd__inv_2 _6227_ (.A(_2233_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _6228_ (.A(_1802_),
    .Y(_2234_));
 sky130_fd_sc_hd__nand2_1 _6229_ (.A(_1801_),
    .B(_1747_),
    .Y(_2236_));
 sky130_fd_sc_hd__nand2_1 _6230_ (.A(_2234_),
    .B(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__mux2_1 _6231_ (.A0(_2237_),
    .A1(_1747_),
    .S(_2098_),
    .X(_2238_));
 sky130_fd_sc_hd__mux2_1 _6232_ (.A0(_2237_),
    .A1(_1747_),
    .S(net132),
    .X(_2239_));
 sky130_fd_sc_hd__a22o_1 _6233_ (.A1(_0075_),
    .A2(_2237_),
    .B1(_2094_),
    .B2(_1747_),
    .X(_2240_));
 sky130_fd_sc_hd__a221o_1 _6234_ (.A1(_2099_),
    .A2(_2238_),
    .B1(_0067_),
    .B2(_2239_),
    .C1(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__nor2_1 _6235_ (.A(net120),
    .B(_2241_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _6236_ (.A(_1803_),
    .Y(_2242_));
 sky130_fd_sc_hd__nand2_1 _6237_ (.A(_2234_),
    .B(_2242_),
    .Y(_2243_));
 sky130_fd_sc_hd__nand2_1 _6238_ (.A(_2243_),
    .B(_1804_),
    .Y(_2244_));
 sky130_fd_sc_hd__mux2_1 _6239_ (.A0(_2244_),
    .A1(_2242_),
    .S(_2736_),
    .X(_2246_));
 sky130_fd_sc_hd__and2_1 _6240_ (.A(_2244_),
    .B(_0075_),
    .X(_2247_));
 sky130_fd_sc_hd__o21a_1 _6241_ (.A1(_2092_),
    .A2(_2094_),
    .B1(_2242_),
    .X(_2248_));
 sky130_fd_sc_hd__a211o_1 _6242_ (.A1(_2117_),
    .A2(_2244_),
    .B1(_2247_),
    .C1(_2248_),
    .X(_2249_));
 sky130_fd_sc_hd__a211o_1 _6243_ (.A1(_2099_),
    .A2(_2246_),
    .B1(_2122_),
    .C1(_2249_),
    .X(_2250_));
 sky130_fd_sc_hd__inv_2 _6244_ (.A(_2250_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_1 _6245_ (.A(_1804_),
    .B(_1746_),
    .Y(_2251_));
 sky130_fd_sc_hd__nand2_1 _6246_ (.A(_2053_),
    .B(_2251_),
    .Y(_2252_));
 sky130_fd_sc_hd__o21a_1 _6247_ (.A1(_2092_),
    .A2(_2094_),
    .B1(_1746_),
    .X(_2253_));
 sky130_fd_sc_hd__a21oi_1 _6248_ (.A1(_2117_),
    .A2(_2252_),
    .B1(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__mux2_1 _6249_ (.A0(_2252_),
    .A1(_1746_),
    .S(_2736_),
    .X(_2256_));
 sky130_fd_sc_hd__nand2_1 _6250_ (.A(_2256_),
    .B(_2099_),
    .Y(_2257_));
 sky130_fd_sc_hd__nand2_1 _6251_ (.A(_2252_),
    .B(_2140_),
    .Y(_2258_));
 sky130_fd_sc_hd__a41o_1 _6252_ (.A1(_2254_),
    .A2(_2257_),
    .A3(_1696_),
    .A4(_2258_),
    .B1(_0001_),
    .X(_0016_));
 sky130_fd_sc_hd__a21o_1 _6253_ (.A1(_2056_),
    .A2(_0079_),
    .B1(_0001_),
    .X(_0017_));
 sky130_fd_sc_hd__a31o_1 _6254_ (.A1(_2047_),
    .A2(_0079_),
    .A3(_2049_),
    .B1(_0001_),
    .X(_0018_));
 sky130_fd_sc_hd__o21ai_1 _6255_ (.A1(net120),
    .A2(_2042_),
    .B1(net117),
    .Y(_0019_));
 sky130_fd_sc_hd__a31o_1 _6256_ (.A1(_2030_),
    .A2(_2036_),
    .A3(_0079_),
    .B1(_0001_),
    .X(_0020_));
 sky130_fd_sc_hd__a21o_1 _6257_ (.A1(_2081_),
    .A2(_0079_),
    .B1(_0001_),
    .X(_0021_));
 sky130_fd_sc_hd__a21o_1 _6258_ (.A1(_2027_),
    .A2(_0079_),
    .B1(_0001_),
    .X(_0022_));
 sky130_fd_sc_hd__a21o_1 _6259_ (.A1(_1958_),
    .A2(_0079_),
    .B1(_0001_),
    .X(_0023_));
 sky130_fd_sc_hd__o21ai_1 _6260_ (.A1(net120),
    .A2(_2019_),
    .B1(net117),
    .Y(_0025_));
 sky130_fd_sc_hd__mux2_1 _6261_ (.A0(_2031_),
    .A1(net122),
    .S(net119),
    .X(_2260_));
 sky130_fd_sc_hd__clkbuf_2 _6262_ (.A(net123),
    .X(_0026_));
 sky130_fd_sc_hd__or4_1 _6263_ (.A(net35),
    .B(net34),
    .C(net64),
    .D(net63),
    .X(_2261_));
 sky130_fd_sc_hd__or4_1 _6264_ (.A(net39),
    .B(net38),
    .C(net37),
    .D(net36),
    .X(_2262_));
 sky130_fd_sc_hd__or4_1 _6265_ (.A(net58),
    .B(net55),
    .C(net44),
    .D(net33),
    .X(_2263_));
 sky130_fd_sc_hd__or4_1 _6266_ (.A(net62),
    .B(net61),
    .C(net60),
    .D(net59),
    .X(_2264_));
 sky130_fd_sc_hd__or4_2 _6267_ (.A(_2261_),
    .B(_2262_),
    .C(_2263_),
    .D(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__or4_1 _6268_ (.A(_1355_),
    .B(_0926_),
    .C(_1058_),
    .D(_0970_),
    .X(_2266_));
 sky130_fd_sc_hd__or3_1 _6269_ (.A(_1300_),
    .B(_1476_),
    .C(_1443_),
    .X(_2268_));
 sky130_fd_sc_hd__nand2_1 _6270_ (.A(_2686_),
    .B(_3241_),
    .Y(_2269_));
 sky130_fd_sc_hd__or4_1 _6271_ (.A(net43),
    .B(net42),
    .C(net41),
    .D(net40),
    .X(_2270_));
 sky130_fd_sc_hd__or4_1 _6272_ (.A(_1014_),
    .B(net47),
    .C(_2269_),
    .D(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__or4_1 _6273_ (.A(_0059_),
    .B(_2266_),
    .C(_2268_),
    .D(_2271_),
    .X(_2272_));
 sky130_fd_sc_hd__nor2_1 _6274_ (.A(_2265_),
    .B(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__or4_1 _6275_ (.A(net3),
    .B(net2),
    .C(net32),
    .D(net31),
    .X(_2274_));
 sky130_fd_sc_hd__or4_1 _6276_ (.A(net7),
    .B(net6),
    .C(net5),
    .D(net4),
    .X(_2275_));
 sky130_fd_sc_hd__or4_1 _6277_ (.A(net26),
    .B(net23),
    .C(net12),
    .D(net1),
    .X(_2276_));
 sky130_fd_sc_hd__or4_1 _6278_ (.A(net30),
    .B(net29),
    .C(net28),
    .D(net27),
    .X(_2277_));
 sky130_fd_sc_hd__or4_2 _6279_ (.A(_2274_),
    .B(_2275_),
    .C(_2276_),
    .D(_2277_),
    .X(_2279_));
 sky130_fd_sc_hd__or4_1 _6280_ (.A(_1377_),
    .B(_0904_),
    .C(_1080_),
    .D(_0992_),
    .X(_2280_));
 sky130_fd_sc_hd__or4_1 _6281_ (.A(net25),
    .B(_1322_),
    .C(_1498_),
    .D(_1421_),
    .X(_2281_));
 sky130_fd_sc_hd__nand2_1 _6282_ (.A(_2705_),
    .B(_3239_),
    .Y(_2282_));
 sky130_fd_sc_hd__or4_1 _6283_ (.A(net11),
    .B(net10),
    .C(net9),
    .D(net8),
    .X(_2283_));
 sky130_fd_sc_hd__or4_1 _6284_ (.A(_1157_),
    .B(net15),
    .C(_2282_),
    .D(_2283_),
    .X(_2284_));
 sky130_fd_sc_hd__or3_1 _6285_ (.A(_2280_),
    .B(_2281_),
    .C(_2284_),
    .X(_2285_));
 sky130_fd_sc_hd__nor2_1 _6286_ (.A(_2279_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__or4_1 _6287_ (.A(net57),
    .B(_2266_),
    .C(_2268_),
    .D(_2271_),
    .X(_2287_));
 sky130_fd_sc_hd__nor2_1 _6288_ (.A(_2265_),
    .B(_2287_),
    .Y(_2288_));
 sky130_fd_sc_hd__or4_1 _6289_ (.A(_1322_),
    .B(_3302_),
    .C(_1498_),
    .D(_1421_),
    .X(_2290_));
 sky130_fd_sc_hd__or3_1 _6290_ (.A(_2280_),
    .B(_2290_),
    .C(_2284_),
    .X(_2291_));
 sky130_fd_sc_hd__nor2_1 _6291_ (.A(_2279_),
    .B(_2291_),
    .Y(_2292_));
 sky130_fd_sc_hd__a22o_1 _6292_ (.A1(_2273_),
    .A2(_2286_),
    .B1(_2288_),
    .B2(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__or4_1 _6293_ (.A(net16),
    .B(net15),
    .C(_2282_),
    .D(_2283_),
    .X(_2294_));
 sky130_fd_sc_hd__or4_1 _6294_ (.A(net20),
    .B(net19),
    .C(net18),
    .D(net17),
    .X(_2295_));
 sky130_fd_sc_hd__or4_1 _6295_ (.A(net21),
    .B(net25),
    .C(net22),
    .D(net24),
    .X(_2296_));
 sky130_fd_sc_hd__or4_1 _6296_ (.A(_2294_),
    .B(_2295_),
    .C(_2296_),
    .D(_2279_),
    .X(_2297_));
 sky130_fd_sc_hd__or4_1 _6297_ (.A(net48),
    .B(net47),
    .C(_2269_),
    .D(_2270_),
    .X(_2298_));
 sky130_fd_sc_hd__or4_1 _6298_ (.A(net52),
    .B(net51),
    .C(net50),
    .D(net49),
    .X(_2299_));
 sky130_fd_sc_hd__or4_1 _6299_ (.A(net53),
    .B(net57),
    .C(net54),
    .D(net56),
    .X(_2301_));
 sky130_fd_sc_hd__or4_1 _6300_ (.A(_2298_),
    .B(_2299_),
    .C(_2301_),
    .D(_2265_),
    .X(_2302_));
 sky130_fd_sc_hd__nor2_1 _6301_ (.A(net25),
    .B(_0059_),
    .Y(_2303_));
 sky130_fd_sc_hd__nor2_1 _6302_ (.A(net57),
    .B(_3302_),
    .Y(_2304_));
 sky130_fd_sc_hd__nor2_4 _6303_ (.A(_2303_),
    .B(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__inv_2 _6304_ (.A(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__and4_1 _6305_ (.A(_3106_),
    .B(_3298_),
    .C(_3282_),
    .D(_3043_),
    .X(_2307_));
 sky130_fd_sc_hd__and3_1 _6306_ (.A(_2307_),
    .B(_3010_),
    .C(_3217_),
    .X(_2308_));
 sky130_fd_sc_hd__or4_1 _6307_ (.A(net53),
    .B(net54),
    .C(_0059_),
    .D(net56),
    .X(_2309_));
 sky130_fd_sc_hd__or4_1 _6308_ (.A(_2298_),
    .B(_2299_),
    .C(_2309_),
    .D(_2265_),
    .X(_2310_));
 sky130_fd_sc_hd__or4_1 _6309_ (.A(net21),
    .B(net22),
    .C(_3302_),
    .D(net24),
    .X(_2312_));
 sky130_fd_sc_hd__or4_1 _6310_ (.A(_2294_),
    .B(_2295_),
    .C(_2312_),
    .D(_2279_),
    .X(_2313_));
 sky130_fd_sc_hd__o2bb2a_1 _6311_ (.A1_N(_2306_),
    .A2_N(_2308_),
    .B1(_2310_),
    .B2(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__o21ai_1 _6312_ (.A1(_2297_),
    .A2(_2302_),
    .B1(_2314_),
    .Y(_2315_));
 sky130_fd_sc_hd__or2b_1 _6313_ (.A(_2293_),
    .B_N(_2315_),
    .X(_2316_));
 sky130_fd_sc_hd__buf_1 _6314_ (.A(_2316_),
    .X(inv_f_c));
 sky130_fd_sc_hd__and2_1 _6315_ (.A(_0073_),
    .B(net67),
    .X(_2317_));
 sky130_fd_sc_hd__nor3_1 _6316_ (.A(_2032_),
    .B(_2305_),
    .C(_2317_),
    .Y(_2318_));
 sky130_fd_sc_hd__a211o_1 _6317_ (.A1(_3302_),
    .A2(_0059_),
    .B1(_2318_),
    .C1(inv_f_c),
    .X(_2319_));
 sky130_fd_sc_hd__inv_2 _6318_ (.A(_2319_),
    .Y(\out_f_c[31] ));
 sky130_fd_sc_hd__nand2_1 _6319_ (.A(_3055_),
    .B(_3308_),
    .Y(\M00[0] ));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(_3067_),
    .B(_3080_),
    .Y(_2321_));
 sky130_fd_sc_hd__xor2_1 _6321_ (.A(_3055_),
    .B(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__xnor2_1 _6322_ (.A(_3308_),
    .B(_2321_),
    .Y(_2323_));
 sky130_fd_sc_hd__inv_2 _6323_ (.A(_3301_),
    .Y(_2324_));
 sky130_fd_sc_hd__clkbuf_4 _6324_ (.A(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__a2bb2o_1 _6325_ (.A1_N(_2322_),
    .A2_N(_0058_),
    .B1(_2323_),
    .B2(_2325_),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _6326_ (.A0(_2326_),
    .A1(_2321_),
    .S(_2305_),
    .X(_2327_));
 sky130_fd_sc_hd__clkbuf_1 _6327_ (.A(_2327_),
    .X(\M00[1] ));
 sky130_fd_sc_hd__clkbuf_4 _6328_ (.A(_2306_),
    .X(_2328_));
 sky130_fd_sc_hd__inv_2 _6329_ (.A(_0058_),
    .Y(_2330_));
 sky130_fd_sc_hd__clkbuf_4 _6330_ (.A(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__clkbuf_4 _6331_ (.A(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__or2_1 _6332_ (.A(_3081_),
    .B(_3043_),
    .X(_2333_));
 sky130_fd_sc_hd__clkbuf_4 _6333_ (.A(_2325_),
    .X(_2334_));
 sky130_fd_sc_hd__xor2_1 _6334_ (.A(_3309_),
    .B(_3043_),
    .X(_2335_));
 sky130_fd_sc_hd__a32o_1 _6335_ (.A1(_2332_),
    .A2(_3082_),
    .A3(_2333_),
    .B1(_2334_),
    .B2(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__clkbuf_4 _6336_ (.A(_2328_),
    .X(_2337_));
 sky130_fd_sc_hd__nand2_1 _6337_ (.A(_2336_),
    .B(_2337_),
    .Y(_2338_));
 sky130_fd_sc_hd__o21ai_1 _6338_ (.A1(_3043_),
    .A2(_2328_),
    .B1(_2338_),
    .Y(\M00[2] ));
 sky130_fd_sc_hd__or2_1 _6339_ (.A(_3106_),
    .B(_3083_),
    .X(_2340_));
 sky130_fd_sc_hd__xor2_1 _6340_ (.A(_3310_),
    .B(_3106_),
    .X(_2341_));
 sky130_fd_sc_hd__a32o_1 _6341_ (.A1(_2332_),
    .A2(_3107_),
    .A3(_2340_),
    .B1(_2334_),
    .B2(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__nand2_1 _6342_ (.A(_3038_),
    .B(_3023_),
    .Y(_2343_));
 sky130_fd_sc_hd__or2_1 _6343_ (.A(_2343_),
    .B(_3106_),
    .X(_2344_));
 sky130_fd_sc_hd__clkbuf_4 _6344_ (.A(_2305_),
    .X(_2345_));
 sky130_fd_sc_hd__nand2_1 _6345_ (.A(_3106_),
    .B(_2343_),
    .Y(_2346_));
 sky130_fd_sc_hd__and3_1 _6346_ (.A(_2344_),
    .B(_2345_),
    .C(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__a21o_1 _6347_ (.A1(_2342_),
    .A2(_2337_),
    .B1(_2347_),
    .X(\M00[3] ));
 sky130_fd_sc_hd__inv_2 _6348_ (.A(_3008_),
    .Y(_2348_));
 sky130_fd_sc_hd__nand2_1 _6349_ (.A(_3108_),
    .B(_2348_),
    .Y(_2350_));
 sky130_fd_sc_hd__or2_1 _6350_ (.A(_2348_),
    .B(_3108_),
    .X(_2351_));
 sky130_fd_sc_hd__or2_1 _6351_ (.A(_2348_),
    .B(_3311_),
    .X(_2352_));
 sky130_fd_sc_hd__nand2_1 _6352_ (.A(_3311_),
    .B(_2348_),
    .Y(_2353_));
 sky130_fd_sc_hd__and2_1 _6353_ (.A(_2352_),
    .B(_2353_),
    .X(_2354_));
 sky130_fd_sc_hd__a32o_1 _6354_ (.A1(_2332_),
    .A2(_2350_),
    .A3(_2351_),
    .B1(_2334_),
    .B2(_2354_),
    .X(_2355_));
 sky130_fd_sc_hd__nand2_1 _6355_ (.A(_3102_),
    .B(_3093_),
    .Y(_2356_));
 sky130_fd_sc_hd__nand2_1 _6356_ (.A(_2344_),
    .B(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__or2_1 _6357_ (.A(_3008_),
    .B(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__nand2_1 _6358_ (.A(_2357_),
    .B(_3008_),
    .Y(_2359_));
 sky130_fd_sc_hd__and3_1 _6359_ (.A(_2358_),
    .B(_2345_),
    .C(_2359_),
    .X(_2361_));
 sky130_fd_sc_hd__a21o_1 _6360_ (.A1(_2355_),
    .A2(_2337_),
    .B1(_2361_),
    .X(\M00[4] ));
 sky130_fd_sc_hd__clkbuf_4 _6361_ (.A(_2305_),
    .X(_2362_));
 sky130_fd_sc_hd__nand2_1 _6362_ (.A(_3005_),
    .B(_2987_),
    .Y(_2363_));
 sky130_fd_sc_hd__nand2_1 _6363_ (.A(_2359_),
    .B(_2363_),
    .Y(_2364_));
 sky130_fd_sc_hd__or2_1 _6364_ (.A(_2969_),
    .B(_2364_),
    .X(_2365_));
 sky130_fd_sc_hd__nand2_1 _6365_ (.A(_2364_),
    .B(_2969_),
    .Y(_2366_));
 sky130_fd_sc_hd__nand2_1 _6366_ (.A(_2350_),
    .B(_3006_),
    .Y(_2367_));
 sky130_fd_sc_hd__xor2_1 _6367_ (.A(_2969_),
    .B(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__nand2_1 _6368_ (.A(_2353_),
    .B(_3007_),
    .Y(_2369_));
 sky130_fd_sc_hd__xnor2_1 _6369_ (.A(_2969_),
    .B(_2369_),
    .Y(_2371_));
 sky130_fd_sc_hd__a2bb2o_1 _6370_ (.A1_N(_2368_),
    .A2_N(_0058_),
    .B1(_2371_),
    .B2(_2324_),
    .X(_2372_));
 sky130_fd_sc_hd__and2_1 _6371_ (.A(_2372_),
    .B(_2328_),
    .X(_2373_));
 sky130_fd_sc_hd__a31o_1 _6372_ (.A1(_2362_),
    .A2(_2365_),
    .A3(_2366_),
    .B1(_2373_),
    .X(\M00[5] ));
 sky130_fd_sc_hd__nand2_1 _6373_ (.A(_2943_),
    .B(_2966_),
    .Y(_2374_));
 sky130_fd_sc_hd__nand2_1 _6374_ (.A(_2366_),
    .B(_2374_),
    .Y(_2375_));
 sky130_fd_sc_hd__or2_1 _6375_ (.A(_2855_),
    .B(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__nand2_1 _6376_ (.A(_2375_),
    .B(_2855_),
    .Y(_2377_));
 sky130_fd_sc_hd__a21bo_1 _6377_ (.A1(_3108_),
    .A2(_3009_),
    .B1_N(_3109_),
    .X(_2378_));
 sky130_fd_sc_hd__inv_2 _6378_ (.A(_2855_),
    .Y(_2379_));
 sky130_fd_sc_hd__nand2_1 _6379_ (.A(_2378_),
    .B(_2379_),
    .Y(_2381_));
 sky130_fd_sc_hd__or2_1 _6380_ (.A(_2379_),
    .B(_2378_),
    .X(_2382_));
 sky130_fd_sc_hd__a21bo_1 _6381_ (.A1(_3311_),
    .A2(_3009_),
    .B1_N(_0036_),
    .X(_2383_));
 sky130_fd_sc_hd__or2_1 _6382_ (.A(_2379_),
    .B(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__nand2_1 _6383_ (.A(_2383_),
    .B(_2379_),
    .Y(_2385_));
 sky130_fd_sc_hd__and2_1 _6384_ (.A(_2384_),
    .B(_2385_),
    .X(_2386_));
 sky130_fd_sc_hd__a32o_1 _6385_ (.A1(_2331_),
    .A2(_2381_),
    .A3(_2382_),
    .B1(_2325_),
    .B2(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__and2_1 _6386_ (.A(_2387_),
    .B(_2328_),
    .X(_2388_));
 sky130_fd_sc_hd__a31o_1 _6387_ (.A1(_2362_),
    .A2(_2376_),
    .A3(_2377_),
    .B1(_2388_),
    .X(\M00[6] ));
 sky130_fd_sc_hd__nand2_1 _6388_ (.A(_2381_),
    .B(_2853_),
    .Y(_2389_));
 sky130_fd_sc_hd__xnor2_1 _6389_ (.A(_2919_),
    .B(_2389_),
    .Y(_2391_));
 sky130_fd_sc_hd__nand2_1 _6390_ (.A(_2385_),
    .B(_2854_),
    .Y(_2392_));
 sky130_fd_sc_hd__xnor2_1 _6391_ (.A(_2919_),
    .B(_2392_),
    .Y(_2393_));
 sky130_fd_sc_hd__a22o_1 _6392_ (.A1(_2332_),
    .A2(_2391_),
    .B1(_2334_),
    .B2(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__nand2_1 _6393_ (.A(_2852_),
    .B(_2796_),
    .Y(_2395_));
 sky130_fd_sc_hd__nand2_1 _6394_ (.A(_2377_),
    .B(_2395_),
    .Y(_2396_));
 sky130_fd_sc_hd__or2_1 _6395_ (.A(_2919_),
    .B(_2396_),
    .X(_2397_));
 sky130_fd_sc_hd__nand2_1 _6396_ (.A(_2396_),
    .B(_2919_),
    .Y(_2398_));
 sky130_fd_sc_hd__and3_1 _6397_ (.A(_2397_),
    .B(_2345_),
    .C(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__a21o_1 _6398_ (.A1(_2394_),
    .A2(_2337_),
    .B1(_2399_),
    .X(\M00[7] ));
 sky130_fd_sc_hd__inv_2 _6399_ (.A(_3193_),
    .Y(_2401_));
 sky130_fd_sc_hd__nand2_1 _6400_ (.A(_3112_),
    .B(_2401_),
    .Y(_2402_));
 sky130_fd_sc_hd__or2_1 _6401_ (.A(_2401_),
    .B(_3112_),
    .X(_2403_));
 sky130_fd_sc_hd__or2_1 _6402_ (.A(_2401_),
    .B(_0039_),
    .X(_2404_));
 sky130_fd_sc_hd__nand2_1 _6403_ (.A(_0039_),
    .B(_2401_),
    .Y(_2405_));
 sky130_fd_sc_hd__and2_1 _6404_ (.A(_2404_),
    .B(_2405_),
    .X(_2406_));
 sky130_fd_sc_hd__a32o_1 _6405_ (.A1(_2332_),
    .A2(_2402_),
    .A3(_2403_),
    .B1(_2334_),
    .B2(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__nand2_1 _6406_ (.A(_2916_),
    .B(_2883_),
    .Y(_2408_));
 sky130_fd_sc_hd__nand2_1 _6407_ (.A(_2398_),
    .B(_2408_),
    .Y(_2409_));
 sky130_fd_sc_hd__or2_1 _6408_ (.A(_3193_),
    .B(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__nand2_1 _6409_ (.A(_2409_),
    .B(_3193_),
    .Y(_2412_));
 sky130_fd_sc_hd__and3_1 _6410_ (.A(_2410_),
    .B(_2345_),
    .C(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__a21o_1 _6411_ (.A1(_2407_),
    .A2(_2337_),
    .B1(_2413_),
    .X(\M00[8] ));
 sky130_fd_sc_hd__nand2_1 _6412_ (.A(_2402_),
    .B(_3191_),
    .Y(_2414_));
 sky130_fd_sc_hd__xnor2_1 _6413_ (.A(_3175_),
    .B(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__nand2_1 _6414_ (.A(_2405_),
    .B(_3192_),
    .Y(_2416_));
 sky130_fd_sc_hd__xnor2_1 _6415_ (.A(_3175_),
    .B(_2416_),
    .Y(_2417_));
 sky130_fd_sc_hd__a22o_1 _6416_ (.A1(_2332_),
    .A2(_2415_),
    .B1(_2334_),
    .B2(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__nand2_1 _6417_ (.A(_3190_),
    .B(_3183_),
    .Y(_2419_));
 sky130_fd_sc_hd__nand2_1 _6418_ (.A(_2412_),
    .B(_2419_),
    .Y(_2420_));
 sky130_fd_sc_hd__or2_1 _6419_ (.A(_3175_),
    .B(_2420_),
    .X(_2422_));
 sky130_fd_sc_hd__nand2_1 _6420_ (.A(_2420_),
    .B(_3175_),
    .Y(_2423_));
 sky130_fd_sc_hd__and3_1 _6421_ (.A(_2422_),
    .B(_2345_),
    .C(_2423_),
    .X(_2424_));
 sky130_fd_sc_hd__a21o_1 _6422_ (.A1(_2418_),
    .A2(_2337_),
    .B1(_2424_),
    .X(\M00[9] ));
 sky130_fd_sc_hd__a21o_1 _6423_ (.A1(_3112_),
    .A2(_3194_),
    .B1(_3218_),
    .X(_2425_));
 sky130_fd_sc_hd__inv_2 _6424_ (.A(_3204_),
    .Y(_2426_));
 sky130_fd_sc_hd__nand2_1 _6425_ (.A(_2425_),
    .B(_2426_),
    .Y(_2427_));
 sky130_fd_sc_hd__or2_1 _6426_ (.A(_2426_),
    .B(_2425_),
    .X(_2428_));
 sky130_fd_sc_hd__a21bo_1 _6427_ (.A1(_0039_),
    .A2(_3194_),
    .B1_N(_0041_),
    .X(_2429_));
 sky130_fd_sc_hd__or2_1 _6428_ (.A(_2426_),
    .B(_2429_),
    .X(_2430_));
 sky130_fd_sc_hd__nand2_1 _6429_ (.A(_2429_),
    .B(_2426_),
    .Y(_2432_));
 sky130_fd_sc_hd__and2_1 _6430_ (.A(_2430_),
    .B(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__a32o_1 _6431_ (.A1(_2332_),
    .A2(_2427_),
    .A3(_2428_),
    .B1(_2334_),
    .B2(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__nand2_1 _6432_ (.A(_3172_),
    .B(_3166_),
    .Y(_2435_));
 sky130_fd_sc_hd__nand2_1 _6433_ (.A(_2423_),
    .B(_2435_),
    .Y(_2436_));
 sky130_fd_sc_hd__or2_1 _6434_ (.A(_3204_),
    .B(_2436_),
    .X(_2437_));
 sky130_fd_sc_hd__nand2_1 _6435_ (.A(_2436_),
    .B(_3204_),
    .Y(_2438_));
 sky130_fd_sc_hd__and3_1 _6436_ (.A(_2437_),
    .B(_2305_),
    .C(_2438_),
    .X(_2439_));
 sky130_fd_sc_hd__a21o_1 _6437_ (.A1(_2434_),
    .A2(_2328_),
    .B1(_2439_),
    .X(\M00[10] ));
 sky130_fd_sc_hd__nand2_1 _6438_ (.A(_2427_),
    .B(_3202_),
    .Y(_2440_));
 sky130_fd_sc_hd__xor2_1 _6439_ (.A(_3214_),
    .B(_2440_),
    .X(_2442_));
 sky130_fd_sc_hd__nand2_1 _6440_ (.A(_2432_),
    .B(_3203_),
    .Y(_2443_));
 sky130_fd_sc_hd__xnor2_1 _6441_ (.A(_3214_),
    .B(_2443_),
    .Y(_2444_));
 sky130_fd_sc_hd__a2bb2o_1 _6442_ (.A1_N(_0058_),
    .A2_N(_2442_),
    .B1(_2325_),
    .B2(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__nand2_1 _6443_ (.A(_3201_),
    .B(_3197_),
    .Y(_2446_));
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(_2438_),
    .B(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__or2_1 _6445_ (.A(_3214_),
    .B(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__nand2_1 _6446_ (.A(_2447_),
    .B(_3214_),
    .Y(_2449_));
 sky130_fd_sc_hd__and3_1 _6447_ (.A(_2448_),
    .B(_2305_),
    .C(_2449_),
    .X(_2450_));
 sky130_fd_sc_hd__a21o_1 _6448_ (.A1(_2337_),
    .A2(_2445_),
    .B1(_2450_),
    .X(\M00[11] ));
 sky130_fd_sc_hd__nand2_1 _6449_ (.A(_3211_),
    .B(_3207_),
    .Y(_2452_));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(_2449_),
    .B(_2452_),
    .Y(_2453_));
 sky130_fd_sc_hd__or2_1 _6451_ (.A(_3138_),
    .B(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__nand2_1 _6452_ (.A(_2453_),
    .B(_3138_),
    .Y(_2455_));
 sky130_fd_sc_hd__inv_2 _6453_ (.A(_3216_),
    .Y(_2456_));
 sky130_fd_sc_hd__a21o_1 _6454_ (.A1(_3112_),
    .A2(_2456_),
    .B1(_3220_),
    .X(_2457_));
 sky130_fd_sc_hd__inv_2 _6455_ (.A(_3138_),
    .Y(_2458_));
 sky130_fd_sc_hd__nand2_1 _6456_ (.A(_2457_),
    .B(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__or2_1 _6457_ (.A(_2458_),
    .B(_2457_),
    .X(_2460_));
 sky130_fd_sc_hd__a21o_1 _6458_ (.A1(_0039_),
    .A2(_2456_),
    .B1(_0043_),
    .X(_2461_));
 sky130_fd_sc_hd__or2_1 _6459_ (.A(_2458_),
    .B(_2461_),
    .X(_2463_));
 sky130_fd_sc_hd__nand2_1 _6460_ (.A(_2461_),
    .B(_2458_),
    .Y(_2464_));
 sky130_fd_sc_hd__and2_1 _6461_ (.A(_2463_),
    .B(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__a32o_1 _6462_ (.A1(_2331_),
    .A2(_2459_),
    .A3(_2460_),
    .B1(_2325_),
    .B2(_2465_),
    .X(_2466_));
 sky130_fd_sc_hd__and2_1 _6463_ (.A(_2466_),
    .B(_2306_),
    .X(_2467_));
 sky130_fd_sc_hd__a31o_1 _6464_ (.A1(_2362_),
    .A2(_2454_),
    .A3(_2455_),
    .B1(_2467_),
    .X(\M00[12] ));
 sky130_fd_sc_hd__nand2_1 _6465_ (.A(_3135_),
    .B(_3130_),
    .Y(_2468_));
 sky130_fd_sc_hd__nand2_1 _6466_ (.A(_2455_),
    .B(_2468_),
    .Y(_2469_));
 sky130_fd_sc_hd__or2_1 _6467_ (.A(_3127_),
    .B(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__nand2_1 _6468_ (.A(_2469_),
    .B(_3127_),
    .Y(_2471_));
 sky130_fd_sc_hd__nand2_1 _6469_ (.A(_2459_),
    .B(_3136_),
    .Y(_2473_));
 sky130_fd_sc_hd__xor2_1 _6470_ (.A(_3127_),
    .B(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__nand2_1 _6471_ (.A(_2464_),
    .B(_3137_),
    .Y(_2475_));
 sky130_fd_sc_hd__xnor2_1 _6472_ (.A(_3127_),
    .B(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__a2bb2o_1 _6473_ (.A1_N(_0058_),
    .A2_N(_2474_),
    .B1(_2324_),
    .B2(_2476_),
    .X(_2477_));
 sky130_fd_sc_hd__and2_1 _6474_ (.A(_2477_),
    .B(_2306_),
    .X(_2478_));
 sky130_fd_sc_hd__a31o_1 _6475_ (.A1(_2470_),
    .A2(_2362_),
    .A3(_2471_),
    .B1(_2478_),
    .X(\M00[13] ));
 sky130_fd_sc_hd__nand2_1 _6476_ (.A(_3124_),
    .B(_3117_),
    .Y(_2479_));
 sky130_fd_sc_hd__nand2_1 _6477_ (.A(_2471_),
    .B(_2479_),
    .Y(_2480_));
 sky130_fd_sc_hd__or2_1 _6478_ (.A(_3149_),
    .B(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__nand2_1 _6479_ (.A(_2480_),
    .B(_3149_),
    .Y(_2483_));
 sky130_fd_sc_hd__inv_2 _6480_ (.A(_3149_),
    .Y(_2484_));
 sky130_fd_sc_hd__a21bo_1 _6481_ (.A1(_2457_),
    .A2(_3139_),
    .B1_N(_3224_),
    .X(_2485_));
 sky130_fd_sc_hd__or2_1 _6482_ (.A(_2484_),
    .B(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__nand2_1 _6483_ (.A(_2485_),
    .B(_2484_),
    .Y(_2487_));
 sky130_fd_sc_hd__and3_1 _6484_ (.A(_2486_),
    .B(_2331_),
    .C(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__a21bo_1 _6485_ (.A1(_2461_),
    .A2(_3139_),
    .B1_N(_0045_),
    .X(_2489_));
 sky130_fd_sc_hd__or2_1 _6486_ (.A(_2484_),
    .B(_2489_),
    .X(_2490_));
 sky130_fd_sc_hd__nand2_1 _6487_ (.A(_2489_),
    .B(_2484_),
    .Y(_2491_));
 sky130_fd_sc_hd__and3_1 _6488_ (.A(_2490_),
    .B(_2325_),
    .C(_2491_),
    .X(_2492_));
 sky130_fd_sc_hd__o21a_1 _6489_ (.A1(_2488_),
    .A2(_2492_),
    .B1(_2328_),
    .X(_2494_));
 sky130_fd_sc_hd__a31o_1 _6490_ (.A1(_2481_),
    .A2(_2362_),
    .A3(_2483_),
    .B1(_2494_),
    .X(\M00[14] ));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(_3146_),
    .B(_3142_),
    .Y(_2495_));
 sky130_fd_sc_hd__nand2_1 _6492_ (.A(_2483_),
    .B(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__or2_1 _6493_ (.A(_3159_),
    .B(_2496_),
    .X(_2497_));
 sky130_fd_sc_hd__nand2_1 _6494_ (.A(_2496_),
    .B(_3159_),
    .Y(_2498_));
 sky130_fd_sc_hd__nand2_1 _6495_ (.A(_2491_),
    .B(_3148_),
    .Y(_2499_));
 sky130_fd_sc_hd__or2_1 _6496_ (.A(_3159_),
    .B(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__nand2_1 _6497_ (.A(_2499_),
    .B(_3159_),
    .Y(_2501_));
 sky130_fd_sc_hd__a21o_1 _6498_ (.A1(_2500_),
    .A2(_2501_),
    .B1(_3301_),
    .X(_2502_));
 sky130_fd_sc_hd__nand2_1 _6499_ (.A(_2502_),
    .B(_0058_),
    .Y(_2504_));
 sky130_fd_sc_hd__nand2_1 _6500_ (.A(_2487_),
    .B(_3147_),
    .Y(_2505_));
 sky130_fd_sc_hd__xor2_1 _6501_ (.A(_3159_),
    .B(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__nand2_1 _6502_ (.A(_2506_),
    .B(_2332_),
    .Y(_2507_));
 sky130_fd_sc_hd__and3_1 _6503_ (.A(_2504_),
    .B(_2306_),
    .C(_2507_),
    .X(_2508_));
 sky130_fd_sc_hd__a31o_1 _6504_ (.A1(_2497_),
    .A2(_2362_),
    .A3(_2498_),
    .B1(_2508_),
    .X(\M00[15] ));
 sky130_fd_sc_hd__nand2_1 _6505_ (.A(_3156_),
    .B(_3152_),
    .Y(_2509_));
 sky130_fd_sc_hd__nand2_1 _6506_ (.A(_2498_),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__or2_1 _6507_ (.A(_3279_),
    .B(_2510_),
    .X(_2511_));
 sky130_fd_sc_hd__nand2_1 _6508_ (.A(_2510_),
    .B(_3279_),
    .Y(_2512_));
 sky130_fd_sc_hd__inv_2 _6509_ (.A(_3279_),
    .Y(_2514_));
 sky130_fd_sc_hd__or2_1 _6510_ (.A(_2514_),
    .B(_3227_),
    .X(_2515_));
 sky130_fd_sc_hd__nand2_1 _6511_ (.A(_3227_),
    .B(_2514_),
    .Y(_2516_));
 sky130_fd_sc_hd__or2_1 _6512_ (.A(_2514_),
    .B(_0047_),
    .X(_2517_));
 sky130_fd_sc_hd__nand2_1 _6513_ (.A(_0047_),
    .B(_2514_),
    .Y(_2518_));
 sky130_fd_sc_hd__and2_1 _6514_ (.A(_2517_),
    .B(_2518_),
    .X(_2519_));
 sky130_fd_sc_hd__a32o_1 _6515_ (.A1(_2331_),
    .A2(_2515_),
    .A3(_2516_),
    .B1(_2325_),
    .B2(_2519_),
    .X(_2520_));
 sky130_fd_sc_hd__and2_1 _6516_ (.A(_2520_),
    .B(_2306_),
    .X(_2521_));
 sky130_fd_sc_hd__a31o_1 _6517_ (.A1(_2511_),
    .A2(_2362_),
    .A3(_2512_),
    .B1(_2521_),
    .X(\M00[16] ));
 sky130_fd_sc_hd__nand2_1 _6518_ (.A(_3276_),
    .B(_3274_),
    .Y(_2522_));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(_2512_),
    .B(_2522_),
    .Y(_2524_));
 sky130_fd_sc_hd__or2_1 _6520_ (.A(_3271_),
    .B(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__nand2_1 _6521_ (.A(_2524_),
    .B(_3271_),
    .Y(_2526_));
 sky130_fd_sc_hd__inv_2 _6522_ (.A(_3271_),
    .Y(_2527_));
 sky130_fd_sc_hd__nand2_1 _6523_ (.A(_2516_),
    .B(_3277_),
    .Y(_2528_));
 sky130_fd_sc_hd__or2_1 _6524_ (.A(_2527_),
    .B(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__nand2_1 _6525_ (.A(_2528_),
    .B(_2527_),
    .Y(_2530_));
 sky130_fd_sc_hd__nand2_1 _6526_ (.A(_2518_),
    .B(_3278_),
    .Y(_2531_));
 sky130_fd_sc_hd__xor2_1 _6527_ (.A(_2527_),
    .B(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__a32o_1 _6528_ (.A1(_2331_),
    .A2(_2529_),
    .A3(_2530_),
    .B1(_2325_),
    .B2(_2532_),
    .X(_2533_));
 sky130_fd_sc_hd__and2_1 _6529_ (.A(_2533_),
    .B(_2306_),
    .X(_2535_));
 sky130_fd_sc_hd__a31o_1 _6530_ (.A1(_2525_),
    .A2(_2362_),
    .A3(_2526_),
    .B1(_2535_),
    .X(\M00[17] ));
 sky130_fd_sc_hd__nand2_1 _6531_ (.A(_3268_),
    .B(_3266_),
    .Y(_2536_));
 sky130_fd_sc_hd__o21a_1 _6532_ (.A1(_2522_),
    .A2(_2527_),
    .B1(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__o21ai_1 _6533_ (.A1(_2527_),
    .A2(_2512_),
    .B1(_2537_),
    .Y(_2538_));
 sky130_fd_sc_hd__or2_1 _6534_ (.A(_3259_),
    .B(_2538_),
    .X(_2539_));
 sky130_fd_sc_hd__nand2_1 _6535_ (.A(_2538_),
    .B(_3259_),
    .Y(_2540_));
 sky130_fd_sc_hd__inv_2 _6536_ (.A(_3259_),
    .Y(_2541_));
 sky130_fd_sc_hd__a21bo_1 _6537_ (.A1(_3227_),
    .A2(_3280_),
    .B1_N(_3287_),
    .X(_2542_));
 sky130_fd_sc_hd__or2_1 _6538_ (.A(_2541_),
    .B(_2542_),
    .X(_2543_));
 sky130_fd_sc_hd__nand2_1 _6539_ (.A(_2542_),
    .B(_2541_),
    .Y(_2545_));
 sky130_fd_sc_hd__and3_1 _6540_ (.A(_2543_),
    .B(_2331_),
    .C(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__a21bo_1 _6541_ (.A1(_0047_),
    .A2(_3280_),
    .B1_N(_0050_),
    .X(_2547_));
 sky130_fd_sc_hd__or2_1 _6542_ (.A(_2541_),
    .B(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__nand2_1 _6543_ (.A(_2547_),
    .B(_2541_),
    .Y(_2549_));
 sky130_fd_sc_hd__and3_1 _6544_ (.A(_2548_),
    .B(_2324_),
    .C(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__o21a_1 _6545_ (.A1(_2546_),
    .A2(_2550_),
    .B1(_2328_),
    .X(_2551_));
 sky130_fd_sc_hd__a31o_1 _6546_ (.A1(_2539_),
    .A2(_2362_),
    .A3(_2540_),
    .B1(_2551_),
    .X(\M00[18] ));
 sky130_fd_sc_hd__inv_2 _6547_ (.A(_3264_),
    .Y(_2552_));
 sky130_fd_sc_hd__nand2_1 _6548_ (.A(_2545_),
    .B(_3257_),
    .Y(_2553_));
 sky130_fd_sc_hd__or2_1 _6549_ (.A(_2552_),
    .B(_2553_),
    .X(_2555_));
 sky130_fd_sc_hd__nand2_1 _6550_ (.A(_2553_),
    .B(_2552_),
    .Y(_2556_));
 sky130_fd_sc_hd__nand2_1 _6551_ (.A(_2549_),
    .B(_3258_),
    .Y(_2557_));
 sky130_fd_sc_hd__xor2_1 _6552_ (.A(_2552_),
    .B(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__a32o_1 _6553_ (.A1(_2555_),
    .A2(_2332_),
    .A3(_2556_),
    .B1(_2334_),
    .B2(_2558_),
    .X(_2559_));
 sky130_fd_sc_hd__or2b_1 _6554_ (.A(_3255_),
    .B_N(_3256_),
    .X(_2560_));
 sky130_fd_sc_hd__a21oi_1 _6555_ (.A1(_2540_),
    .A2(_2560_),
    .B1(_2552_),
    .Y(_2561_));
 sky130_fd_sc_hd__a31o_1 _6556_ (.A1(_2540_),
    .A2(_2552_),
    .A3(_2560_),
    .B1(_2306_),
    .X(_2562_));
 sky130_fd_sc_hd__o2bb2ai_1 _6557_ (.A1_N(_2337_),
    .A2_N(_2559_),
    .B1(_2561_),
    .B2(_2562_),
    .Y(\M00[19] ));
 sky130_fd_sc_hd__and4_1 _6558_ (.A(_3264_),
    .B(_3279_),
    .C(_3259_),
    .D(_3271_),
    .X(_2563_));
 sky130_fd_sc_hd__nand2_1 _6559_ (.A(_2510_),
    .B(_2563_),
    .Y(_2565_));
 sky130_fd_sc_hd__or2b_1 _6560_ (.A(_3260_),
    .B_N(_3261_),
    .X(_2566_));
 sky130_fd_sc_hd__or2_1 _6561_ (.A(_2560_),
    .B(_2552_),
    .X(_2567_));
 sky130_fd_sc_hd__o311a_1 _6562_ (.A1(_2552_),
    .A2(_2541_),
    .A3(_2537_),
    .B1(_2566_),
    .C1(_2567_),
    .X(_2568_));
 sky130_fd_sc_hd__nand2_1 _6563_ (.A(_2565_),
    .B(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__or2_1 _6564_ (.A(_3237_),
    .B(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__nand2_1 _6565_ (.A(_2569_),
    .B(_3237_),
    .Y(_2571_));
 sky130_fd_sc_hd__inv_2 _6566_ (.A(_3237_),
    .Y(_2572_));
 sky130_fd_sc_hd__inv_2 _6567_ (.A(_3281_),
    .Y(_2573_));
 sky130_fd_sc_hd__a21bo_1 _6568_ (.A1(_3227_),
    .A2(_2573_),
    .B1_N(_3288_),
    .X(_2574_));
 sky130_fd_sc_hd__or2_1 _6569_ (.A(_2572_),
    .B(_2574_),
    .X(_2576_));
 sky130_fd_sc_hd__nand2_1 _6570_ (.A(_2574_),
    .B(_2572_),
    .Y(_2577_));
 sky130_fd_sc_hd__and3_1 _6571_ (.A(_2576_),
    .B(_2331_),
    .C(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__a21bo_1 _6572_ (.A1(_0047_),
    .A2(_2573_),
    .B1_N(_0051_),
    .X(_2579_));
 sky130_fd_sc_hd__or2_1 _6573_ (.A(_2572_),
    .B(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__nand2_1 _6574_ (.A(_2579_),
    .B(_2572_),
    .Y(_2581_));
 sky130_fd_sc_hd__and3_1 _6575_ (.A(_2580_),
    .B(_2324_),
    .C(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__o21a_1 _6576_ (.A1(_2578_),
    .A2(_2582_),
    .B1(_2328_),
    .X(_2583_));
 sky130_fd_sc_hd__a31o_1 _6577_ (.A1(_2570_),
    .A2(_2345_),
    .A3(_2571_),
    .B1(_2583_),
    .X(\M00[20] ));
 sky130_fd_sc_hd__or2b_1 _6578_ (.A(_3233_),
    .B_N(_3234_),
    .X(_2584_));
 sky130_fd_sc_hd__nand2_1 _6579_ (.A(_2571_),
    .B(_2584_),
    .Y(_2586_));
 sky130_fd_sc_hd__or2_1 _6580_ (.A(_3232_),
    .B(_2586_),
    .X(_2587_));
 sky130_fd_sc_hd__nand2_1 _6581_ (.A(_2586_),
    .B(_3232_),
    .Y(_2588_));
 sky130_fd_sc_hd__inv_2 _6582_ (.A(_3232_),
    .Y(_2589_));
 sky130_fd_sc_hd__nand2_1 _6583_ (.A(_2577_),
    .B(_3235_),
    .Y(_2590_));
 sky130_fd_sc_hd__or2_1 _6584_ (.A(_2589_),
    .B(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__nand2_1 _6585_ (.A(_2590_),
    .B(_2589_),
    .Y(_2592_));
 sky130_fd_sc_hd__nand2_1 _6586_ (.A(_2581_),
    .B(_3236_),
    .Y(_2593_));
 sky130_fd_sc_hd__xor2_1 _6587_ (.A(_2589_),
    .B(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__a32o_1 _6588_ (.A1(_2591_),
    .A2(_2331_),
    .A3(_2592_),
    .B1(_2325_),
    .B2(_2594_),
    .X(_2595_));
 sky130_fd_sc_hd__and2_1 _6589_ (.A(_2595_),
    .B(_2306_),
    .X(_2597_));
 sky130_fd_sc_hd__a31o_1 _6590_ (.A1(_2587_),
    .A2(_2345_),
    .A3(_2588_),
    .B1(_2597_),
    .X(\M00[21] ));
 sky130_fd_sc_hd__nand3_1 _6591_ (.A(_2569_),
    .B(_3232_),
    .C(_3237_),
    .Y(_2598_));
 sky130_fd_sc_hd__or2b_1 _6592_ (.A(_3228_),
    .B_N(_3229_),
    .X(_2599_));
 sky130_fd_sc_hd__o21a_1 _6593_ (.A1(_2584_),
    .A2(_2589_),
    .B1(_2599_),
    .X(_2600_));
 sky130_fd_sc_hd__nand2_1 _6594_ (.A(_2598_),
    .B(_2600_),
    .Y(_2601_));
 sky130_fd_sc_hd__or2_1 _6595_ (.A(_3246_),
    .B(_2601_),
    .X(_2602_));
 sky130_fd_sc_hd__nand2_1 _6596_ (.A(_2601_),
    .B(_3246_),
    .Y(_2603_));
 sky130_fd_sc_hd__inv_2 _6597_ (.A(_3246_),
    .Y(_2604_));
 sky130_fd_sc_hd__a21bo_1 _6598_ (.A1(_2579_),
    .A2(_3238_),
    .B1_N(_0049_),
    .X(_2605_));
 sky130_fd_sc_hd__or2_1 _6599_ (.A(_2604_),
    .B(_2605_),
    .X(_2607_));
 sky130_fd_sc_hd__nand2_1 _6600_ (.A(_2605_),
    .B(_2604_),
    .Y(_2608_));
 sky130_fd_sc_hd__a21bo_1 _6601_ (.A1(_2574_),
    .A2(_3238_),
    .B1_N(_3285_),
    .X(_2609_));
 sky130_fd_sc_hd__nand2_1 _6602_ (.A(_2609_),
    .B(_2604_),
    .Y(_2610_));
 sky130_fd_sc_hd__and2_1 _6603_ (.A(_2610_),
    .B(_2330_),
    .X(_2611_));
 sky130_fd_sc_hd__or2_1 _6604_ (.A(_2604_),
    .B(_2609_),
    .X(_2612_));
 sky130_fd_sc_hd__a32o_1 _6605_ (.A1(_2607_),
    .A2(_2324_),
    .A3(_2608_),
    .B1(_2611_),
    .B2(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__and2_1 _6606_ (.A(_2613_),
    .B(_2306_),
    .X(_2614_));
 sky130_fd_sc_hd__a31o_1 _6607_ (.A1(_2602_),
    .A2(_2345_),
    .A3(_2603_),
    .B1(_2614_),
    .X(\M00[22] ));
 sky130_fd_sc_hd__or2_1 _6608_ (.A(_3240_),
    .B(_3242_),
    .X(_2615_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(_2603_),
    .B(_2615_),
    .Y(_2617_));
 sky130_fd_sc_hd__nand2_1 _6610_ (.A(_2617_),
    .B(_3252_),
    .Y(_2618_));
 sky130_fd_sc_hd__inv_2 _6611_ (.A(_3252_),
    .Y(_2619_));
 sky130_fd_sc_hd__nand3_1 _6612_ (.A(_2603_),
    .B(_2619_),
    .C(_2615_),
    .Y(_2620_));
 sky130_fd_sc_hd__nand2_1 _6613_ (.A(_2618_),
    .B(_2620_),
    .Y(_2621_));
 sky130_fd_sc_hd__nand2_1 _6614_ (.A(_2610_),
    .B(_3244_),
    .Y(_2622_));
 sky130_fd_sc_hd__or2_1 _6615_ (.A(_2619_),
    .B(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__nand2_1 _6616_ (.A(_2622_),
    .B(_2619_),
    .Y(_2624_));
 sky130_fd_sc_hd__nand2_1 _6617_ (.A(_2608_),
    .B(_3245_),
    .Y(_2625_));
 sky130_fd_sc_hd__xor2_1 _6618_ (.A(_2619_),
    .B(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__a32o_1 _6619_ (.A1(_2623_),
    .A2(_2332_),
    .A3(_2624_),
    .B1(_2334_),
    .B2(_2626_),
    .X(_2628_));
 sky130_fd_sc_hd__nand2_1 _6620_ (.A(_2628_),
    .B(_2337_),
    .Y(_2629_));
 sky130_fd_sc_hd__o21ai_1 _6621_ (.A1(_2328_),
    .A2(_2621_),
    .B1(_2629_),
    .Y(\M00[23] ));
 sky130_fd_sc_hd__nor2_1 _6622_ (.A(_2604_),
    .B(_2619_),
    .Y(_2630_));
 sky130_fd_sc_hd__and3_1 _6623_ (.A(_2630_),
    .B(_3232_),
    .C(_3237_),
    .X(_2631_));
 sky130_fd_sc_hd__nand3_1 _6624_ (.A(_2510_),
    .B(_2563_),
    .C(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__or2_1 _6625_ (.A(_3247_),
    .B(_3248_),
    .X(_2633_));
 sky130_fd_sc_hd__o21a_1 _6626_ (.A1(_2615_),
    .A2(_2619_),
    .B1(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__or2b_1 _6627_ (.A(_2568_),
    .B_N(_2631_),
    .X(_2635_));
 sky130_fd_sc_hd__o311a_1 _6628_ (.A1(_2619_),
    .A2(_2604_),
    .A3(_2600_),
    .B1(_2634_),
    .C1(_2635_),
    .X(_2636_));
 sky130_fd_sc_hd__nand2_1 _6629_ (.A(_2632_),
    .B(_2636_),
    .Y(_2638_));
 sky130_fd_sc_hd__or2_1 _6630_ (.A(_3297_),
    .B(_2638_),
    .X(_2639_));
 sky130_fd_sc_hd__nand2_1 _6631_ (.A(_2638_),
    .B(_3297_),
    .Y(_2640_));
 sky130_fd_sc_hd__inv_2 _6632_ (.A(_3297_),
    .Y(_2641_));
 sky130_fd_sc_hd__or2_1 _6633_ (.A(_2641_),
    .B(_3291_),
    .X(_2642_));
 sky130_fd_sc_hd__nand2_1 _6634_ (.A(_3291_),
    .B(_2641_),
    .Y(_2643_));
 sky130_fd_sc_hd__and3_1 _6635_ (.A(_2331_),
    .B(_2642_),
    .C(_2643_),
    .X(_2644_));
 sky130_fd_sc_hd__or2_1 _6636_ (.A(_2641_),
    .B(_0054_),
    .X(_2645_));
 sky130_fd_sc_hd__nand2_1 _6637_ (.A(_0054_),
    .B(_2641_),
    .Y(_2646_));
 sky130_fd_sc_hd__and3_1 _6638_ (.A(_2325_),
    .B(_2645_),
    .C(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__o21a_1 _6639_ (.A1(_2644_),
    .A2(_2647_),
    .B1(_2328_),
    .X(_2649_));
 sky130_fd_sc_hd__a31o_1 _6640_ (.A1(_2639_),
    .A2(_2345_),
    .A3(_2640_),
    .B1(_2649_),
    .X(\M00[24] ));
 sky130_fd_sc_hd__nand3_1 _6641_ (.A(_2643_),
    .B(_1652_),
    .C(_3296_),
    .Y(_2650_));
 sky130_fd_sc_hd__inv_2 _6642_ (.A(_1652_),
    .Y(_2651_));
 sky130_fd_sc_hd__nand2_1 _6643_ (.A(_2646_),
    .B(_3295_),
    .Y(_2652_));
 sky130_fd_sc_hd__xor2_1 _6644_ (.A(_2651_),
    .B(_2652_),
    .X(_2653_));
 sky130_fd_sc_hd__a22oi_1 _6645_ (.A1(_2697_),
    .A2(_2650_),
    .B1(_2653_),
    .B2(_2334_),
    .Y(_2654_));
 sky130_fd_sc_hd__or2b_1 _6646_ (.A(_3294_),
    .B_N(_3292_),
    .X(_2655_));
 sky130_fd_sc_hd__nand2_1 _6647_ (.A(_2640_),
    .B(_2655_),
    .Y(_2656_));
 sky130_fd_sc_hd__nor2_1 _6648_ (.A(_2651_),
    .B(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__and2_1 _6649_ (.A(_2656_),
    .B(_2651_),
    .X(_2659_));
 sky130_fd_sc_hd__o21ai_1 _6650_ (.A1(_2657_),
    .A2(_2659_),
    .B1(_2362_),
    .Y(_2660_));
 sky130_fd_sc_hd__o21ai_1 _6651_ (.A1(_2345_),
    .A2(_2654_),
    .B1(_2660_),
    .Y(\M00[25] ));
 sky130_fd_sc_hd__nor2_1 _6652_ (.A(_2337_),
    .B(_2657_),
    .Y(\M00[26] ));
 sky130_fd_sc_hd__or3_1 _6653_ (.A(_2286_),
    .B(_2288_),
    .C(_2315_),
    .X(_2661_));
 sky130_fd_sc_hd__clkbuf_1 _6654_ (.A(_2661_),
    .X(forward_c));
 sky130_fd_sc_hd__dfrtp_1 _6655_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0002_),
    .RESET_B(net109),
    .Q(net72));
 sky130_fd_sc_hd__dfrtp_1 _6656_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0013_),
    .RESET_B(net109),
    .Q(net83));
 sky130_fd_sc_hd__dfrtp_1 _6657_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0024_),
    .RESET_B(net109),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 _6658_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0027_),
    .RESET_B(net109),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 _6659_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0028_),
    .RESET_B(net109),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_1 _6660_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0029_),
    .RESET_B(net109),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_1 _6661_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0030_),
    .RESET_B(net109),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_1 _6662_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0031_),
    .RESET_B(net109),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 _6663_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0032_),
    .RESET_B(net109),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 _6664_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0033_),
    .RESET_B(net109),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_1 _6665_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0003_),
    .RESET_B(net110),
    .Q(net73));
 sky130_fd_sc_hd__dfrtp_1 _6666_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0004_),
    .RESET_B(net110),
    .Q(net74));
 sky130_fd_sc_hd__dfrtp_1 _6667_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0005_),
    .RESET_B(net110),
    .Q(net75));
 sky130_fd_sc_hd__dfrtp_1 _6668_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0006_),
    .RESET_B(net110),
    .Q(net76));
 sky130_fd_sc_hd__dfrtp_1 _6669_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0007_),
    .RESET_B(net110),
    .Q(net77));
 sky130_fd_sc_hd__dfrtp_1 _6670_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0008_),
    .RESET_B(net110),
    .Q(net78));
 sky130_fd_sc_hd__dfrtp_1 _6671_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0009_),
    .RESET_B(net110),
    .Q(net79));
 sky130_fd_sc_hd__dfrtp_1 _6672_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0010_),
    .RESET_B(net110),
    .Q(net80));
 sky130_fd_sc_hd__dfrtp_1 _6673_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0011_),
    .RESET_B(net110),
    .Q(net81));
 sky130_fd_sc_hd__dfrtp_1 _6674_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0012_),
    .RESET_B(net112),
    .Q(net82));
 sky130_fd_sc_hd__dfrtp_1 _6675_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0014_),
    .RESET_B(net112),
    .Q(net84));
 sky130_fd_sc_hd__dfrtp_1 _6676_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0015_),
    .RESET_B(net112),
    .Q(net85));
 sky130_fd_sc_hd__dfrtp_1 _6677_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0016_),
    .RESET_B(net112),
    .Q(net86));
 sky130_fd_sc_hd__dfrtp_1 _6678_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0017_),
    .RESET_B(net112),
    .Q(net87));
 sky130_fd_sc_hd__dfrtp_1 _6679_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0018_),
    .RESET_B(net112),
    .Q(net88));
 sky130_fd_sc_hd__dfrtp_1 _6680_ (.CLK(clknet_3_6__leaf_clk),
    .D(net121),
    .RESET_B(net112),
    .Q(net89));
 sky130_fd_sc_hd__dfrtp_1 _6681_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0020_),
    .RESET_B(net112),
    .Q(net90));
 sky130_fd_sc_hd__dfrtp_1 _6682_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0021_),
    .RESET_B(net111),
    .Q(net91));
 sky130_fd_sc_hd__dfrtp_1 _6683_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0022_),
    .RESET_B(net111),
    .Q(net92));
 sky130_fd_sc_hd__dfrtp_1 _6684_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0023_),
    .RESET_B(net111),
    .Q(net93));
 sky130_fd_sc_hd__dfrtp_1 _6685_ (.CLK(clknet_3_7__leaf_clk),
    .D(net118),
    .RESET_B(net111),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_1 _6686_ (.CLK(clknet_3_7__leaf_clk),
    .D(net124),
    .RESET_B(net111),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_1 _6687_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0034_),
    .RESET_B(net111),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 _6688_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0035_),
    .RESET_B(net111),
    .Q(net105));
 sky130_fd_sc_hd__dfstp_1 _6689_ (.CLK(clknet_3_7__leaf_clk),
    .D(net185),
    .SET_B(net111),
    .Q(net69));
 sky130_fd_sc_hd__dfrtp_1 _6690_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0001_),
    .RESET_B(net111),
    .Q(net71));
 sky130_fd_sc_hd__dfrtp_1 _6691_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0000_),
    .RESET_B(net111),
    .Q(net70));
 sky130_fd_sc_hd__dfrtp_1 _6692_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[0] ),
    .RESET_B(net107),
    .Q(\M000[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6693_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[1] ),
    .RESET_B(net107),
    .Q(\M000[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6694_ (.CLK(clknet_3_0__leaf_clk),
    .D(\M00[2] ),
    .RESET_B(net106),
    .Q(\M000[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6695_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[3] ),
    .RESET_B(net106),
    .Q(\M000[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6696_ (.CLK(clknet_3_0__leaf_clk),
    .D(\M00[4] ),
    .RESET_B(net106),
    .Q(\M000[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6697_ (.CLK(clknet_3_0__leaf_clk),
    .D(\M00[5] ),
    .RESET_B(net106),
    .Q(\M000[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6698_ (.CLK(clknet_3_0__leaf_clk),
    .D(\M00[6] ),
    .RESET_B(net106),
    .Q(\M000[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6699_ (.CLK(clknet_3_0__leaf_clk),
    .D(\M00[7] ),
    .RESET_B(net106),
    .Q(\M000[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6700_ (.CLK(clknet_3_0__leaf_clk),
    .D(\M00[8] ),
    .RESET_B(net106),
    .Q(\M000[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6701_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[9] ),
    .RESET_B(net106),
    .Q(\M000[9] ));
 sky130_fd_sc_hd__dfrtp_1 _6702_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[10] ),
    .RESET_B(net106),
    .Q(\M000[10] ));
 sky130_fd_sc_hd__dfrtp_1 _6703_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[11] ),
    .RESET_B(net106),
    .Q(\M000[11] ));
 sky130_fd_sc_hd__dfrtp_1 _6704_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[12] ),
    .RESET_B(net107),
    .Q(\M000[12] ));
 sky130_fd_sc_hd__dfrtp_1 _6705_ (.CLK(clknet_3_0__leaf_clk),
    .D(\M00[13] ),
    .RESET_B(net107),
    .Q(\M000[13] ));
 sky130_fd_sc_hd__dfrtp_1 _6706_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[14] ),
    .RESET_B(net107),
    .Q(\M000[14] ));
 sky130_fd_sc_hd__dfrtp_1 _6707_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[15] ),
    .RESET_B(net107),
    .Q(\M000[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6708_ (.CLK(clknet_3_1__leaf_clk),
    .D(\M00[16] ),
    .RESET_B(net107),
    .Q(\M000[16] ));
 sky130_fd_sc_hd__dfrtp_1 _6709_ (.CLK(clknet_3_3__leaf_clk),
    .D(\M00[17] ),
    .RESET_B(net107),
    .Q(\M000[17] ));
 sky130_fd_sc_hd__dfrtp_1 _6710_ (.CLK(clknet_3_3__leaf_clk),
    .D(\M00[18] ),
    .RESET_B(net107),
    .Q(\M000[18] ));
 sky130_fd_sc_hd__dfrtp_1 _6711_ (.CLK(clknet_3_3__leaf_clk),
    .D(\M00[19] ),
    .RESET_B(net108),
    .Q(\M000[19] ));
 sky130_fd_sc_hd__dfrtp_1 _6712_ (.CLK(clknet_3_2__leaf_clk),
    .D(\M00[20] ),
    .RESET_B(net108),
    .Q(\M000[20] ));
 sky130_fd_sc_hd__dfrtp_1 _6713_ (.CLK(clknet_3_2__leaf_clk),
    .D(\M00[21] ),
    .RESET_B(net108),
    .Q(\M000[21] ));
 sky130_fd_sc_hd__dfrtp_1 _6714_ (.CLK(clknet_3_2__leaf_clk),
    .D(\M00[22] ),
    .RESET_B(net108),
    .Q(\M000[22] ));
 sky130_fd_sc_hd__dfrtp_1 _6715_ (.CLK(clknet_3_3__leaf_clk),
    .D(\M00[23] ),
    .RESET_B(net108),
    .Q(\M000[23] ));
 sky130_fd_sc_hd__dfrtp_1 _6716_ (.CLK(clknet_3_2__leaf_clk),
    .D(\M00[24] ),
    .RESET_B(net108),
    .Q(\M000[24] ));
 sky130_fd_sc_hd__dfrtp_1 _6717_ (.CLK(clknet_3_3__leaf_clk),
    .D(\M00[25] ),
    .RESET_B(net108),
    .Q(\M000[25] ));
 sky130_fd_sc_hd__dfrtp_1 _6718_ (.CLK(clknet_3_3__leaf_clk),
    .D(\M00[26] ),
    .RESET_B(net108),
    .Q(\M000[26] ));
 sky130_fd_sc_hd__dfrtp_1 _6719_ (.CLK(clknet_3_7__leaf_clk),
    .D(net114),
    .RESET_B(net112),
    .Q(done0_r));
 sky130_fd_sc_hd__conb_1 _6719__114 (.HI(net114));
 sky130_fd_sc_hd__dfrtp_1 _6720_ (.CLK(clknet_3_2__leaf_clk),
    .D(inv_f_c),
    .RESET_B(net108),
    .Q(inv_f));
 sky130_fd_sc_hd__dfrtp_1 _6721_ (.CLK(clknet_3_3__leaf_clk),
    .D(\out_f_c[31] ),
    .RESET_B(net108),
    .Q(\out_f[31] ));
 sky130_fd_sc_hd__dfrtp_1 _6722_ (.CLK(clknet_3_2__leaf_clk),
    .D(forward_c),
    .RESET_B(net113),
    .Q(forward));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(net113),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net113),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net113),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(net113),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net113),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net68),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net184),
    .X(net115));
 sky130_fd_sc_hd__buf_1 hold10 (.A(_0026_),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(forward),
    .X(net125));
 sky130_fd_sc_hd__buf_2 hold12 (.A(net119),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0080_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\M000[0] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0750_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_2720_),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_2721_),
    .X(net131));
 sky130_fd_sc_hd__buf_2 hold18 (.A(_0068_),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_2152_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(inv_f),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_2153_),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\M000[2] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0717_),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0794_),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 hold24 (.A(_0882_),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\M000[3] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_2723_),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_2724_),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_2727_),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_2 hold29 (.A(_2734_),
    .X(net143));
 sky130_fd_sc_hd__buf_1 hold3 (.A(net127),
    .X(net117));
 sky130_fd_sc_hd__buf_1 hold30 (.A(\M000[24] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_2729_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_2730_),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_2731_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\M000[4] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_1174_),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_1246_),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_1316_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_1405_),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_1506_),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0025_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 hold40 (.A(_1763_),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_2118_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_2119_),
    .X(net156));
 sky130_fd_sc_hd__buf_1 hold43 (.A(\M000[26] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0838_),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\M000[5] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_1098_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_1100_),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_1103_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_1105_),
    .X(net163));
 sky130_fd_sc_hd__buf_4 hold5 (.A(net125),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\M000[20] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0204_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0206_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0208_),
    .X(net167));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold54 (.A(_0211_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 hold55 (.A(_0236_),
    .X(net169));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold56 (.A(_1765_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\M000[23] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0133_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0178_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 hold6 (.A(_2073_),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0180_),
    .X(net174));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold61 (.A(_0182_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0275_),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0298_),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_1770_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\M000[25] ),
    .X(net179));
 sky130_fd_sc_hd__buf_1 hold66 (.A(_1760_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\M000[19] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0288_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0377_),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0019_),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net186),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net115),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(done0_r),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\out_f[31] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_2260_),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in1[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(in1[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(in1[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(in1[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(in1[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(in1[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(in1[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(in1[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(in1[24]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(in1[25]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(in1[26]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(in1[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(in1[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(in1[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(in1[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(in1[2]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(in1[30]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(in1[31]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(in1[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(in1[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(in1[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(in1[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(in1[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(in1[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(in1[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(in1[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(in2[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(in2[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(in2[11]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(in2[12]),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(in2[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(in2[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(in2[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(in1[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(in2[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(in2[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(in2[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(in2[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(in2[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(in2[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(in2[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(in2[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(in2[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(in2[24]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(in1[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(in2[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(in2[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(in2[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(in2[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(in2[29]),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(in2[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(in2[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(in2[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(in2[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(in2[4]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input6 (.A(in1[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(in2[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(in2[6]),
    .X(net61));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(in2[7]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input63 (.A(in2[8]),
    .X(net63));
 sky130_fd_sc_hd__dlymetal6s2s_1 input64 (.A(in2[9]),
    .X(net64));
 sky130_fd_sc_hd__dlymetal6s2s_1 input65 (.A(round_m[0]),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(round_m[1]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(round_m[2]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(rst),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(in1[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(in1[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(in1[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(out[6]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(out[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(out[8]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(out[9]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(ov));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(un));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(done));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(inexact));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(inv));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(out[0]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(out[10]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(out[11]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(out[12]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(out[13]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(out[14]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(out[15]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(out[16]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(out[17]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(out[18]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(out[19]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(out[20]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(out[21]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(out[22]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(out[23]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(out[24]));
 sky130_fd_sc_hd__clkbuf_4 output89 (.A(net89),
    .X(out[25]));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(out[26]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(out[27]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(out[28]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(out[29]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(out[2]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(out[30]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(out[31]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(out[3]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(out[4]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(out[5]));
endmodule

